module b10_C( R_BUTTON, G_BUTTON, KEY, START, TEST, RTS, RTR, VOTO0_REG_SCAN_IN, V_IN_3_, V_IN_2_, V_IN_1_, V_IN_0_, STATO_REG_3__SCAN_IN, STATO_REG_2__SCAN_IN, STATO_REG_1__SCAN_IN, STATO_REG_0__SCAN_IN, V_OUT_REG_3__SCAN_IN, V_OUT_REG_2__SCAN_IN, V_OUT_REG_1__SCAN_IN, V_OUT_REG_0__SCAN_IN, SIGN_REG_3__SCAN_IN, VOTO1_REG_SCAN_IN, CTR_REG_SCAN_IN, VOTO3_REG_SCAN_IN, LAST_R_REG_SCAN_IN, CTS_REG_SCAN_IN, VOTO2_REG_SCAN_IN, LAST_G_REG_SCAN_IN, U207, U208, U209, U210, U211, U212, U233, U234, U235, U236, U237, U238, U239, U240, U241, U242, U243); 
input R_BUTTON, G_BUTTON, KEY, START, TEST, RTS, RTR, VOTO0_REG_SCAN_IN, V_IN_3_, V_IN_2_, V_IN_1_, V_IN_0_, STATO_REG_3__SCAN_IN, STATO_REG_2__SCAN_IN, STATO_REG_1__SCAN_IN, STATO_REG_0__SCAN_IN, V_OUT_REG_3__SCAN_IN, V_OUT_REG_2__SCAN_IN, V_OUT_REG_1__SCAN_IN, V_OUT_REG_0__SCAN_IN, SIGN_REG_3__SCAN_IN, VOTO1_REG_SCAN_IN, CTR_REG_SCAN_IN, VOTO3_REG_SCAN_IN, LAST_R_REG_SCAN_IN, CTS_REG_SCAN_IN, VOTO2_REG_SCAN_IN, LAST_G_REG_SCAN_IN; 
output U207, U208, U209, U210, U211, U212, U233, U234, U235, U236, U237, U238, U239, U240, U241, U242, U243; 
wire U200, U201, U202, U203, U204, U205, U206, U213, U214, U215, U216, U217, U218, U219, U220, U221, U222, U223, U224, U225, U226, U227, U228, U229, U230, U231, U232, U244, U245, U246, U247, U248, U249, U250, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, U280, U281, U282, U283, U284, U285, U286, U287, U288, U289, U290, U291, U292, U293, U294, U295, U296, U297, U298, U299, U300, U301, U302, U303, U304, U305, U306, U307, U308, U309, U310, U311, U312, U313, U314, U315, U316, U317, U318, U319, U320, U321, U322, U323, U324, U325, U326, U327, U328, U329, U330, U331, U332, U333, U334, U335, U336, U337, U338, U339, U340, U341, U342, U343, U344, U345, U346, U347, U348, U349, U350, U351, U352, U353, U354, U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U365, U366, U367, U368, U369, U370, U371; 
assign U200 = ~(STATO_REG_3__SCAN_IN | STATO_REG_2__SCAN_IN); 
assign U213 = ~STATO_REG_0__SCAN_IN; 
assign U215 = ~STATO_REG_2__SCAN_IN; 
assign U216 = ~RTR; 
assign U217 = ~STATO_REG_1__SCAN_IN; 
assign U219 = ~RTS; 
assign U221 = ~STATO_REG_3__SCAN_IN; 
assign U222 = ~START; 
assign U224 = ~(STATO_REG_1__SCAN_IN & STATO_REG_0__SCAN_IN); 
assign U226 = ~VOTO1_REG_SCAN_IN; 
assign U227 = ~VOTO2_REG_SCAN_IN; 
assign U230 = ~SIGN_REG_3__SCAN_IN; 
assign U232 = ~KEY; 
assign U247 = ~VOTO3_REG_SCAN_IN; 
assign U248 = ~VOTO0_REG_SCAN_IN; 
assign U251 = ~LAST_R_REG_SCAN_IN; 
assign U254 = ~LAST_G_REG_SCAN_IN; 
assign U257 = ~TEST; 
assign U270 = RTR | STATO_REG_1__SCAN_IN; 
assign U290 = ~(STATO_REG_3__SCAN_IN & STATO_REG_0__SCAN_IN); 
assign U310 = STATO_REG_3__SCAN_IN | STATO_REG_0__SCAN_IN; 
assign U331 = ~(V_IN_3_ & V_IN_2_ & V_IN_0_ & V_IN_1_); 
assign U201 = U213 & STATO_REG_2__SCAN_IN; 
assign U214 = ~(U217 & STATO_REG_0__SCAN_IN); 
assign U220 = ~(U200 & U213); 
assign U223 = ~(START & U200); 
assign U225 = ~(U221 & STATO_REG_1__SCAN_IN); 
assign U228 = ~(U247 & U248 & VOTO1_REG_SCAN_IN & VOTO2_REG_SCAN_IN); 
assign U231 = ~(U215 & STATO_REG_1__SCAN_IN); 
assign U266 = ~U224; 
assign U299 = ~(U217 & STATO_REG_2__SCAN_IN); 
assign U302 = ~(START & U232); 
assign U311 = ~(RTR & U310); 
assign U313 = ~(U213 & STATO_REG_1__SCAN_IN); 
assign U326 = ~(U230 & STATO_REG_3__SCAN_IN); 
assign U333 = ~(U331 & STATO_REG_0__SCAN_IN); 
assign U337 = ~(U213 & STATO_REG_3__SCAN_IN); 
assign U338 = ~(U221 & STATO_REG_0__SCAN_IN); 
assign U354 = ~(U217 & STATO_REG_3__SCAN_IN); 
assign U355 = ~(U219 & STATO_REG_1__SCAN_IN); 
assign U356 = ~(U248 & VOTO2_REG_SCAN_IN); 
assign U357 = ~(U227 & VOTO0_REG_SCAN_IN); 
assign U206 = U231 & U299; 
assign U218 = ~(U201 & STATO_REG_1__SCAN_IN); 
assign U245 = ~(U357 & U356); 
assign U246 = ~(RTR & U217 & U201); 
assign U256 = ~U228; 
assign U258 = ~U220; 
assign U262 = ~U223; 
assign U264 = ~U214; 
assign U265 = ~U231; 
assign U271 = ~U225; 
assign U281 = ~(U213 & U228); 
assign U303 = ~(U224 & U302); 
assign U315 = ~(U217 & U201 & STATO_REG_3__SCAN_IN); 
assign U334 = ~(U270 & U231 & U213); 
assign U336 = ~(U266 & U216 & STATO_REG_2__SCAN_IN); 
assign U339 = ~(U338 & U337); 
assign U202 = START & U258; 
assign U259 = ~U218; 
assign U260 = ~(U219 & U264 & STATO_REG_2__SCAN_IN); 
assign U261 = ~(U215 & U264 & STATO_REG_3__SCAN_IN); 
assign U267 = ~U246; 
assign U269 = ~(U258 & U217); 
assign U272 = ~(U334 & U333 & STATO_REG_3__SCAN_IN); 
assign U273 = ~(U262 & STATO_REG_0__SCAN_IN); 
assign U275 = ~(U256 & U201); 
assign U276 = ~(U258 & U257); 
assign U283 = ~(U339 & STATO_REG_1__SCAN_IN); 
assign U285 = ~(U256 & U221); 
assign U288 = ~(U257 & U217 & U258); 
assign U291 = ~(START & U215 & U264); 
assign U296 = ~(KEY & U226 & U265); 
assign U300 = ~(U355 & U354 & U213 & U206); 
assign U304 = ~(U200 & U303); 
assign U312 = ~(U264 & STATO_REG_3__SCAN_IN); 
assign U316 = ~(RTR & U200 & U264); 
assign U320 = ~(KEY & U227 & U265); 
assign U323 = ~(U265 & U339); 
assign U325 = ~(KEY & U258); 
assign U335 = ~(U271 & U222 & U215); 
assign U341 = ~(U271 & U213); 
assign U344 = ~(U246 & V_OUT_REG_3__SCAN_IN); 
assign U346 = ~(U246 & V_OUT_REG_2__SCAN_IN); 
assign U348 = ~(U246 & V_OUT_REG_1__SCAN_IN); 
assign U350 = ~(U246 & V_OUT_REG_0__SCAN_IN); 
assign U358 = ~U245; 
assign U360 = ~(U245 & U226); 
assign U244 = U336 & U335 & U273; 
assign U252 = ~(KEY & U202 & STATO_REG_1__SCAN_IN); 
assign U263 = ~(U202 & U232); 
assign U268 = ~(RTS & U259); 
assign U277 = ~(U276 & U275); 
assign U286 = ~(U213 & U217 & U285); 
assign U289 = ~(U288 & SIGN_REG_3__SCAN_IN); 
assign U292 = ~(G_BUTTON & U254 & U202); 
assign U294 = ~(U259 & U221); 
assign U301 = ~(U300 & CTR_REG_SCAN_IN); 
assign U314 = ~(U206 & U313 & U312 & U311); 
assign U318 = ~(R_BUTTON & U251 & U202); 
assign U327 = ~(U326 & U325); 
assign U345 = ~(U267 & VOTO3_REG_SCAN_IN); 
assign U347 = ~(U267 & VOTO2_REG_SCAN_IN); 
assign U349 = ~(U267 & VOTO1_REG_SCAN_IN); 
assign U351 = ~(U267 & VOTO0_REG_SCAN_IN); 
assign U359 = ~(U358 & VOTO1_REG_SCAN_IN); 
assign U203 = U269 & U268; 
assign U208 = ~(U260 & U301); 
assign U209 = ~(U290 & U289); 
assign U234 = ~(U345 & U344); 
assign U235 = ~(U347 & U346); 
assign U236 = ~(U349 & U348); 
assign U237 = ~(U351 & U350); 
assign U287 = ~(U218 & U220 & U286); 
assign U295 = ~(U261 & U294); 
assign U309 = ~U252; 
assign U317 = ~(U314 & CTS_REG_SCAN_IN); 
assign U328 = ~(U327 & STATO_REG_1__SCAN_IN); 
assign U361 = ~(U360 & U359); 
assign U364 = ~(U252 & LAST_R_REG_SCAN_IN); 
assign U368 = ~(U252 & LAST_G_REG_SCAN_IN); 
assign U204 = U203 & U261; 
assign U207 = ~(U315 & U246 & U316 & U317); 
assign U229 = ~(U246 & U260 & U272 & U244 & U203); 
assign U297 = ~(V_IN_1_ & U295); 
assign U306 = ~(U266 & U361); 
assign U307 = ~(V_IN_3_ & U295); 
assign U321 = ~(V_IN_2_ & U295); 
assign U329 = ~(V_IN_0_ & U295); 
assign U365 = ~(U309 & R_BUTTON); 
assign U369 = ~(U309 & G_BUTTON); 
assign U205 = U204 & U291; 
assign U240 = ~(U365 & U364); 
assign U242 = ~(U369 & U368); 
assign U255 = ~(U323 & U223 & U204); 
assign U274 = ~U229; 
assign U278 = ~(U213 & U229); 
assign U279 = ~(U277 & U217 & U229); 
assign U282 = ~(U281 & U214 & U229); 
assign U298 = ~(U297 & U296); 
assign U308 = ~(U307 & U306); 
assign U322 = ~(U321 & U320); 
assign U330 = ~(U329 & U328); 
assign U340 = ~(U229 & U225 & STATO_REG_0__SCAN_IN); 
assign U343 = ~(U287 & U229); 
assign U249 = ~(U292 & U263 & U205); 
assign U250 = ~(U205 & U304); 
assign U253 = ~(U318 & U263 & U205); 
assign U280 = ~(U278 & STATO_REG_3__SCAN_IN); 
assign U284 = ~(U282 & STATO_REG_2__SCAN_IN); 
assign U324 = ~U255; 
assign U332 = ~(U274 & STATO_REG_1__SCAN_IN); 
assign U342 = ~(U274 & STATO_REG_0__SCAN_IN); 
assign U371 = ~(U330 & U255); 
assign U210 = ~(U332 & U218 & U341 & U340); 
assign U211 = ~(U283 & U218 & U284); 
assign U212 = ~(U280 & U279); 
assign U233 = ~(U343 & U342); 
assign U293 = ~U249; 
assign U305 = ~U250; 
assign U319 = ~U253; 
assign U353 = ~(U298 & U249); 
assign U363 = ~(U308 & U250); 
assign U367 = ~(U322 & U253); 
assign U370 = ~(U324 & VOTO0_REG_SCAN_IN); 
assign U243 = ~(U371 & U370); 
assign U352 = ~(U293 & VOTO1_REG_SCAN_IN); 
assign U362 = ~(U305 & VOTO3_REG_SCAN_IN); 
assign U366 = ~(U319 & VOTO2_REG_SCAN_IN); 
assign U238 = ~(U353 & U352); 
assign U239 = ~(U363 & U362); 
assign U241 = ~(U367 & U366); 
endmodule 
