module b11_C( X_IN_5_, X_IN_4_, X_IN_3_, X_IN_2_, X_IN_1_, X_IN_0_, STBI, STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, STATO_REG_2__SCAN_IN, STATO_REG_3__SCAN_IN, X_OUT_REG_0__SCAN_IN, X_OUT_REG_1__SCAN_IN, X_OUT_REG_2__SCAN_IN, X_OUT_REG_3__SCAN_IN, X_OUT_REG_4__SCAN_IN, X_OUT_REG_5__SCAN_IN, CONT1_REG_0__SCAN_IN, CONT1_REG_1__SCAN_IN, R_IN_REG_5__SCAN_IN, R_IN_REG_4__SCAN_IN, R_IN_REG_3__SCAN_IN, R_IN_REG_2__SCAN_IN, R_IN_REG_1__SCAN_IN, R_IN_REG_0__SCAN_IN, CONT_REG_5__SCAN_IN, CONT_REG_4__SCAN_IN, CONT_REG_3__SCAN_IN, CONT_REG_2__SCAN_IN, CONT_REG_1__SCAN_IN, CONT_REG_0__SCAN_IN, CONT1_REG_8__SCAN_IN, CONT1_REG_7__SCAN_IN, CONT1_REG_6__SCAN_IN, CONT1_REG_5__SCAN_IN, CONT1_REG_4__SCAN_IN, CONT1_REG_3__SCAN_IN, CONT1_REG_2__SCAN_IN, U360, U361, U362, U363, U364, U365, U366, U367, U368, U369, U370, U371, U372, U373, U374, U375, U376, U377, U378, U379, U380, U381, U382, U383, U384, U404, U405, U406, U407, U408, U409); 
input X_IN_5_, X_IN_4_, X_IN_3_, X_IN_2_, X_IN_1_, X_IN_0_, STBI, STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, STATO_REG_2__SCAN_IN, STATO_REG_3__SCAN_IN, X_OUT_REG_0__SCAN_IN, X_OUT_REG_1__SCAN_IN, X_OUT_REG_2__SCAN_IN, X_OUT_REG_3__SCAN_IN, X_OUT_REG_4__SCAN_IN, X_OUT_REG_5__SCAN_IN, CONT1_REG_0__SCAN_IN, CONT1_REG_1__SCAN_IN, R_IN_REG_5__SCAN_IN, R_IN_REG_4__SCAN_IN, R_IN_REG_3__SCAN_IN, R_IN_REG_2__SCAN_IN, R_IN_REG_1__SCAN_IN, R_IN_REG_0__SCAN_IN, CONT_REG_5__SCAN_IN, CONT_REG_4__SCAN_IN, CONT_REG_3__SCAN_IN, CONT_REG_2__SCAN_IN, CONT_REG_1__SCAN_IN, CONT_REG_0__SCAN_IN, CONT1_REG_8__SCAN_IN, CONT1_REG_7__SCAN_IN, CONT1_REG_6__SCAN_IN, CONT1_REG_5__SCAN_IN, CONT1_REG_4__SCAN_IN, CONT1_REG_3__SCAN_IN, CONT1_REG_2__SCAN_IN; 
output U360, U361, U362, U363, U364, U365, U366, U367, U368, U369, U370, U371, U372, U373, U374, U375, U376, U377, U378, U379, U380, U381, U382, U383, U384, U404, U405, U406, U407, U408, U409; 
wire U309, U310, U311, U312, U313, U314, U315, U316, U317, U318, U319, U320, U321, U322, U323, U324, U325, U326, U327, U328, U329, U330, U331, U332, U333, U334, U335, U336, U337, U338, U339, U340, U341, U342, U343, U344, U345, U346, U347, U348, U349, U350, U351, U352, U353, U354, U355, U356, U357, U358, U359, U385, U386, U387, U388, U389, U390, U391, U392, U393, U394, U395, U396, U397, U398, U399, U400, U401, U402, U403, U410, U411, U412, U413, U414, U415, U416, U417, U418, U419, U420, U421, U422, U423, U424, U425, U426, U427, U428, U429, U430, U431, U432, U433, U434, U435, U436, U437, U438, U439, U440, U441, U442, U443, U444, U445, U446, U447, U448, U449, U450, U451, U452, U453, U454, U455, U456, U457, U458, U459, U460, U461, U462, U463, U464, U465, U466, U467, U468, U469, U470, U471, U472, U473, U474, U475, U476, U477, U478, U479, U480, U481, U482, U483, U484, U485, U486, U487, U488, U489, U490, U491, U492, U493, U494, U495, U496, U497, U498, U499, U500, U501, U502, U503, U504, U505, U506, U507, U508, U509, U510, U511, U512, U513, U514, U515, U516, U517, U518, U519, U520, U521, U522, U523, U524, U525, U526, U527, U528, U529, U530, U531, U532, U533, U534, U535, U536, U537, U538, U539, U540, U541, U542, U543, U544, U545, U546, U547, U548, U549, U550, U551, U552, U553, U554, U555, U556, U557, U558, U559, U560, U561, U562, U563, U564, U565, U566, U567, U568, U569, U570, U571, U572, U573, U574, R229_U4, R229_U5, R229_U6, R229_U7, R229_U8, R229_U9, R229_U10, R229_U11, R229_U12, R229_U13, R229_U14, R229_U15, R229_U16, R229_U17, R229_U18, R229_U19, R229_U20, R229_U21, R229_U22, R229_U23, R229_U24, R229_U25, R229_U26, R229_U27, R229_U28, R229_U29, R229_U30, R229_U31, R229_U32, R229_U33, R229_U34, R229_U35, R229_U36, R229_U37, R229_U38, R229_U39, R229_U40, R229_U41, R229_U42, R229_U43, R229_U44, R229_U45, R229_U46, R229_U47, R229_U48, R229_U49, R229_U50, R229_U51, R229_U52, R229_U53, R229_U54, R229_U55, R229_U56, R229_U57, R229_U58, R229_U59, R229_U60, R229_U61, R229_U62, R229_U63, R229_U64, R229_U65, R229_U66, R229_U67, R229_U68, R229_U69, R229_U70, R229_U71, R229_U72, R229_U73, R229_U74, R229_U75, R229_U76, R229_U77, R229_U78, R229_U79, R229_U80, R229_U81, R229_U82, R229_U83, R229_U84, R229_U85, R229_U86, R229_U87, R229_U88, R229_U89, R229_U90, R229_U91, R229_U92, R229_U93, R229_U94, R229_U95, R229_U96, R229_U97, R229_U98, R229_U99, R229_U100, R229_U101, R229_U102, R229_U103, R229_U104, R229_U105, R229_U106, R229_U107, R229_U108, R229_U109, R229_U110, R229_U111, R229_U112, R229_U113, R229_U114, R229_U115, R229_U116, R229_U117, R229_U118, R229_U119, R229_U120, R229_U121, R229_U122, R229_U123, R229_U124, R229_U125, R229_U126, R229_U127, R229_U128, R248_U6, R248_U7, R248_U8, R248_U9, R248_U10, R248_U11, R248_U12, R248_U13, R248_U14, R248_U15, R248_U16, R248_U17, R248_U18, R248_U19, R248_U20, R248_U21, R248_U22, R248_U23, R248_U24, R248_U25, R248_U26, R248_U27, R248_U28, R248_U29, R248_U30, R248_U31, R248_U32, R248_U33, R248_U34, R248_U35, R248_U36, R248_U37, R248_U38, R248_U39, R248_U40, R248_U41, R248_U42, R248_U43, R248_U44, R248_U45, R248_U46, R248_U47, R248_U48, R248_U49, R248_U50, R248_U51, R248_U52, R248_U53, R248_U54, R248_U55, R248_U56, R248_U57, R248_U58, R248_U59, R248_U60, R248_U61, R248_U62, R248_U63, R248_U64, R248_U65, R248_U66, R248_U67, R248_U68, R248_U69, R248_U70, R248_U71, R248_U72, R248_U73, R248_U74, R248_U75, R248_U76, R248_U77, R248_U78, R248_U79, R248_U80, R248_U81, R248_U82, R248_U83, R248_U84, R248_U85, R248_U86, R248_U87, R248_U88, R248_U89, R248_U90, R248_U91, R248_U92, R248_U93, R248_U94, R248_U95, R248_U96, R248_U97, R248_U98, R248_U99, R248_U100, R248_U101, R248_U102, R248_U103, R248_U104, R248_U105, R248_U106, R248_U107, R248_U108, R248_U109, R248_U110, R248_U111, R248_U112, R248_U113, R248_U114, R248_U115, GT_80_U6, GT_80_U7, GT_80_U8, GT_80_U9, GT_80_U10, GT_87_U6, GT_87_U7, R259_U6, R259_U7, R259_U8, R259_U9, R259_U10, R259_U11, R259_U12, R259_U13, R259_U14, R259_U15, R259_U16, R259_U17, R259_U18, R259_U19, R259_U20, R259_U21, R259_U22, R259_U23, R259_U24, R259_U25, R259_U26, R259_U27, R259_U28, R259_U29, R259_U30, R259_U31, R259_U32, R259_U33, ADD_53_U5, ADD_53_U6, ADD_53_U7, ADD_53_U8, ADD_53_U9, ADD_53_U10, ADD_53_U11, ADD_53_U12, ADD_53_U13, ADD_53_U14, ADD_53_U15, ADD_53_U16, ADD_53_U17, ADD_53_U18, ADD_53_U19, ADD_53_U20, ADD_53_U21, ADD_53_U22, ADD_53_U23, ADD_53_U24, ADD_53_U25, ADD_53_U26, ADD_53_U27, ADD_53_U28, ADD_53_U29, ADD_53_U30, ADD_53_U31, ADD_53_U32, ADD_53_U33, ADD_88_U5, ADD_88_U6, ADD_88_U7, ADD_88_U8, ADD_88_U9, ADD_88_U10, ADD_88_U11, ADD_88_U12, ADD_88_U13, ADD_88_U14, ADD_88_U15, ADD_88_U16, ADD_88_U17, ADD_88_U18, ADD_88_U19, ADD_88_U20, ADD_88_U21, ADD_88_U22, ADD_88_U23, ADD_88_U24, ADD_88_U25, ADD_88_U26, ADD_88_U27, ADD_88_U28, ADD_88_U29, ADD_88_U30, ADD_88_U31, ADD_88_U32, ADD_88_U33, ADD_88_U34, ADD_88_U35, ADD_88_U36, ADD_88_U37, ADD_88_U38, ADD_88_U39, ADD_88_U40, ADD_88_U41, R254_U5, R254_U6, R254_U7, R254_U8, R254_U9, R254_U10, R254_U11, R254_U12, R254_U13, R254_U14, R254_U15, R254_U16, R254_U17, R254_U18, R254_U19, R254_U20, R254_U21, R254_U22, R254_U23, R254_U24, R254_U25, R254_U26, R254_U27, R254_U28, R254_U29, R254_U30, R254_U31, R254_U32, R254_U33, R254_U34, R254_U35, R254_U36, R254_U37, R254_U38, R254_U39, R254_U40, R254_U41, R254_U42, R254_U43, R254_U44, R254_U45, R254_U46, R254_U47, R254_U48, R254_U49, R254_U50, R254_U51, R254_U52, R254_U53, R254_U54, R254_U55, R254_U56, R254_U57, R254_U58, R254_U59, R254_U60, R254_U61, R254_U62, R254_U63, R254_U64, R254_U65, R254_U66, R254_U67, R254_U68, R254_U69, R254_U70, R254_U71, R254_U72, R254_U73, R254_U74, R254_U75, R254_U76, R254_U77, R254_U78, R254_U79, R254_U80, R254_U81, R254_U82, R254_U83, R254_U84, R254_U85, R254_U86, R254_U87, R254_U88, R254_U89, R254_U90, R254_U91, R254_U92, R254_U93, R254_U94, R254_U95, R254_U96, R254_U97, R254_U98, R254_U99, R254_U100, R254_U101, R254_U102, R254_U103, R254_U104, R254_U105, R254_U106, R254_U107, R254_U108, R254_U109, R254_U110, R254_U111, R254_U112, R254_U113, R254_U114, R254_U115, R254_U116, R254_U117, R254_U118, R254_U119, R254_U120, R254_U121, R254_U122, R254_U123, R254_U124, R254_U125, R254_U126, R254_U127, R254_U128; 
assign U310 = CONT1_REG_5__SCAN_IN & STATO_REG_3__SCAN_IN; 
assign U311 = CONT1_REG_2__SCAN_IN & STATO_REG_3__SCAN_IN; 
assign U312 = CONT1_REG_0__SCAN_IN & STATO_REG_3__SCAN_IN; 
assign U324 = STATO_REG_2__SCAN_IN & STATO_REG_1__SCAN_IN; 
assign U330 = ~(STATO_REG_2__SCAN_IN | STATO_REG_1__SCAN_IN); 
assign U331 = ~R_IN_REG_1__SCAN_IN; 
assign U358 = ~R_IN_REG_2__SCAN_IN; 
assign U359 = ~R_IN_REG_3__SCAN_IN; 
assign U386 = ~STATO_REG_1__SCAN_IN; 
assign U387 = ~STATO_REG_2__SCAN_IN; 
assign U388 = ~STATO_REG_0__SCAN_IN; 
assign U389 = ~R_IN_REG_5__SCAN_IN; 
assign U390 = ~R_IN_REG_4__SCAN_IN; 
assign U391 = ~R_IN_REG_0__SCAN_IN; 
assign U395 = ~CONT_REG_4__SCAN_IN; 
assign U396 = ~CONT_REG_3__SCAN_IN; 
assign U397 = ~CONT_REG_1__SCAN_IN; 
assign U399 = ~CONT1_REG_4__SCAN_IN; 
assign U400 = ~CONT1_REG_3__SCAN_IN; 
assign U401 = ~CONT1_REG_1__SCAN_IN; 
assign U402 = ~STATO_REG_3__SCAN_IN; 
assign U403 = ~CONT1_REG_8__SCAN_IN; 
assign U418 = ~STBI; 
assign U424 = ~(STATO_REG_1__SCAN_IN & STATO_REG_0__SCAN_IN); 
assign U452 = ~(STATO_REG_1__SCAN_IN & STATO_REG_0__SCAN_IN); 
assign U551 = STBI | STATO_REG_2__SCAN_IN; 
assign U552 = R_IN_REG_1__SCAN_IN | STATO_REG_0__SCAN_IN; 
assign R229_U5 = ~CONT1_REG_0__SCAN_IN; 
assign R229_U7 = ~CONT1_REG_1__SCAN_IN; 
assign R229_U8 = ~CONT1_REG_2__SCAN_IN; 
assign R229_U9 = ~CONT1_REG_3__SCAN_IN; 
assign R229_U10 = ~CONT1_REG_4__SCAN_IN; 
assign R229_U12 = ~CONT1_REG_5__SCAN_IN; 
assign R229_U14 = ~CONT1_REG_6__SCAN_IN; 
assign R229_U16 = ~CONT1_REG_7__SCAN_IN; 
assign R229_U31 = ~CONT1_REG_8__SCAN_IN; 
assign GT_80_U7 = CONT1_REG_1__SCAN_IN & CONT1_REG_0__SCAN_IN; 
assign GT_87_U7 = ~(CONT1_REG_7__SCAN_IN | CONT1_REG_6__SCAN_IN); 
assign ADD_53_U5 = ~CONT_REG_0__SCAN_IN; 
assign ADD_53_U6 = ~CONT_REG_1__SCAN_IN; 
assign ADD_53_U7 = ~(CONT_REG_1__SCAN_IN & CONT_REG_0__SCAN_IN); 
assign ADD_53_U8 = ~CONT_REG_2__SCAN_IN; 
assign ADD_53_U10 = ~CONT_REG_3__SCAN_IN; 
assign ADD_53_U12 = ~CONT_REG_4__SCAN_IN; 
assign ADD_53_U18 = ~CONT_REG_5__SCAN_IN; 
assign ADD_88_U5 = ~CONT1_REG_1__SCAN_IN; 
assign ADD_88_U8 = ~CONT1_REG_2__SCAN_IN; 
assign ADD_88_U10 = ~CONT1_REG_5__SCAN_IN; 
assign ADD_88_U12 = ~CONT1_REG_6__SCAN_IN; 
assign ADD_88_U14 = ~CONT1_REG_7__SCAN_IN; 
assign ADD_88_U15 = ~CONT1_REG_3__SCAN_IN; 
assign ADD_88_U21 = ~CONT1_REG_8__SCAN_IN; 
assign ADD_88_U23 = ~CONT1_REG_4__SCAN_IN; 
assign ADD_88_U24 = ~(CONT1_REG_2__SCAN_IN & CONT1_REG_1__SCAN_IN); 
assign ADD_88_U31 = ~(CONT1_REG_3__SCAN_IN & CONT1_REG_2__SCAN_IN & CONT1_REG_1__SCAN_IN); 
assign R254_U5 = ~R_IN_REG_0__SCAN_IN; 
assign R254_U6 = ~R_IN_REG_2__SCAN_IN; 
assign R254_U7 = ~R_IN_REG_3__SCAN_IN; 
assign R254_U8 = ~R_IN_REG_4__SCAN_IN; 
assign R254_U9 = ~R_IN_REG_5__SCAN_IN; 
assign R254_U22 = ~CONT1_REG_7__SCAN_IN; 
assign R254_U23 = ~CONT1_REG_0__SCAN_IN; 
assign R254_U24 = ~CONT1_REG_1__SCAN_IN; 
assign R254_U25 = ~CONT1_REG_2__SCAN_IN; 
assign R254_U26 = ~CONT1_REG_3__SCAN_IN; 
assign R254_U27 = ~CONT1_REG_4__SCAN_IN; 
assign R254_U28 = ~CONT1_REG_5__SCAN_IN; 
assign R254_U29 = ~CONT1_REG_6__SCAN_IN; 
assign R254_U30 = ~CONT1_REG_8__SCAN_IN; 
assign R254_U73 = ~(R_IN_REG_1__SCAN_IN & CONT1_REG_7__SCAN_IN); 
assign R254_U76 = ~(R_IN_REG_1__SCAN_IN & CONT1_REG_0__SCAN_IN); 
assign R254_U78 = ~(R_IN_REG_1__SCAN_IN & CONT1_REG_0__SCAN_IN); 
assign R254_U81 = ~(R_IN_REG_1__SCAN_IN & CONT1_REG_1__SCAN_IN); 
assign R254_U83 = ~(R_IN_REG_1__SCAN_IN & CONT1_REG_1__SCAN_IN); 
assign R254_U86 = ~(R_IN_REG_1__SCAN_IN & CONT1_REG_2__SCAN_IN); 
assign R254_U88 = ~(R_IN_REG_1__SCAN_IN & CONT1_REG_2__SCAN_IN); 
assign R254_U91 = ~(R_IN_REG_1__SCAN_IN & CONT1_REG_3__SCAN_IN); 
assign R254_U93 = ~(R_IN_REG_1__SCAN_IN & CONT1_REG_3__SCAN_IN); 
assign R254_U96 = ~(R_IN_REG_1__SCAN_IN & CONT1_REG_4__SCAN_IN); 
assign R254_U98 = ~(R_IN_REG_1__SCAN_IN & CONT1_REG_4__SCAN_IN); 
assign R254_U101 = ~(R_IN_REG_1__SCAN_IN & CONT1_REG_5__SCAN_IN); 
assign R254_U103 = ~(R_IN_REG_1__SCAN_IN & CONT1_REG_5__SCAN_IN); 
assign R254_U106 = ~(R_IN_REG_1__SCAN_IN & CONT1_REG_6__SCAN_IN); 
assign R254_U109 = ~(R_IN_REG_1__SCAN_IN & CONT1_REG_8__SCAN_IN); 
assign U325 = U387 & STATO_REG_1__SCAN_IN; 
assign U344 = U402 & CONT1_REG_8__SCAN_IN; 
assign U345 = U402 & CONT1_REG_7__SCAN_IN; 
assign U346 = U402 & CONT1_REG_6__SCAN_IN; 
assign U347 = U402 & CONT1_REG_5__SCAN_IN; 
assign U348 = U402 & CONT1_REG_4__SCAN_IN; 
assign U349 = U402 & CONT1_REG_3__SCAN_IN; 
assign U350 = U402 & CONT1_REG_2__SCAN_IN; 
assign U351 = U402 & CONT1_REG_1__SCAN_IN; 
assign U352 = U402 & CONT1_REG_0__SCAN_IN; 
assign U353 = ~(U399 & STATO_REG_3__SCAN_IN); 
assign U354 = ~(U400 & STATO_REG_3__SCAN_IN); 
assign U355 = ~(U401 & STATO_REG_3__SCAN_IN); 
assign U356 = ~(U359 & R_IN_REG_2__SCAN_IN); 
assign U393 = ~(U330 & U388); 
assign U417 = ~(U330 & U402); 
assign U422 = ~(U324 & STATO_REG_0__SCAN_IN); 
assign U425 = ~(U424 & STATO_REG_2__SCAN_IN); 
assign U427 = ~(U418 & U330 & STATO_REG_0__SCAN_IN); 
assign U433 = ~(U551 & U386 & U552); 
assign U548 = ~(U358 & R_IN_REG_3__SCAN_IN); 
assign U555 = ~(U331 & R_IN_REG_3__SCAN_IN); 
assign U556 = ~(U358 & R_IN_REG_1__SCAN_IN); 
assign U557 = ~(U389 & R_IN_REG_4__SCAN_IN); 
assign U558 = ~(U359 & R_IN_REG_5__SCAN_IN); 
assign U559 = ~(U390 & R_IN_REG_0__SCAN_IN); 
assign U560 = ~(U391 & R_IN_REG_2__SCAN_IN); 
assign U562 = ~(U386 & U388 & R_IN_REG_1__SCAN_IN); 
assign R229_U4 = ~U359; 
assign R229_U78 = ~(U359 & U358); 
assign R229_U84 = ~(U359 & R229_U31); 
assign R229_U89 = ~(U359 & R229_U16); 
assign R229_U94 = ~(U359 & R229_U14); 
assign R229_U124 = ~(U359 & R229_U5); 
assign R248_U7 = ~U312; 
assign R248_U11 = ~U311; 
assign R248_U18 = ~U310; 
assign GT_80_U10 = GT_80_U7 | CONT1_REG_2__SCAN_IN; 
assign GT_87_U6 = ~(GT_87_U7 | CONT1_REG_8__SCAN_IN); 
assign ADD_53_U20 = ~ADD_53_U7; 
assign ADD_53_U30 = ~(ADD_53_U7 & CONT_REG_2__SCAN_IN); 
assign ADD_53_U32 = ~(ADD_53_U5 & CONT_REG_1__SCAN_IN); 
assign ADD_53_U33 = ~(ADD_53_U6 & CONT_REG_0__SCAN_IN); 
assign ADD_88_U9 = ~(ADD_88_U15 & ADD_88_U24); 
assign ADD_88_U40 = ~(ADD_88_U8 & CONT1_REG_1__SCAN_IN); 
assign ADD_88_U41 = ~(ADD_88_U5 & CONT1_REG_2__SCAN_IN); 
assign R254_U72 = ~(U331 & R254_U22); 
assign R254_U75 = ~(U331 & R254_U23); 
assign R254_U77 = ~(U331 & R254_U23); 
assign R254_U80 = ~(U331 & R254_U24); 
assign R254_U82 = ~(U331 & R254_U24); 
assign R254_U85 = ~(U331 & R254_U25); 
assign R254_U87 = ~(U331 & R254_U25); 
assign R254_U90 = ~(U331 & R254_U26); 
assign R254_U92 = ~(U331 & R254_U26); 
assign R254_U95 = ~(U331 & R254_U27); 
assign R254_U97 = ~(U331 & R254_U27); 
assign R254_U100 = ~(U331 & R254_U28); 
assign R254_U102 = ~(U331 & R254_U28); 
assign R254_U105 = ~(U331 & R254_U29); 
assign R254_U108 = ~(U331 & R254_U30); 
assign U309 = U325 & U388; 
assign U357 = ~(U356 & U548); 
assign U410 = U560 & U559 & U558 & U557; 
assign U419 = ~GT_87_U6; 
assign U426 = ~(U325 & STATO_REG_0__SCAN_IN); 
assign U430 = ~U393; 
assign U434 = ~U417; 
assign U531 = ~(U393 & X_OUT_REG_5__SCAN_IN); 
assign U534 = ~(U393 & X_OUT_REG_4__SCAN_IN); 
assign U537 = ~(U393 & X_OUT_REG_3__SCAN_IN); 
assign U540 = ~(U393 & X_OUT_REG_2__SCAN_IN); 
assign U543 = ~(U393 & X_OUT_REG_1__SCAN_IN); 
assign U546 = ~(U393 & X_OUT_REG_0__SCAN_IN); 
assign U547 = ~U356; 
assign U563 = ~(U417 & R_IN_REG_5__SCAN_IN); 
assign U565 = ~(U417 & R_IN_REG_4__SCAN_IN); 
assign U567 = ~(U417 & R_IN_REG_3__SCAN_IN); 
assign U569 = ~(U417 & R_IN_REG_2__SCAN_IN); 
assign U571 = ~(U417 & R_IN_REG_1__SCAN_IN); 
assign U573 = ~(U417 & R_IN_REG_0__SCAN_IN); 
assign R229_U79 = ~(R229_U4 & R_IN_REG_2__SCAN_IN); 
assign R229_U81 = ~(U359 & U356); 
assign R229_U85 = ~(R229_U4 & CONT1_REG_8__SCAN_IN); 
assign R229_U90 = ~(R229_U4 & CONT1_REG_7__SCAN_IN); 
assign R229_U95 = ~(R229_U4 & CONT1_REG_6__SCAN_IN); 
assign R229_U125 = ~(R229_U4 & CONT1_REG_0__SCAN_IN); 
assign R248_U8 = ~U355; 
assign R248_U9 = ~U351; 
assign R248_U12 = ~U350; 
assign R248_U13 = ~U354; 
assign R248_U14 = ~U349; 
assign R248_U16 = ~U353; 
assign R248_U17 = ~U348; 
assign R248_U19 = ~U347; 
assign R248_U20 = ~U346; 
assign R248_U22 = ~U345; 
assign R248_U23 = ~U352; 
assign R248_U40 = ~U344; 
assign R248_U65 = ~(U347 & R248_U18); 
assign R248_U69 = ~(U346 & R248_U18); 
assign R248_U75 = ~(U352 & R248_U7); 
assign R248_U76 = ~(U344 & R248_U18); 
assign R248_U81 = ~(U345 & R248_U18); 
assign R248_U86 = ~(U346 & R248_U18); 
assign R248_U91 = ~(U347 & R248_U18); 
assign R248_U106 = ~(U350 & R248_U11); 
assign GT_80_U8 = GT_80_U10 & CONT1_REG_4__SCAN_IN & CONT1_REG_3__SCAN_IN; 
assign ADD_53_U9 = ~(ADD_53_U20 & CONT_REG_2__SCAN_IN); 
assign ADD_53_U17 = ~(ADD_53_U33 & ADD_53_U32); 
assign ADD_53_U31 = ~(ADD_53_U20 & ADD_53_U8); 
assign ADD_88_U7 = ~(ADD_88_U9 & ADD_88_U31); 
assign ADD_88_U20 = ~(ADD_88_U41 & ADD_88_U40); 
assign ADD_88_U25 = ~ADD_88_U9; 
assign ADD_88_U38 = ~(ADD_88_U9 & CONT1_REG_4__SCAN_IN); 
assign R254_U11 = ~(R254_U73 & R254_U72); 
assign R254_U12 = ~(R254_U106 & R254_U105); 
assign R254_U21 = ~(R254_U109 & R254_U108); 
assign R254_U41 = ~(R254_U76 & R254_U75 & R254_U5); 
assign R254_U45 = ~(R254_U81 & R254_U80 & U331); 
assign R254_U49 = ~(R254_U86 & R254_U85 & R254_U6); 
assign R254_U53 = ~(R254_U91 & R254_U90 & R254_U7); 
assign R254_U57 = ~(R254_U96 & R254_U95 & R254_U8); 
assign R254_U61 = ~(R254_U101 & R254_U100 & R254_U9); 
assign R254_U79 = ~(R254_U78 & R254_U77); 
assign R254_U84 = ~(R254_U83 & R254_U82); 
assign R254_U89 = ~(R254_U88 & R254_U87); 
assign R254_U94 = ~(R254_U93 & R254_U92); 
assign R254_U99 = ~(R254_U98 & R254_U97); 
assign R254_U104 = ~(R254_U103 & R254_U102); 
assign U316 = U430 & STATO_REG_3__SCAN_IN; 
assign U329 = U430 & U403; 
assign U361 = ~(U426 & U425); 
assign U385 = ~(U556 & U555 & U410); 
assign U431 = ~(U388 & U324 & U419); 
assign U435 = ~(U430 & U402); 
assign U549 = ~U357; 
assign U553 = ~(U419 & STATO_REG_1__SCAN_IN); 
assign U564 = ~(X_IN_5_ & U434); 
assign U566 = ~(X_IN_4_ & U434); 
assign U568 = ~(X_IN_3_ & U434); 
assign U570 = ~(X_IN_2_ & U434); 
assign U572 = ~(X_IN_1_ & U434); 
assign U574 = ~(X_IN_0_ & U434); 
assign R229_U18 = ~(R229_U79 & R229_U78); 
assign R229_U22 = ~(R229_U85 & R229_U84); 
assign R229_U23 = ~(R229_U90 & R229_U89); 
assign R229_U24 = ~(R229_U95 & R229_U94); 
assign R229_U30 = ~(R229_U125 & R229_U124); 
assign R229_U76 = ~(U357 & R229_U4); 
assign R229_U82 = ~(U547 & R229_U4); 
assign R248_U45 = ~(U312 & R248_U23); 
assign R248_U47 = ~(U355 & R248_U9); 
assign R248_U49 = ~(U351 & R248_U8); 
assign R248_U55 = ~(U354 & R248_U14); 
assign R248_U57 = ~(U349 & R248_U13); 
assign R248_U63 = ~(U310 & R248_U19); 
assign R248_U67 = ~(U310 & R248_U20); 
assign R248_U77 = ~(U310 & R248_U40); 
assign R248_U82 = ~(U310 & R248_U22); 
assign R248_U87 = ~(U310 & R248_U20); 
assign R248_U92 = ~(U310 & R248_U19); 
assign R248_U96 = ~(U348 & R248_U16); 
assign R248_U97 = ~(U353 & R248_U17); 
assign R248_U101 = ~(U349 & R248_U13); 
assign R248_U102 = ~(U354 & R248_U14); 
assign R248_U107 = ~(U311 & R248_U12); 
assign R248_U111 = ~(U351 & R248_U8); 
assign R248_U112 = ~(U355 & R248_U9); 
assign GT_80_U9 = ~(GT_80_U8 | CONT1_REG_7__SCAN_IN | CONT1_REG_6__SCAN_IN | CONT1_REG_5__SCAN_IN); 
assign ADD_53_U16 = ~(ADD_53_U31 & ADD_53_U30); 
assign ADD_53_U21 = ~ADD_53_U9; 
assign ADD_53_U28 = ~(ADD_53_U9 & CONT_REG_3__SCAN_IN); 
assign ADD_88_U26 = ~(ADD_88_U25 & ADD_88_U23); 
assign ADD_88_U30 = ~(ADD_88_U23 & ADD_88_U10 & ADD_88_U25); 
assign ADD_88_U39 = ~(ADD_88_U25 & ADD_88_U23); 
assign R254_U42 = ~(R254_U79 & R_IN_REG_0__SCAN_IN); 
assign R254_U43 = ~(U331 & R254_U41); 
assign R254_U46 = ~(R254_U84 & R_IN_REG_1__SCAN_IN); 
assign R254_U50 = ~(R254_U89 & R_IN_REG_2__SCAN_IN); 
assign R254_U54 = ~(R254_U94 & R_IN_REG_3__SCAN_IN); 
assign R254_U58 = ~(R254_U99 & R_IN_REG_4__SCAN_IN); 
assign R254_U62 = ~(R254_U104 & R_IN_REG_5__SCAN_IN); 
assign R254_U74 = ~R254_U11; 
assign R254_U107 = ~R254_U12; 
assign R254_U110 = ~R254_U21; 
assign U323 = U316 & CONT1_REG_8__SCAN_IN; 
assign U328 = U316 & U403; 
assign U332 = U385 & R_IN_REG_5__SCAN_IN; 
assign U333 = ~(U385 & U390); 
assign U334 = ~(U385 & U359); 
assign U335 = U385 & R_IN_REG_2__SCAN_IN; 
assign U336 = U385 & R_IN_REG_1__SCAN_IN; 
assign U337 = ~(U385 & U391); 
assign U404 = ~(U564 & U563); 
assign U405 = ~(U566 & U565); 
assign U406 = ~(U568 & U567); 
assign U407 = ~(U570 & U569); 
assign U408 = ~(U572 & U571); 
assign U409 = ~(U574 & U573); 
assign U421 = ~U385; 
assign U432 = ~(U309 & U385); 
assign U529 = ~(U310 & U329); 
assign U538 = ~(U311 & U329); 
assign U544 = ~(U312 & U329); 
assign R229_U19 = ~(R229_U82 & R229_U81); 
assign R229_U43 = ~(R229_U18 & R229_U5); 
assign R229_U57 = ~(R229_U18 & CONT1_REG_3__SCAN_IN); 
assign R229_U75 = ~(U359 & U549); 
assign R229_U80 = ~R229_U18; 
assign R229_U86 = ~R229_U22; 
assign R229_U91 = ~R229_U23; 
assign R229_U96 = ~R229_U24; 
assign R229_U110 = ~(R229_U18 & R229_U9); 
assign R229_U126 = ~R229_U30; 
assign R248_U6 = ~(R248_U45 & R248_U75); 
assign R248_U32 = ~(R248_U77 & R248_U76); 
assign R248_U33 = ~(R248_U82 & R248_U81); 
assign R248_U34 = ~(R248_U87 & R248_U86); 
assign R248_U35 = ~(R248_U92 & R248_U91); 
assign R248_U36 = ~(R248_U97 & R248_U96); 
assign R248_U37 = ~(R248_U102 & R248_U101); 
assign R248_U38 = ~(R248_U107 & R248_U106); 
assign R248_U39 = ~(R248_U112 & R248_U111); 
assign R248_U46 = ~R248_U45; 
assign R248_U48 = ~(R248_U47 & R248_U45); 
assign GT_80_U6 = ~(GT_80_U9 | CONT1_REG_8__SCAN_IN); 
assign ADD_53_U11 = ~(ADD_53_U21 & CONT_REG_3__SCAN_IN); 
assign ADD_53_U29 = ~(ADD_53_U21 & ADD_53_U10); 
assign ADD_88_U11 = ~(ADD_88_U26 & CONT1_REG_5__SCAN_IN); 
assign ADD_88_U19 = ~(ADD_88_U39 & ADD_88_U38); 
assign R254_U38 = ~(R254_U42 & R254_U43); 
assign R254_U39 = ~(R254_U41 & R254_U42); 
assign R254_U67 = ~(R254_U62 & R254_U61); 
assign R254_U68 = ~(R254_U58 & R254_U57); 
assign R254_U69 = ~(R254_U54 & R254_U53); 
assign R254_U70 = ~(R254_U50 & R254_U49); 
assign R254_U71 = ~(R254_U46 & R254_U45); 
assign U338 = U421 & CONT_REG_5__SCAN_IN; 
assign U339 = ~(U395 & U421); 
assign U340 = ~(U396 & U421); 
assign U341 = U421 & CONT_REG_2__SCAN_IN; 
assign U342 = ~(U397 & U421); 
assign U343 = U421 & CONT_REG_0__SCAN_IN; 
assign U363 = ~(U433 & U432 & U431 & U393); 
assign U420 = ~GT_80_U6; 
assign U423 = ~(U309 & U421); 
assign U436 = ~(U309 & U421); 
assign U450 = ~(U325 & U421); 
assign U532 = ~(U328 & CONT1_REG_4__SCAN_IN); 
assign U535 = ~(U328 & CONT1_REG_3__SCAN_IN); 
assign U541 = ~(U328 & CONT1_REG_1__SCAN_IN); 
assign U545 = ~(U323 & R248_U6); 
assign U550 = GT_80_U6 | STATO_REG_1__SCAN_IN; 
assign R229_U17 = ~(R229_U76 & R229_U75); 
assign R229_U44 = ~(U359 & R229_U43); 
assign R229_U45 = ~(R229_U80 & CONT1_REG_0__SCAN_IN); 
assign R229_U51 = ~(R229_U19 & R229_U8); 
assign R229_U55 = ~(R229_U80 & R229_U9); 
assign R229_U83 = ~R229_U19; 
assign R229_U100 = ~(R229_U19 & R229_U12); 
assign R229_U109 = ~(R229_U80 & CONT1_REG_3__SCAN_IN); 
assign R229_U115 = ~(R229_U19 & R229_U8); 
assign R229_U127 = ~(R229_U18 & R229_U126); 
assign R229_U128 = ~(R229_U30 & R229_U80); 
assign R248_U10 = ~(R248_U49 & R248_U48); 
assign R248_U78 = ~R248_U32; 
assign R248_U83 = ~R248_U33; 
assign R248_U88 = ~R248_U34; 
assign R248_U93 = ~R248_U35; 
assign R248_U98 = ~R248_U36; 
assign R248_U103 = ~R248_U37; 
assign R248_U108 = ~R248_U38; 
assign R248_U113 = ~R248_U39; 
assign R248_U115 = ~(R248_U39 & R248_U45); 
assign R259_U7 = ~U332; 
assign R259_U10 = ~U336; 
assign R259_U11 = ~U335; 
assign R259_U14 = ~U334; 
assign R259_U15 = ~U333; 
assign ADD_53_U15 = ~(ADD_53_U29 & ADD_53_U28); 
assign ADD_53_U22 = ~ADD_53_U11; 
assign ADD_53_U26 = ~(ADD_53_U11 & CONT_REG_4__SCAN_IN); 
assign ADD_88_U6 = ADD_88_U30 & ADD_88_U11; 
assign ADD_88_U27 = ~ADD_88_U11; 
assign ADD_88_U36 = ~(ADD_88_U11 & CONT1_REG_6__SCAN_IN); 
assign R254_U44 = ~R254_U38; 
assign R254_U47 = ~(R254_U45 & R254_U38); 
assign R254_U66 = ~R254_U39; 
assign R254_U125 = ~(R254_U71 & R254_U38); 
assign R254_U127 = ~(U331 & R254_U39); 
assign U360 = ~(U423 & U422); 
assign U364 = ~(U546 & U544 & U545); 
assign U394 = ~(U436 & U435); 
assign U554 = ~(U420 & STATO_REG_0__SCAN_IN); 
assign U561 = ~(U550 & STATO_REG_0__SCAN_IN); 
assign R229_U6 = ~(R229_U45 & R229_U44); 
assign R229_U27 = ~(R229_U110 & R229_U109); 
assign R229_U42 = R229_U128 & R229_U127; 
assign R229_U53 = ~(R229_U83 & CONT1_REG_2__SCAN_IN); 
assign R229_U59 = ~(R229_U17 & R229_U10); 
assign R229_U77 = ~R229_U17; 
assign R229_U99 = ~(R229_U83 & CONT1_REG_5__SCAN_IN); 
assign R229_U105 = ~(R229_U17 & R229_U10); 
assign R229_U114 = ~(R229_U83 & CONT1_REG_2__SCAN_IN); 
assign R229_U120 = ~(R229_U17 & R229_U7); 
assign R248_U50 = ~R248_U10; 
assign R248_U53 = ~(R248_U10 & R248_U11); 
assign R248_U110 = ~(R248_U38 & R248_U10); 
assign R248_U114 = ~(R248_U46 & R248_U113); 
assign R259_U8 = ~U339; 
assign R259_U9 = ~U342; 
assign R259_U12 = ~U341; 
assign R259_U13 = ~U340; 
assign R259_U16 = ~U338; 
assign R259_U17 = ~U343; 
assign R259_U19 = ~(U342 & R259_U10); 
assign R259_U24 = ~(U341 & R259_U11); 
assign R259_U25 = ~(U340 & R259_U14); 
assign R259_U30 = ~(U339 & R259_U15); 
assign R259_U33 = ~(U338 & R259_U7); 
assign ADD_53_U19 = ~(ADD_53_U22 & CONT_REG_4__SCAN_IN); 
assign ADD_53_U27 = ~(ADD_53_U22 & ADD_53_U12); 
assign ADD_88_U13 = ~(ADD_88_U27 & CONT1_REG_6__SCAN_IN); 
assign ADD_88_U37 = ~(ADD_88_U27 & ADD_88_U12); 
assign R254_U37 = ~(R254_U46 & R254_U47); 
assign R254_U126 = ~(R254_U46 & R254_U45 & R254_U44); 
assign R254_U128 = ~(R254_U66 & R_IN_REG_1__SCAN_IN); 
assign U428 = ~(U562 & U561 & STATO_REG_2__SCAN_IN); 
assign U437 = ~U394; 
assign U451 = ~(U553 & U554 & STATO_REG_2__SCAN_IN); 
assign R229_U25 = ~(R229_U100 & R229_U99); 
assign R229_U28 = ~(R229_U115 & R229_U114); 
assign R229_U46 = ~R229_U6; 
assign R229_U49 = ~(R229_U17 & R229_U6); 
assign R229_U61 = ~(R229_U77 & CONT1_REG_4__SCAN_IN); 
assign R229_U104 = ~(R229_U77 & CONT1_REG_4__SCAN_IN); 
assign R229_U111 = ~R229_U27; 
assign R229_U119 = ~(R229_U77 & CONT1_REG_1__SCAN_IN); 
assign R248_U31 = ~(R248_U115 & R248_U114); 
assign R248_U51 = ~(U311 & R248_U50); 
assign R248_U109 = ~(R248_U108 & R248_U50); 
assign R259_U18 = ~(U332 & R259_U16); 
assign R259_U20 = ~(U337 & R259_U17 & R259_U19); 
assign R259_U21 = ~(U336 & R259_U9); 
assign R259_U22 = ~(U335 & R259_U12); 
assign R259_U27 = ~(U334 & R259_U13); 
assign R259_U28 = ~(U333 & R259_U8); 
assign ADD_53_U14 = ~(ADD_53_U27 & ADD_53_U26); 
assign ADD_53_U23 = ~ADD_53_U19; 
assign ADD_53_U24 = ~(ADD_53_U19 & CONT_REG_5__SCAN_IN); 
assign ADD_88_U18 = ~(ADD_88_U37 & ADD_88_U36); 
assign ADD_88_U28 = ~ADD_88_U13; 
assign ADD_88_U34 = ~(ADD_88_U13 & CONT1_REG_7__SCAN_IN); 
assign R254_U15 = ~(R254_U128 & R254_U127); 
assign R254_U20 = ~(R254_U126 & R254_U125); 
assign R254_U48 = ~R254_U37; 
assign R254_U51 = ~(R254_U49 & R254_U37); 
assign R254_U123 = ~(R254_U70 & R254_U37); 
assign U398 = ~(U452 & U450 & U451); 
assign U439 = ~(U437 & CONT_REG_5__SCAN_IN); 
assign U441 = ~(U437 & CONT_REG_4__SCAN_IN); 
assign U443 = ~(U437 & CONT_REG_3__SCAN_IN); 
assign U445 = ~(U437 & CONT_REG_2__SCAN_IN); 
assign U447 = ~(U437 & CONT_REG_1__SCAN_IN); 
assign U449 = ~(U437 & CONT_REG_0__SCAN_IN); 
assign U542 = ~(U323 & R248_U31); 
assign R229_U26 = ~(R229_U105 & R229_U104); 
assign R229_U29 = ~(R229_U120 & R229_U119); 
assign R229_U47 = ~(R229_U46 & R229_U77); 
assign R229_U101 = ~R229_U25; 
assign R229_U116 = ~R229_U28; 
assign R248_U30 = ~(R248_U110 & R248_U109); 
assign R248_U52 = ~(U350 & R248_U51); 
assign R259_U23 = ~(R259_U21 & R259_U22 & R259_U20); 
assign ADD_53_U25 = ~(ADD_53_U23 & ADD_53_U18); 
assign ADD_88_U22 = ~(ADD_88_U28 & CONT1_REG_7__SCAN_IN); 
assign ADD_88_U35 = ~(ADD_88_U28 & ADD_88_U14); 
assign R254_U36 = ~(R254_U50 & R254_U51); 
assign R254_U124 = ~(R254_U50 & R254_U49 & R254_U48); 
assign U313 = U324 & U398; 
assign U315 = U398 & U386; 
assign U320 = U398 & U387; 
assign U365 = ~(U543 & U541 & U542); 
assign U453 = ~U398; 
assign U539 = ~(U323 & R248_U30); 
assign R229_U48 = ~(R229_U47 & CONT1_REG_1__SCAN_IN); 
assign R229_U106 = ~R229_U26; 
assign R229_U121 = ~R229_U29; 
assign R229_U123 = ~(R229_U29 & R229_U6); 
assign R248_U44 = ~(R248_U53 & R248_U52); 
assign R259_U26 = ~(R259_U24 & R259_U25 & R259_U23); 
assign ADD_53_U13 = ~(ADD_53_U25 & ADD_53_U24); 
assign ADD_88_U17 = ~(ADD_88_U35 & ADD_88_U34); 
assign ADD_88_U29 = ~ADD_88_U22; 
assign ADD_88_U32 = ~(ADD_88_U22 & CONT1_REG_8__SCAN_IN); 
assign R254_U19 = ~(R254_U124 & R254_U123); 
assign R254_U52 = ~R254_U36; 
assign R254_U55 = ~(R254_U53 & R254_U36); 
assign R254_U121 = ~(R254_U69 & R254_U36); 
assign U314 = U320 & STATO_REG_0__SCAN_IN; 
assign U318 = U313 & STATO_REG_0__SCAN_IN; 
assign U319 = U315 & STATO_REG_0__SCAN_IN; 
assign U326 = U313 & U388; 
assign U327 = U315 & U388; 
assign U366 = ~(U540 & U538 & U539); 
assign U458 = ~(U453 & CONT1_REG_8__SCAN_IN); 
assign U463 = ~(U453 & CONT1_REG_7__SCAN_IN); 
assign U469 = ~(U453 & CONT1_REG_6__SCAN_IN); 
assign U470 = ~(U320 & R_IN_REG_5__SCAN_IN); 
assign U472 = ~(ADD_88_U6 & U313); 
assign U479 = ~(U453 & CONT1_REG_5__SCAN_IN); 
assign U480 = ~(U320 & R_IN_REG_4__SCAN_IN); 
assign U482 = ~(ADD_88_U19 & U313); 
assign U489 = ~(U453 & CONT1_REG_4__SCAN_IN); 
assign U490 = ~(U320 & R_IN_REG_3__SCAN_IN); 
assign U492 = ~(ADD_88_U7 & U313); 
assign U499 = ~(U453 & CONT1_REG_3__SCAN_IN); 
assign U500 = ~(U320 & R_IN_REG_2__SCAN_IN); 
assign U501 = ~(R254_U19 & U315); 
assign U502 = ~(ADD_88_U20 & U313); 
assign U509 = ~(U453 & CONT1_REG_2__SCAN_IN); 
assign U510 = ~(U320 & R_IN_REG_1__SCAN_IN); 
assign U511 = ~(R254_U20 & U315); 
assign U512 = ~(ADD_88_U5 & U313); 
assign U519 = ~(U453 & CONT1_REG_1__SCAN_IN); 
assign U520 = ~(U320 & R_IN_REG_0__SCAN_IN); 
assign U521 = ~(R254_U15 & U315); 
assign U522 = ~(U313 & CONT1_REG_0__SCAN_IN); 
assign U528 = ~(U453 & CONT1_REG_0__SCAN_IN); 
assign R229_U40 = ~(R229_U49 & R229_U48); 
assign R229_U122 = ~(R229_U121 & R229_U46); 
assign R248_U54 = ~R248_U44; 
assign R248_U56 = ~(R248_U55 & R248_U44); 
assign R248_U105 = ~(R248_U37 & R248_U44); 
assign R259_U29 = ~(R259_U27 & R259_U28 & R259_U26); 
assign ADD_88_U33 = ~(ADD_88_U29 & ADD_88_U21); 
assign R254_U35 = ~(R254_U54 & R254_U55); 
assign R254_U122 = ~(R254_U54 & R254_U53 & R254_U52); 
assign U321 = U314 & R_IN_REG_0__SCAN_IN; 
assign U322 = U314 & U391; 
assign U460 = ~(ADD_88_U17 & U326); 
assign U465 = ~(ADD_88_U18 & U326); 
assign U503 = ~(U502 & U500 & U501); 
assign U506 = ~(R248_U30 & U319); 
assign U513 = ~(U511 & U510 & U512); 
assign U516 = ~(R248_U31 & U319); 
assign U523 = ~(U521 & U520 & U522); 
assign U525 = ~(R248_U6 & U319); 
assign U526 = ~(R229_U42 & U318); 
assign R229_U41 = R229_U123 & R229_U122; 
assign R229_U50 = ~R229_U40; 
assign R229_U52 = ~(R229_U51 & R229_U40); 
assign R229_U118 = ~(R229_U28 & R229_U40); 
assign R248_U15 = ~(R248_U57 & R248_U56); 
assign R248_U104 = ~(R248_U54 & R248_U103); 
assign R259_U31 = ~(R259_U29 & R259_U30); 
assign ADD_88_U16 = ~(ADD_88_U33 & ADD_88_U32); 
assign R254_U18 = ~(R254_U122 & R254_U121); 
assign R254_U56 = ~R254_U35; 
assign R254_U59 = ~(R254_U57 & R254_U35); 
assign R254_U119 = ~(R254_U68 & R254_U35); 
assign U455 = ~(ADD_88_U16 & U326); 
assign U466 = ~(U321 & CONT_REG_5__SCAN_IN); 
assign U474 = ~(U322 & CONT_REG_5__SCAN_IN); 
assign U475 = ~(U321 & CONT_REG_4__SCAN_IN); 
assign U484 = ~(U322 & CONT_REG_4__SCAN_IN); 
assign U485 = ~(U321 & CONT_REG_3__SCAN_IN); 
assign U491 = ~(R254_U18 & U315); 
assign U494 = ~(U322 & CONT_REG_3__SCAN_IN); 
assign U495 = ~(U321 & CONT_REG_2__SCAN_IN); 
assign U504 = ~(U322 & CONT_REG_2__SCAN_IN); 
assign U505 = ~(U321 & CONT_REG_1__SCAN_IN); 
assign U508 = ~(U503 & U388); 
assign U514 = ~(U322 & CONT_REG_1__SCAN_IN); 
assign U515 = ~(U321 & CONT_REG_0__SCAN_IN); 
assign U517 = ~(R229_U41 & U318); 
assign U518 = ~(U513 & U388); 
assign U524 = ~(U322 & CONT_REG_0__SCAN_IN); 
assign U527 = ~(U523 & U388); 
assign R229_U38 = ~(R229_U53 & R229_U52); 
assign R229_U117 = ~(R229_U50 & R229_U116); 
assign R248_U29 = ~(R248_U105 & R248_U104); 
assign R248_U58 = ~R248_U15; 
assign R248_U61 = ~(R248_U15 & R248_U16); 
assign R248_U100 = ~(R248_U36 & R248_U15); 
assign R259_U32 = ~(R259_U31 & R259_U18); 
assign R254_U34 = ~(R254_U58 & R254_U59); 
assign R254_U120 = ~(R254_U58 & R254_U57 & R254_U56); 
assign U370 = ~(U525 & U526 & U524 & U528 & U527); 
assign U416 = U519 & U517; 
assign U493 = ~(U492 & U490 & U491); 
assign U496 = ~(R248_U29 & U319); 
assign U536 = ~(U323 & R248_U29); 
assign R229_U21 = ~(R229_U118 & R229_U117); 
assign R229_U54 = ~R229_U38; 
assign R229_U56 = ~(R229_U55 & R229_U38); 
assign R229_U113 = ~(R229_U27 & R229_U38); 
assign R248_U59 = ~(U353 & R248_U58); 
assign R248_U99 = ~(R248_U98 & R248_U58); 
assign R259_U6 = ~(R259_U33 & R259_U32); 
assign R254_U17 = ~(R254_U120 & R254_U119); 
assign R254_U60 = ~R254_U34; 
assign R254_U63 = ~(R254_U61 & R254_U34); 
assign R254_U117 = ~(R254_U67 & R254_U34); 
assign U367 = ~(U537 & U535 & U536); 
assign U371 = ~(U515 & U514 & U516 & U416 & U518); 
assign U392 = ~R259_U6; 
assign U429 = ~(U309 & U385 & R259_U6); 
assign U481 = ~(R254_U17 & U315); 
assign U498 = ~(U493 & U388); 
assign U507 = ~(R229_U21 & U318); 
assign R229_U37 = ~(R229_U57 & R229_U56); 
assign R229_U112 = ~(R229_U54 & R229_U111); 
assign R248_U28 = ~(R248_U100 & R248_U99); 
assign R248_U60 = ~(U348 & R248_U59); 
assign R254_U32 = ~(R254_U62 & R254_U63); 
assign R254_U118 = ~(R254_U62 & R254_U61 & R254_U60); 
assign U317 = U394 & U392 & STATO_REG_1__SCAN_IN; 
assign U362 = ~(U428 & U427 & U429); 
assign U415 = U509 & U507; 
assign U483 = ~(U482 & U480 & U481); 
assign U486 = ~(R248_U28 & U319); 
assign U533 = ~(U323 & R248_U28); 
assign R229_U39 = R229_U113 & R229_U112; 
assign R229_U58 = ~R229_U37; 
assign R229_U60 = ~(R229_U59 & R229_U37); 
assign R229_U108 = ~(R229_U26 & R229_U37); 
assign R248_U43 = ~(R248_U61 & R248_U60); 
assign R254_U10 = ~(R254_U12 & R254_U32); 
assign R254_U16 = ~(R254_U118 & R254_U117); 
assign R254_U64 = ~R254_U32; 
assign R254_U116 = ~(R254_U12 & R254_U32); 
assign U368 = ~(U534 & U532 & U533); 
assign U372 = ~(U505 & U504 & U506 & U415 & U508); 
assign U438 = ~(ADD_53_U13 & U317); 
assign U440 = ~(ADD_53_U14 & U317); 
assign U442 = ~(ADD_53_U15 & U317); 
assign U444 = ~(ADD_53_U16 & U317); 
assign U446 = ~(ADD_53_U17 & U317); 
assign U448 = ~(ADD_53_U5 & U317); 
assign U471 = ~(R254_U16 & U315); 
assign U488 = ~(U483 & U388); 
assign U497 = ~(R229_U39 & U318); 
assign R229_U11 = ~(R229_U61 & R229_U60); 
assign R229_U107 = ~(R229_U58 & R229_U106); 
assign R248_U62 = ~R248_U43; 
assign R248_U64 = ~(R248_U63 & R248_U43); 
assign R248_U95 = ~(R248_U35 & R248_U43); 
assign R254_U40 = ~R254_U10; 
assign R254_U114 = ~(R254_U11 & R254_U10); 
assign R254_U115 = ~(R254_U64 & R254_U107); 
assign U379 = ~(U449 & U448); 
assign U380 = ~(U447 & U446); 
assign U381 = ~(U445 & U444); 
assign U382 = ~(U443 & U442); 
assign U383 = ~(U441 & U440); 
assign U384 = ~(U439 & U438); 
assign U414 = U499 & U497; 
assign U473 = ~(U472 & U470 & U471); 
assign R229_U20 = ~(R229_U108 & R229_U107); 
assign R229_U62 = ~R229_U11; 
assign R229_U65 = ~(R229_U11 & CONT1_REG_5__SCAN_IN); 
assign R229_U103 = ~(R229_U25 & R229_U11); 
assign R248_U42 = ~(R248_U65 & R248_U64); 
assign R248_U94 = ~(R248_U62 & R248_U93); 
assign R254_U31 = ~(R254_U40 & R254_U11); 
assign R254_U33 = R254_U116 & R254_U115; 
assign R254_U113 = ~(R254_U74 & R254_U40); 
assign U373 = ~(U495 & U494 & U496 & U414 & U498); 
assign U464 = ~(R254_U33 & U327); 
assign U478 = ~(U473 & U388); 
assign U487 = ~(R229_U20 & U318); 
assign R229_U63 = ~(R229_U62 & R229_U12); 
assign R229_U102 = ~(R229_U101 & R229_U62); 
assign R248_U27 = ~(R248_U95 & R248_U94); 
assign R248_U66 = ~R248_U42; 
assign R248_U68 = ~(R248_U67 & R248_U42); 
assign R248_U90 = ~(R248_U34 & R248_U42); 
assign R254_U14 = ~(R254_U114 & R254_U113); 
assign R254_U65 = ~R254_U31; 
assign R254_U112 = ~(R254_U21 & R254_U31); 
assign U413 = U489 & U487; 
assign U459 = ~(R254_U14 & U327); 
assign U476 = ~(R248_U27 & U319); 
assign U530 = ~(U323 & R248_U27); 
assign R229_U36 = R229_U103 & R229_U102; 
assign R229_U64 = ~(R229_U19 & R229_U63); 
assign R248_U21 = ~(R248_U69 & R248_U68); 
assign R248_U89 = ~(R248_U66 & R248_U88); 
assign R254_U111 = ~(R254_U65 & R254_U110); 
assign U369 = ~(U531 & U529 & U530); 
assign U374 = ~(U485 & U484 & U486 & U413 & U488); 
assign U477 = ~(R229_U36 & U318); 
assign R229_U13 = ~(R229_U65 & R229_U64); 
assign R248_U26 = ~(R248_U90 & R248_U89); 
assign R248_U70 = ~R248_U21; 
assign R248_U73 = ~(R248_U21 & R248_U18); 
assign R248_U85 = ~(R248_U33 & R248_U21); 
assign R254_U13 = ~(R254_U112 & R254_U111); 
assign U412 = U479 & U477; 
assign U454 = ~(R254_U13 & U327); 
assign U467 = ~(R248_U26 & U319); 
assign R229_U66 = ~R229_U13; 
assign R229_U69 = ~(R229_U13 & CONT1_REG_6__SCAN_IN); 
assign R229_U98 = ~(R229_U24 & R229_U13); 
assign R248_U71 = ~(R248_U70 & U310); 
assign R248_U84 = ~(R248_U83 & R248_U70); 
assign U375 = ~(U475 & U474 & U476 & U412 & U478); 
assign R229_U67 = ~(R229_U66 & R229_U14); 
assign R229_U97 = ~(R229_U96 & R229_U66); 
assign R248_U25 = ~(R248_U85 & R248_U84); 
assign R248_U72 = ~(U345 & R248_U71); 
assign U461 = ~(R248_U25 & U319); 
assign R229_U35 = R229_U98 & R229_U97; 
assign R229_U68 = ~(U359 & R229_U67); 
assign R248_U41 = ~(R248_U73 & R248_U72); 
assign U468 = ~(R229_U35 & U318); 
assign R229_U15 = ~(R229_U69 & R229_U68); 
assign R248_U74 = ~R248_U41; 
assign R248_U80 = ~(R248_U32 & R248_U41); 
assign U411 = U469 & U467 & U468; 
assign R229_U70 = ~R229_U15; 
assign R229_U73 = ~(R229_U15 & CONT1_REG_7__SCAN_IN); 
assign R229_U93 = ~(R229_U23 & R229_U15); 
assign R248_U79 = ~(R248_U74 & R248_U78); 
assign U376 = ~(U465 & U466 & U464 & U411); 
assign R229_U71 = ~(R229_U70 & R229_U16); 
assign R229_U92 = ~(R229_U91 & R229_U70); 
assign R248_U24 = ~(R248_U80 & R248_U79); 
assign U456 = ~(R248_U24 & U319); 
assign R229_U34 = R229_U93 & R229_U92; 
assign R229_U72 = ~(U359 & R229_U71); 
assign U462 = ~(R229_U34 & U318); 
assign R229_U32 = ~(R229_U73 & R229_U72); 
assign U377 = ~(U460 & U461 & U463 & U459 & U462); 
assign R229_U74 = ~R229_U32; 
assign R229_U88 = ~(R229_U22 & R229_U32); 
assign R229_U87 = ~(R229_U74 & R229_U86); 
assign R229_U33 = R229_U88 & R229_U87; 
assign U457 = ~(R229_U33 & U318); 
assign U378 = ~(U455 & U456 & U458 & U454 & U457); 
endmodule 
