module b04_C( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_, DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_, STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN, DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN, DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN, DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN, DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN, REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN, RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN, RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN, RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN, RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN, RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN, RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN, RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN, RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN, REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN, REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN, REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U281, U282, U283, U284, U285, U286, U287, U288, U289, U290, U291, U292, U293, U294, U295, U296, U297, U298, U299, U300, U301, U302, U303, U304, U305, U306, U307, U308, U309, U310, U311, U312, U313, U314, U315, U316, U317, U318, U319, U320, U321, U322, U323, U324, U325, U326, U327, U328, U329, U330, U331, U332, U333, U334, U335, U336, U337, U338, U339, U340, U341, U342, U343, U344, U375); 
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_, DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_, STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN, DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN, DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN, DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN, DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN, REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN, RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN, RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN, RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN, RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN, RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN, RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN, RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN, RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN, REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN, REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN, REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN; 
output U281, U282, U283, U284, U285, U286, U287, U288, U289, U290, U291, U292, U293, U294, U295, U296, U297, U298, U299, U300, U301, U302, U303, U304, U305, U306, U307, U308, U309, U310, U311, U312, U313, U314, U315, U316, U317, U318, U319, U320, U321, U322, U323, U324, U325, U326, U327, U328, U329, U330, U331, U332, U333, U334, U335, U336, U337, U338, U339, U340, U341, U342, U343, U344, U375; 
wire U272, U273, U274, U275, U276, U277, U278, U279, U280, U345, U346, U347, U348, U349, U350, U351, U352, U353, U354, U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U365, U366, U367, U368, U369, U370, U371, U372, U373, U374, U376, U377, U378, U379, U380, U381, U382, U383, U384, U385, U386, U387, U388, U389, U390, U391, U392, U393, U394, U395, U396, U397, U398, U399, U400, U401, U402, U403, U404, U405, U406, U407, U408, U409, U410, U411, U412, U413, U414, U415, U416, U417, U418, U419, U420, U421, U422, U423, U424, U425, U426, U427, U428, U429, U430, U431, U432, U433, U434, U435, U436, U437, U438, U439, U440, U441, U442, U443, U444, U445, U446, U447, U448, U449, U450, U451, U452, U453, U454, U455, U456, U457, U458, U459, U460, U461, U462, U463, U464, U465, U466, U467, U468, U469, U470, U471, U472, U473, U474, U475, U476, U477, U478, U479, U480, U481, U482, U483, U484, U485, U486, U487, U488, U489, U490, U491, U492, U493, U494, U495, U496, U497, U498, U499, U500, U501, U502, U503, U504, U505, U506, U507, U508, U509, U510, U511, U512, U513, U514, U515, U516, U517, U518, U519, U520, U521, U522, U523, U524, U525, U526, U527, U528, U529, U530, U531, U532, U533, U534, U535, U536, U537, U538, U539, U540, U541, U542, U543, U544, U545, U546, U547, U548, U549, U550, U551, U552, U553, U554, U555, U556, U557, U558, U559, U560, U561, U562, U563, U564, U565, U566, U567, U568, U569, U570, U571, U572, U573, U574, U575, U576, U577, U578, GTE_67_U6, SUB_82_U6, SUB_82_U7, SUB_82_U8, SUB_82_U9, SUB_82_U10, SUB_82_U11, SUB_82_U12, SUB_82_U13, SUB_82_U14, SUB_82_U15, SUB_82_U16, SUB_82_U17, SUB_82_U18, SUB_82_U19, SUB_82_U20, SUB_82_U21, SUB_82_U22, SUB_82_U23, SUB_82_U24, SUB_82_U25, SUB_82_U26, SUB_82_U27, SUB_82_U28, SUB_82_U29, SUB_82_U30, SUB_82_U31, SUB_82_U32, SUB_82_U33, SUB_82_U34, SUB_82_U35, ADD_65_U4, ADD_65_U5, ADD_65_U6, ADD_65_U7, ADD_65_U8, ADD_65_U9, ADD_65_U10, ADD_65_U11, ADD_65_U12, ADD_65_U13, ADD_65_U14, ADD_65_U15, ADD_65_U16, ADD_65_U17, ADD_65_U18, ADD_65_U19, ADD_65_U20, ADD_65_U21, ADD_65_U22, ADD_65_U23, ADD_65_U24, ADD_65_U25, ADD_65_U26, ADD_65_U27, ADD_65_U28, ADD_65_U29, ADD_65_U30, ADD_65_U31, ADD_77_U4, ADD_77_U5, ADD_77_U6, ADD_77_U7, ADD_77_U8, ADD_77_U9, ADD_77_U10, ADD_77_U11, ADD_77_U12, ADD_77_U13, ADD_77_U14, ADD_77_U15, ADD_77_U16, ADD_77_U17, ADD_77_U18, ADD_77_U19, ADD_77_U20, ADD_77_U21, ADD_77_U22, ADD_77_U23, ADD_77_U24, ADD_77_U25, ADD_77_U26, ADD_77_U27, ADD_77_U28, ADD_77_U29, ADD_77_U30, ADD_77_U31, SUB_70_166_U6, SUB_70_166_U7, SUB_70_166_U8, SUB_70_166_U9, SUB_70_166_U10, SUB_70_166_U11, SUB_70_166_U12, SUB_70_166_U13, SUB_70_166_U14, SUB_70_166_U15, SUB_70_166_U16, SUB_70_166_U17, SUB_70_166_U18, SUB_70_166_U19, SUB_70_166_U20, SUB_70_166_U21, SUB_70_166_U22, SUB_70_166_U23, SUB_70_166_U24, SUB_70_166_U25, SUB_70_166_U26, SUB_70_166_U27, SUB_70_166_U28, SUB_70_166_U29, SUB_70_166_U30, SUB_70_166_U31, SUB_70_166_U32, SUB_70_166_U33, SUB_70_166_U34, SUB_70_166_U35, LT_90_U6, LT_90_U7, LT_90_U8, LT_90_U9, LT_90_U10, LT_90_U11, LT_90_U12, LT_90_U13, LT_90_U14, LT_90_U15, LT_90_U16, LT_90_U17, LT_90_U18, LT_90_U19, LT_90_U20, LT_90_U21, LT_90_U22, LT_90_U23, LT_90_U24, LT_90_U25, LT_90_U26, LT_90_U27, LT_90_U28, LT_90_U29, LT_90_U30, LT_90_U31, LT_90_U32, LT_90_U33, LT_90_U34, LT_90_U35, LT_90_U36, LT_90_U37, LT_90_U38, LT_90_U39, LT_90_U40, LT_90_U41, LT_90_U42, GT_88_U6, GT_88_U7, GT_88_U8, GT_88_U9, GT_88_U10, GT_88_U11, GT_88_U12, GT_88_U13, GT_88_U14, GT_88_U15, GT_88_U16, GT_88_U17, GT_88_U18, GT_88_U19, GT_88_U20, GT_88_U21, GT_88_U22, GT_88_U23, GT_88_U24, GT_88_U25, GT_88_U26, GT_88_U27, GT_88_U28, GT_88_U29, GT_88_U30, GT_88_U31, GT_88_U32, GT_88_U33, GT_88_U34, GT_88_U35, GT_88_U36, GT_88_U37, GT_88_U38, GT_88_U39, GT_88_U40, GT_88_U41, GT_88_U42, SUB_82_165_U6, SUB_82_165_U7, SUB_82_165_U8, SUB_82_165_U9, SUB_82_165_U10, SUB_82_165_U11, SUB_82_165_U12, SUB_82_165_U13, SUB_82_165_U14, SUB_82_165_U15, SUB_82_165_U16, SUB_82_165_U17, SUB_82_165_U18, SUB_82_165_U19, SUB_82_165_U20, SUB_82_165_U21, SUB_82_165_U22, SUB_82_165_U23, SUB_82_165_U24, SUB_82_165_U25, SUB_82_165_U26, SUB_82_165_U27, SUB_82_165_U28, SUB_82_165_U29, SUB_82_165_U30, SUB_82_165_U31, SUB_82_165_U32, SUB_82_165_U33, SUB_82_165_U34, SUB_82_165_U35, GTE_79_U6, R179_U4, R179_U5, R179_U6, R179_U7, R179_U8, R179_U9, R179_U10, R179_U11, R179_U12, R179_U13, R179_U14, R179_U15, R179_U16, R179_U17, R179_U18, R179_U19, R179_U20, R179_U21, R179_U22, R179_U23, R179_U24, R179_U25, R179_U26, R179_U27, R179_U28, R179_U29, R179_U30, R179_U31, R179_U32, R179_U33, R179_U34, R179_U35, R179_U36, R179_U37, R179_U38, R179_U39, R179_U40, R179_U41, R179_U42, R179_U43, R179_U44, R179_U45, R179_U46, R179_U47, R179_U48, R179_U49, R179_U50, R179_U51, R179_U52, R179_U53, R179_U54, R179_U55, R179_U56, R179_U57, R179_U58, R179_U59, R179_U60, R179_U61, R179_U62, R179_U63, R179_U64, R179_U65, R179_U66, R179_U67, R179_U68, R179_U69, R179_U70, R179_U71, R179_U72, R179_U73, R179_U74, R179_U75, R179_U76, R179_U77, R179_U78, R179_U79, R179_U80, R179_U81, R179_U82, R179_U83, R179_U84, R179_U85, R179_U86, R179_U87, R179_U88, R179_U89, R179_U90, R179_U91, R179_U92, R179_U93, R179_U94, R179_U95, R179_U96, SUB_70_U6, SUB_70_U7, SUB_70_U8, SUB_70_U9, SUB_70_U10, SUB_70_U11, SUB_70_U12, SUB_70_U13, SUB_70_U14, SUB_70_U15, SUB_70_U16, SUB_70_U17, SUB_70_U18, SUB_70_U19, SUB_70_U20, SUB_70_U21, SUB_70_U22, SUB_70_U23, SUB_70_U24, SUB_70_U25, SUB_70_U26, SUB_70_U27, SUB_70_U28, SUB_70_U29, SUB_70_U30, SUB_70_U31, SUB_70_U32, SUB_70_U33, SUB_70_U34, SUB_70_U35; 
assign U345 = ~STATO_REG_0__SCAN_IN; 
assign U346 = ~STATO_REG_1__SCAN_IN; 
assign U349 = ~AVERAGE; 
assign U350 = ~ENABLE; 
assign U351 = ~RESTART; 
assign U374 = STATO_REG_1__SCAN_IN | STATO_REG_0__SCAN_IN; 
assign U420 = ENABLE | STATO_REG_0__SCAN_IN; 
assign U552 = ~(RESTART & RMAX_REG_6__SCAN_IN); 
assign U554 = ~(RESTART & RMAX_REG_5__SCAN_IN); 
assign U556 = ~(RESTART & RMAX_REG_4__SCAN_IN); 
assign U558 = ~(RESTART & RMAX_REG_3__SCAN_IN); 
assign U560 = ~(RESTART & RMAX_REG_2__SCAN_IN); 
assign U562 = ~(RESTART & RMAX_REG_1__SCAN_IN); 
assign U564 = ~(RESTART & RMAX_REG_0__SCAN_IN); 
assign U566 = ~(RESTART & RMIN_REG_6__SCAN_IN); 
assign U568 = ~(RESTART & RMIN_REG_5__SCAN_IN); 
assign U570 = ~(RESTART & RMIN_REG_4__SCAN_IN); 
assign U572 = ~(RESTART & RMIN_REG_3__SCAN_IN); 
assign U574 = ~(RESTART & RMIN_REG_2__SCAN_IN); 
assign U576 = ~(RESTART & RMIN_REG_1__SCAN_IN); 
assign U578 = ~(RESTART & RMIN_REG_0__SCAN_IN); 
assign ADD_65_U6 = ~RMAX_REG_6__SCAN_IN; 
assign ADD_65_U8 = RMAX_REG_5__SCAN_IN | RMIN_REG_5__SCAN_IN; 
assign ADD_65_U9 = ~(RMAX_REG_1__SCAN_IN & RMIN_REG_1__SCAN_IN); 
assign ADD_65_U10 = ~(RMAX_REG_0__SCAN_IN & RMIN_REG_0__SCAN_IN); 
assign ADD_65_U12 = RMAX_REG_1__SCAN_IN | RMIN_REG_1__SCAN_IN; 
assign ADD_65_U13 = RMAX_REG_2__SCAN_IN | RMIN_REG_2__SCAN_IN; 
assign ADD_65_U15 = ~(RMAX_REG_3__SCAN_IN & RMIN_REG_3__SCAN_IN); 
assign ADD_65_U16 = ~(RMAX_REG_2__SCAN_IN & RMIN_REG_2__SCAN_IN); 
assign ADD_65_U18 = RMAX_REG_3__SCAN_IN | RMIN_REG_3__SCAN_IN; 
assign ADD_65_U19 = RMAX_REG_4__SCAN_IN | RMIN_REG_4__SCAN_IN; 
assign ADD_65_U21 = ~(RMAX_REG_4__SCAN_IN & RMIN_REG_4__SCAN_IN); 
assign ADD_65_U24 = ~(RMAX_REG_5__SCAN_IN & RMIN_REG_5__SCAN_IN); 
assign ADD_65_U29 = RMAX_REG_7__SCAN_IN | RMIN_REG_7__SCAN_IN; 
assign ADD_65_U30 = ~(RMAX_REG_7__SCAN_IN & RMIN_REG_7__SCAN_IN); 
assign ADD_77_U6 = ~DATA_IN_6_; 
assign ADD_77_U8 = DATA_IN_5_ | REG4_REG_5__SCAN_IN; 
assign ADD_77_U9 = ~(DATA_IN_1_ & REG4_REG_1__SCAN_IN); 
assign ADD_77_U10 = ~(DATA_IN_0_ & REG4_REG_0__SCAN_IN); 
assign ADD_77_U12 = DATA_IN_1_ | REG4_REG_1__SCAN_IN; 
assign ADD_77_U13 = DATA_IN_2_ | REG4_REG_2__SCAN_IN; 
assign ADD_77_U15 = ~(DATA_IN_3_ & REG4_REG_3__SCAN_IN); 
assign ADD_77_U16 = ~(DATA_IN_2_ & REG4_REG_2__SCAN_IN); 
assign ADD_77_U18 = DATA_IN_3_ | REG4_REG_3__SCAN_IN; 
assign ADD_77_U19 = DATA_IN_4_ | REG4_REG_4__SCAN_IN; 
assign ADD_77_U21 = ~(DATA_IN_4_ & REG4_REG_4__SCAN_IN); 
assign ADD_77_U24 = ~(DATA_IN_5_ & REG4_REG_5__SCAN_IN); 
assign ADD_77_U29 = DATA_IN_7_ | REG4_REG_7__SCAN_IN; 
assign ADD_77_U30 = ~(DATA_IN_7_ & REG4_REG_7__SCAN_IN); 
assign LT_90_U7 = ~DATA_IN_7_; 
assign LT_90_U8 = ~DATA_IN_1_; 
assign LT_90_U9 = ~RMIN_REG_1__SCAN_IN; 
assign LT_90_U10 = ~RMIN_REG_2__SCAN_IN; 
assign LT_90_U11 = ~DATA_IN_2_; 
assign LT_90_U12 = ~DATA_IN_3_; 
assign LT_90_U13 = ~RMIN_REG_3__SCAN_IN; 
assign LT_90_U14 = ~RMIN_REG_4__SCAN_IN; 
assign LT_90_U15 = ~DATA_IN_4_; 
assign LT_90_U16 = ~DATA_IN_5_; 
assign LT_90_U17 = ~RMIN_REG_5__SCAN_IN; 
assign LT_90_U18 = ~RMIN_REG_6__SCAN_IN; 
assign LT_90_U19 = ~DATA_IN_6_; 
assign LT_90_U20 = ~RMIN_REG_7__SCAN_IN; 
assign LT_90_U21 = ~DATA_IN_0_; 
assign GT_88_U7 = ~RMAX_REG_7__SCAN_IN; 
assign GT_88_U8 = ~RMAX_REG_1__SCAN_IN; 
assign GT_88_U9 = ~DATA_IN_1_; 
assign GT_88_U10 = ~DATA_IN_2_; 
assign GT_88_U11 = ~RMAX_REG_2__SCAN_IN; 
assign GT_88_U12 = ~RMAX_REG_3__SCAN_IN; 
assign GT_88_U13 = ~DATA_IN_3_; 
assign GT_88_U14 = ~DATA_IN_4_; 
assign GT_88_U15 = ~RMAX_REG_4__SCAN_IN; 
assign GT_88_U16 = ~RMAX_REG_5__SCAN_IN; 
assign GT_88_U17 = ~DATA_IN_5_; 
assign GT_88_U18 = ~DATA_IN_6_; 
assign GT_88_U19 = ~RMAX_REG_6__SCAN_IN; 
assign GT_88_U20 = ~DATA_IN_7_; 
assign GT_88_U21 = ~RMAX_REG_0__SCAN_IN; 
assign U278 = U420 & STATO_REG_1__SCAN_IN; 
assign U348 = ~(U345 & STATO_REG_1__SCAN_IN); 
assign U375 = ~U374; 
assign U377 = ~(U346 & STATO_REG_0__SCAN_IN); 
assign U421 = ~(U374 & U420); 
assign U551 = ~(DATA_IN_6_ & U351); 
assign U553 = ~(DATA_IN_5_ & U351); 
assign U555 = ~(DATA_IN_4_ & U351); 
assign U557 = ~(DATA_IN_3_ & U351); 
assign U559 = ~(DATA_IN_2_ & U351); 
assign U561 = ~(DATA_IN_1_ & U351); 
assign U563 = ~(DATA_IN_0_ & U351); 
assign U565 = ~(U351 & REG4_REG_6__SCAN_IN); 
assign U567 = ~(U351 & REG4_REG_5__SCAN_IN); 
assign U569 = ~(U351 & REG4_REG_4__SCAN_IN); 
assign U571 = ~(U351 & REG4_REG_3__SCAN_IN); 
assign U573 = ~(U351 & REG4_REG_2__SCAN_IN); 
assign U575 = ~(U351 & REG4_REG_1__SCAN_IN); 
assign U577 = ~(U351 & REG4_REG_0__SCAN_IN); 
assign ADD_65_U11 = ~(ADD_65_U10 & ADD_65_U9); 
assign ADD_77_U11 = ~(ADD_77_U10 & ADD_77_U9); 
assign LT_90_U22 = ~(DATA_IN_1_ & LT_90_U9); 
assign LT_90_U24 = ~(LT_90_U8 & RMIN_REG_1__SCAN_IN); 
assign LT_90_U25 = ~(LT_90_U11 & RMIN_REG_2__SCAN_IN); 
assign LT_90_U27 = ~(DATA_IN_2_ & LT_90_U10); 
assign LT_90_U28 = ~(DATA_IN_3_ & LT_90_U13); 
assign LT_90_U30 = ~(LT_90_U12 & RMIN_REG_3__SCAN_IN); 
assign LT_90_U31 = ~(LT_90_U15 & RMIN_REG_4__SCAN_IN); 
assign LT_90_U33 = ~(DATA_IN_4_ & LT_90_U14); 
assign LT_90_U34 = ~(DATA_IN_5_ & LT_90_U17); 
assign LT_90_U36 = ~(LT_90_U16 & RMIN_REG_5__SCAN_IN); 
assign LT_90_U37 = ~(LT_90_U19 & RMIN_REG_6__SCAN_IN); 
assign LT_90_U39 = ~(DATA_IN_6_ & LT_90_U18); 
assign LT_90_U40 = ~(LT_90_U7 & RMIN_REG_7__SCAN_IN); 
assign LT_90_U42 = ~(DATA_IN_7_ & LT_90_U20); 
assign GT_88_U22 = ~(GT_88_U9 & RMAX_REG_1__SCAN_IN); 
assign GT_88_U24 = ~(DATA_IN_1_ & GT_88_U8); 
assign GT_88_U25 = ~(DATA_IN_2_ & GT_88_U11); 
assign GT_88_U27 = ~(GT_88_U10 & RMAX_REG_2__SCAN_IN); 
assign GT_88_U28 = ~(GT_88_U13 & RMAX_REG_3__SCAN_IN); 
assign GT_88_U30 = ~(DATA_IN_3_ & GT_88_U12); 
assign GT_88_U31 = ~(DATA_IN_4_ & GT_88_U15); 
assign GT_88_U33 = ~(GT_88_U14 & RMAX_REG_4__SCAN_IN); 
assign GT_88_U34 = ~(GT_88_U17 & RMAX_REG_5__SCAN_IN); 
assign GT_88_U36 = ~(DATA_IN_5_ & GT_88_U16); 
assign GT_88_U37 = ~(DATA_IN_6_ & GT_88_U19); 
assign GT_88_U39 = ~(GT_88_U18 & RMAX_REG_6__SCAN_IN); 
assign GT_88_U40 = ~(DATA_IN_7_ & GT_88_U7); 
assign GT_88_U42 = ~(GT_88_U20 & RMAX_REG_7__SCAN_IN); 
assign U280 = ~(U348 & U377); 
assign U353 = ~(U552 & U551); 
assign U354 = ~(U554 & U553); 
assign U355 = ~(U556 & U555); 
assign U356 = ~(U558 & U557); 
assign U357 = ~(U560 & U559); 
assign U358 = ~(U562 & U561); 
assign U359 = ~(U564 & U563); 
assign U360 = ~(U566 & U565); 
assign U361 = ~(U568 & U567); 
assign U362 = ~(U570 & U569); 
assign U363 = ~(U572 & U571); 
assign U364 = ~(U574 & U573); 
assign U365 = ~(U576 & U575); 
assign U366 = ~(U578 & U577); 
assign U376 = ~U348; 
assign U422 = ~(U278 & DATA_IN_7_); 
assign U423 = ~(U421 & RLAST_REG_7__SCAN_IN); 
assign U424 = ~(U278 & DATA_IN_6_); 
assign U425 = ~(U421 & RLAST_REG_6__SCAN_IN); 
assign U426 = ~(U278 & DATA_IN_5_); 
assign U427 = ~(U421 & RLAST_REG_5__SCAN_IN); 
assign U428 = ~(U278 & DATA_IN_4_); 
assign U429 = ~(U421 & RLAST_REG_4__SCAN_IN); 
assign U430 = ~(U278 & DATA_IN_3_); 
assign U431 = ~(U421 & RLAST_REG_3__SCAN_IN); 
assign U432 = ~(U278 & DATA_IN_2_); 
assign U433 = ~(U421 & RLAST_REG_2__SCAN_IN); 
assign U434 = ~(U278 & DATA_IN_1_); 
assign U435 = ~(U421 & RLAST_REG_1__SCAN_IN); 
assign U436 = ~(U278 & DATA_IN_0_); 
assign U437 = ~(U421 & RLAST_REG_0__SCAN_IN); 
assign ADD_65_U14 = ~(ADD_65_U12 & ADD_65_U13 & ADD_65_U11); 
assign ADD_77_U14 = ~(ADD_77_U12 & ADD_77_U13 & ADD_77_U11); 
assign LT_90_U23 = ~(LT_90_U21 & LT_90_U22 & RMIN_REG_0__SCAN_IN); 
assign GT_88_U23 = ~(DATA_IN_0_ & GT_88_U21 & GT_88_U22); 
assign U279 = U280 & STATO_REG_1__SCAN_IN; 
assign U321 = ~(U437 & U436); 
assign U322 = ~(U435 & U434); 
assign U323 = ~(U433 & U432); 
assign U324 = ~(U431 & U430); 
assign U325 = ~(U429 & U428); 
assign U326 = ~(U427 & U426); 
assign U327 = ~(U425 & U424); 
assign U328 = ~(U423 & U422); 
assign U378 = ~U280; 
assign U438 = ~(U376 & DATA_IN_7_); 
assign U440 = ~(U376 & DATA_IN_6_); 
assign U442 = ~(U376 & DATA_IN_5_); 
assign U444 = ~(U376 & DATA_IN_4_); 
assign U446 = ~(U376 & DATA_IN_3_); 
assign U448 = ~(U376 & DATA_IN_2_); 
assign U450 = ~(U376 & DATA_IN_1_); 
assign U452 = ~(U376 & DATA_IN_0_); 
assign U454 = ~(U376 & REG1_REG_7__SCAN_IN); 
assign U456 = ~(U376 & REG1_REG_6__SCAN_IN); 
assign U458 = ~(U376 & REG1_REG_5__SCAN_IN); 
assign U460 = ~(U376 & REG1_REG_4__SCAN_IN); 
assign U462 = ~(U376 & REG1_REG_3__SCAN_IN); 
assign U464 = ~(U376 & REG1_REG_2__SCAN_IN); 
assign U466 = ~(U376 & REG1_REG_1__SCAN_IN); 
assign U468 = ~(U376 & REG1_REG_0__SCAN_IN); 
assign U470 = ~(U376 & REG2_REG_7__SCAN_IN); 
assign U472 = ~(U376 & REG2_REG_6__SCAN_IN); 
assign U474 = ~(U376 & REG2_REG_5__SCAN_IN); 
assign U476 = ~(U376 & REG2_REG_4__SCAN_IN); 
assign U478 = ~(U376 & REG2_REG_3__SCAN_IN); 
assign U480 = ~(U376 & REG2_REG_2__SCAN_IN); 
assign U482 = ~(U376 & REG2_REG_1__SCAN_IN); 
assign U484 = ~(U376 & REG2_REG_0__SCAN_IN); 
assign U486 = ~(U376 & REG3_REG_7__SCAN_IN); 
assign U488 = ~(U376 & REG3_REG_6__SCAN_IN); 
assign U490 = ~(U376 & REG3_REG_5__SCAN_IN); 
assign U492 = ~(U376 & REG3_REG_4__SCAN_IN); 
assign U494 = ~(U376 & REG3_REG_3__SCAN_IN); 
assign U496 = ~(U376 & REG3_REG_2__SCAN_IN); 
assign U498 = ~(U376 & REG3_REG_1__SCAN_IN); 
assign U500 = ~(U376 & REG3_REG_0__SCAN_IN); 
assign ADD_65_U17 = ~(ADD_65_U15 & ADD_65_U16 & ADD_65_U14); 
assign ADD_77_U17 = ~(ADD_77_U15 & ADD_77_U16 & ADD_77_U14); 
assign LT_90_U26 = ~(LT_90_U24 & LT_90_U25 & LT_90_U23); 
assign GT_88_U26 = ~(GT_88_U24 & GT_88_U25 & GT_88_U23); 
assign R179_U6 = ~U359; 
assign R179_U7 = ~U366; 
assign R179_U8 = ~U365; 
assign R179_U9 = ~(U366 & U359); 
assign R179_U10 = ~U358; 
assign R179_U11 = ~U357; 
assign R179_U12 = ~U364; 
assign R179_U13 = ~U356; 
assign R179_U14 = ~U363; 
assign R179_U15 = ~U355; 
assign R179_U16 = ~U362; 
assign R179_U17 = ~U354; 
assign R179_U18 = ~U361; 
assign R179_U25 = ~U360; 
assign R179_U26 = ~U353; 
assign R179_U36 = U357 | U364; 
assign R179_U38 = ~(U364 & U357); 
assign R179_U40 = U356 | U363; 
assign R179_U42 = ~(U363 & U356); 
assign R179_U44 = U355 | U362; 
assign R179_U46 = ~(U362 & U355); 
assign R179_U48 = U354 | U361; 
assign R179_U50 = ~(U361 & U354); 
assign R179_U52 = ~(U361 & U354); 
assign R179_U54 = U361 | U354; 
assign U272 = U279 & U351; 
assign U439 = ~(U378 & REG1_REG_7__SCAN_IN); 
assign U441 = ~(U378 & REG1_REG_6__SCAN_IN); 
assign U443 = ~(U378 & REG1_REG_5__SCAN_IN); 
assign U445 = ~(U378 & REG1_REG_4__SCAN_IN); 
assign U447 = ~(U378 & REG1_REG_3__SCAN_IN); 
assign U449 = ~(U378 & REG1_REG_2__SCAN_IN); 
assign U451 = ~(U378 & REG1_REG_1__SCAN_IN); 
assign U453 = ~(U378 & REG1_REG_0__SCAN_IN); 
assign U455 = ~(U378 & REG2_REG_7__SCAN_IN); 
assign U457 = ~(U378 & REG2_REG_6__SCAN_IN); 
assign U459 = ~(U378 & REG2_REG_5__SCAN_IN); 
assign U461 = ~(U378 & REG2_REG_4__SCAN_IN); 
assign U463 = ~(U378 & REG2_REG_3__SCAN_IN); 
assign U465 = ~(U378 & REG2_REG_2__SCAN_IN); 
assign U467 = ~(U378 & REG2_REG_1__SCAN_IN); 
assign U469 = ~(U378 & REG2_REG_0__SCAN_IN); 
assign U471 = ~(U378 & REG3_REG_7__SCAN_IN); 
assign U473 = ~(U378 & REG3_REG_6__SCAN_IN); 
assign U475 = ~(U378 & REG3_REG_5__SCAN_IN); 
assign U477 = ~(U378 & REG3_REG_4__SCAN_IN); 
assign U479 = ~(U378 & REG3_REG_3__SCAN_IN); 
assign U481 = ~(U378 & REG3_REG_2__SCAN_IN); 
assign U483 = ~(U378 & REG3_REG_1__SCAN_IN); 
assign U485 = ~(U378 & REG3_REG_0__SCAN_IN); 
assign U487 = ~(U378 & REG4_REG_7__SCAN_IN); 
assign U489 = ~(U378 & REG4_REG_6__SCAN_IN); 
assign U491 = ~(U378 & REG4_REG_5__SCAN_IN); 
assign U493 = ~(U378 & REG4_REG_4__SCAN_IN); 
assign U495 = ~(U378 & REG4_REG_3__SCAN_IN); 
assign U497 = ~(U378 & REG4_REG_2__SCAN_IN); 
assign U499 = ~(U378 & REG4_REG_1__SCAN_IN); 
assign U501 = ~(U378 & REG4_REG_0__SCAN_IN); 
assign U506 = ~(U378 & DATA_OUT_REG_7__SCAN_IN); 
assign U511 = ~(U378 & DATA_OUT_REG_6__SCAN_IN); 
assign U517 = ~(U378 & DATA_OUT_REG_5__SCAN_IN); 
assign U523 = ~(U378 & DATA_OUT_REG_4__SCAN_IN); 
assign U529 = ~(U378 & DATA_OUT_REG_3__SCAN_IN); 
assign U535 = ~(U378 & DATA_OUT_REG_2__SCAN_IN); 
assign U541 = ~(U378 & DATA_OUT_REG_1__SCAN_IN); 
assign U547 = ~(U378 & DATA_OUT_REG_0__SCAN_IN); 
assign ADD_65_U20 = ~(ADD_65_U18 & ADD_65_U19 & ADD_65_U17); 
assign ADD_77_U20 = ~(ADD_77_U18 & ADD_77_U19 & ADD_77_U17); 
assign LT_90_U29 = ~(LT_90_U27 & LT_90_U28 & LT_90_U26); 
assign GT_88_U29 = ~(GT_88_U27 & GT_88_U28 & GT_88_U26); 
assign R179_U32 = ~R179_U9; 
assign R179_U33 = ~(R179_U10 & R179_U9); 
assign R179_U57 = ~(U360 & R179_U26); 
assign R179_U58 = ~(U353 & R179_U25); 
assign R179_U59 = ~(U360 & R179_U26); 
assign R179_U60 = ~(U353 & R179_U25); 
assign R179_U62 = ~(U361 & R179_U17); 
assign R179_U63 = ~(U354 & R179_U18); 
assign R179_U64 = ~(U361 & R179_U17); 
assign R179_U65 = ~(U354 & R179_U18); 
assign R179_U69 = ~(U362 & R179_U15); 
assign R179_U70 = ~(U355 & R179_U16); 
assign R179_U71 = ~(U362 & R179_U15); 
assign R179_U72 = ~(U355 & R179_U16); 
assign R179_U76 = ~(U363 & R179_U13); 
assign R179_U77 = ~(U356 & R179_U14); 
assign R179_U78 = ~(U363 & R179_U13); 
assign R179_U79 = ~(U356 & R179_U14); 
assign R179_U83 = ~(U364 & R179_U11); 
assign R179_U84 = ~(U357 & R179_U12); 
assign R179_U85 = ~(U364 & R179_U11); 
assign R179_U86 = ~(U357 & R179_U12); 
assign R179_U90 = ~(U365 & R179_U9); 
assign R179_U93 = ~(U358 & R179_U9 & R179_U8); 
assign R179_U95 = ~(U366 & R179_U6); 
assign R179_U96 = ~(U359 & R179_U7); 
assign U275 = AVERAGE & ENABLE & U272; 
assign U277 = U272 & U350; 
assign U289 = ~(U501 & U500); 
assign U290 = ~(U499 & U498); 
assign U291 = ~(U497 & U496); 
assign U292 = ~(U495 & U494); 
assign U293 = ~(U493 & U492); 
assign U294 = ~(U491 & U490); 
assign U295 = ~(U489 & U488); 
assign U296 = ~(U487 & U486); 
assign U297 = ~(U485 & U484); 
assign U298 = ~(U483 & U482); 
assign U299 = ~(U481 & U480); 
assign U300 = ~(U479 & U478); 
assign U301 = ~(U477 & U476); 
assign U302 = ~(U475 & U474); 
assign U303 = ~(U473 & U472); 
assign U304 = ~(U471 & U470); 
assign U305 = ~(U469 & U468); 
assign U306 = ~(U467 & U466); 
assign U307 = ~(U465 & U464); 
assign U308 = ~(U463 & U462); 
assign U309 = ~(U461 & U460); 
assign U310 = ~(U459 & U458); 
assign U311 = ~(U457 & U456); 
assign U312 = ~(U455 & U454); 
assign U313 = ~(U453 & U452); 
assign U314 = ~(U451 & U450); 
assign U315 = ~(U449 & U448); 
assign U316 = ~(U447 & U446); 
assign U317 = ~(U445 & U444); 
assign U318 = ~(U443 & U442); 
assign U319 = ~(U441 & U440); 
assign U320 = ~(U439 & U438); 
assign ADD_65_U22 = ~(ADD_65_U20 & ADD_65_U21); 
assign ADD_77_U22 = ~(ADD_77_U20 & ADD_77_U21); 
assign LT_90_U32 = ~(LT_90_U30 & LT_90_U31 & LT_90_U29); 
assign GT_88_U32 = ~(GT_88_U30 & GT_88_U31 & GT_88_U29); 
assign R179_U20 = ~(R179_U96 & R179_U95); 
assign R179_U30 = ~(U358 & R179_U32); 
assign R179_U34 = ~(U365 & R179_U33); 
assign R179_U61 = ~(R179_U60 & R179_U59); 
assign R179_U66 = ~(R179_U65 & R179_U64); 
assign R179_U73 = ~(R179_U72 & R179_U71); 
assign R179_U80 = ~(R179_U79 & R179_U78); 
assign R179_U87 = ~(R179_U86 & R179_U85); 
assign R179_U91 = ~(R179_U32 & R179_U8); 
assign U502 = ~(U277 & RLAST_REG_7__SCAN_IN); 
assign U503 = ~(U275 & REG4_REG_7__SCAN_IN); 
assign U507 = ~(U277 & RLAST_REG_6__SCAN_IN); 
assign U508 = ~(U275 & REG4_REG_6__SCAN_IN); 
assign U512 = ~(U277 & RLAST_REG_5__SCAN_IN); 
assign U514 = ~(U275 & REG4_REG_5__SCAN_IN); 
assign U518 = ~(U277 & RLAST_REG_4__SCAN_IN); 
assign U520 = ~(U275 & REG4_REG_4__SCAN_IN); 
assign U524 = ~(U277 & RLAST_REG_3__SCAN_IN); 
assign U526 = ~(U275 & REG4_REG_3__SCAN_IN); 
assign U530 = ~(U277 & RLAST_REG_2__SCAN_IN); 
assign U532 = ~(U275 & REG4_REG_2__SCAN_IN); 
assign U536 = ~(U277 & RLAST_REG_1__SCAN_IN); 
assign U538 = ~(U275 & REG4_REG_1__SCAN_IN); 
assign U542 = ~(U277 & RLAST_REG_0__SCAN_IN); 
assign U544 = ~(U275 & REG4_REG_0__SCAN_IN); 
assign SUB_82_U21 = ~R179_U20; 
assign ADD_65_U23 = ~(ADD_65_U22 & ADD_65_U8); 
assign ADD_77_U23 = ~(ADD_77_U22 & ADD_77_U8); 
assign LT_90_U35 = ~(LT_90_U33 & LT_90_U34 & LT_90_U32); 
assign GT_88_U35 = ~(GT_88_U33 & GT_88_U34 & GT_88_U32); 
assign R179_U29 = ~(R179_U30 & R179_U34); 
assign R179_U31 = ~R179_U30; 
assign R179_U92 = ~(R179_U91 & R179_U90); 
assign SUB_70_U21 = ~R179_U20; 
assign U370 = U532 & U530; 
assign U371 = U538 & U536; 
assign U372 = U544 & U542; 
assign ADD_65_U7 = ~(ADD_65_U24 & ADD_65_U23); 
assign ADD_77_U7 = ~(ADD_77_U24 & ADD_77_U23); 
assign LT_90_U38 = ~(LT_90_U36 & LT_90_U37 & LT_90_U35); 
assign GT_88_U38 = ~(GT_88_U36 & GT_88_U37 & GT_88_U35); 
assign R179_U35 = ~R179_U29; 
assign R179_U37 = ~(R179_U36 & R179_U29); 
assign R179_U56 = ~(R179_U92 & R179_U10); 
assign R179_U88 = ~(R179_U84 & R179_U83 & R179_U29); 
assign R179_U94 = ~(R179_U31 & U365); 
assign ADD_65_U4 = ADD_65_U7 & RMAX_REG_6__SCAN_IN; 
assign ADD_65_U25 = ~ADD_65_U7; 
assign ADD_77_U4 = DATA_IN_6_ & ADD_77_U7; 
assign ADD_77_U25 = ~ADD_77_U7; 
assign LT_90_U41 = ~(LT_90_U39 & LT_90_U40 & LT_90_U38); 
assign GT_88_U41 = ~(GT_88_U39 & GT_88_U40 & GT_88_U38); 
assign R179_U5 = ~(R179_U94 & R179_U93 & R179_U56); 
assign R179_U28 = ~(R179_U38 & R179_U37); 
assign R179_U89 = ~(R179_U35 & R179_U87); 
assign SUB_82_U20 = ~R179_U5; 
assign SUB_82_U28 = R179_U5 | R179_U20; 
assign SUB_82_U34 = ~(R179_U5 & SUB_82_U21); 
assign ADD_65_U26 = ADD_65_U4 | RMIN_REG_6__SCAN_IN; 
assign ADD_65_U27 = ~(ADD_65_U25 & ADD_65_U6); 
assign ADD_77_U26 = ADD_77_U4 | REG4_REG_6__SCAN_IN; 
assign ADD_77_U27 = ~(ADD_77_U25 & ADD_77_U6); 
assign LT_90_U6 = ~(LT_90_U41 & LT_90_U42); 
assign GT_88_U6 = ~(GT_88_U41 & GT_88_U42); 
assign R179_U24 = ~(R179_U89 & R179_U88); 
assign R179_U39 = ~R179_U28; 
assign R179_U41 = ~(R179_U40 & R179_U28); 
assign R179_U81 = ~(R179_U77 & R179_U76 & R179_U28); 
assign SUB_70_U20 = ~R179_U5; 
assign SUB_70_U28 = R179_U5 | R179_U20; 
assign SUB_70_U34 = ~(R179_U5 & SUB_70_U21); 
assign U347 = ~GT_88_U6; 
assign U379 = ~(GT_88_U6 & STATO_REG_1__SCAN_IN); 
assign U381 = GT_88_U6 | STATO_REG_0__SCAN_IN; 
assign SUB_82_U10 = R179_U5 | R179_U20 | R179_U24; 
assign SUB_82_U29 = ~(R179_U24 & SUB_82_U28); 
assign SUB_82_U35 = ~(R179_U20 & SUB_82_U20); 
assign ADD_65_U28 = ~(ADD_65_U27 & ADD_65_U26); 
assign ADD_77_U28 = ~(ADD_77_U27 & ADD_77_U26); 
assign R179_U27 = ~(R179_U42 & R179_U41); 
assign R179_U82 = ~(R179_U39 & R179_U80); 
assign SUB_70_U10 = R179_U5 | R179_U20 | R179_U24; 
assign SUB_70_U29 = ~(R179_U24 & SUB_70_U28); 
assign SUB_70_U35 = ~(R179_U20 & SUB_70_U20); 
assign U380 = ~(U345 & U379); 
assign U382 = ~(U374 & U381); 
assign U399 = ~(LT_90_U6 & U347); 
assign U402 = ~(U347 & LT_90_U6 & STATO_REG_1__SCAN_IN); 
assign SUB_82_U6 = SUB_82_U29 & SUB_82_U10; 
assign SUB_82_U15 = ~(SUB_82_U35 & SUB_82_U34); 
assign SUB_82_U22 = ~SUB_82_U10; 
assign ADD_65_U31 = ~(ADD_65_U29 & ADD_65_U28); 
assign ADD_77_U31 = ~(ADD_77_U29 & ADD_77_U28); 
assign R179_U23 = ~(R179_U82 & R179_U81); 
assign R179_U43 = ~R179_U27; 
assign R179_U45 = ~(R179_U44 & R179_U27); 
assign R179_U74 = ~(R179_U70 & R179_U69 & R179_U27); 
assign SUB_70_U6 = SUB_70_U29 & SUB_70_U10; 
assign SUB_70_U15 = ~(SUB_70_U35 & SUB_70_U34); 
assign SUB_70_U22 = ~SUB_70_U10; 
assign U383 = ~(U382 & RMAX_REG_7__SCAN_IN); 
assign U384 = ~(DATA_IN_7_ & U380); 
assign U385 = ~(U382 & RMAX_REG_6__SCAN_IN); 
assign U386 = ~(DATA_IN_6_ & U380); 
assign U387 = ~(U382 & RMAX_REG_5__SCAN_IN); 
assign U388 = ~(DATA_IN_5_ & U380); 
assign U389 = ~(U382 & RMAX_REG_4__SCAN_IN); 
assign U390 = ~(DATA_IN_4_ & U380); 
assign U391 = ~(U382 & RMAX_REG_3__SCAN_IN); 
assign U392 = ~(DATA_IN_3_ & U380); 
assign U393 = ~(U382 & RMAX_REG_2__SCAN_IN); 
assign U394 = ~(DATA_IN_2_ & U380); 
assign U395 = ~(U382 & RMAX_REG_1__SCAN_IN); 
assign U396 = ~(DATA_IN_1_ & U380); 
assign U397 = ~(U382 & RMAX_REG_0__SCAN_IN); 
assign U398 = ~(DATA_IN_0_ & U380); 
assign U400 = ~(U399 & U345); 
assign U403 = ~(U345 & U402); 
assign SUB_82_U18 = ~R179_U23; 
assign SUB_82_U32 = ~(R179_U23 & SUB_82_U10); 
assign ADD_65_U5 = ~(ADD_65_U31 & ADD_65_U30); 
assign ADD_77_U5 = ~(ADD_77_U31 & ADD_77_U30); 
assign SUB_70_166_U19 = ~SUB_70_U6; 
assign SUB_70_166_U20 = ~SUB_70_U15; 
assign SUB_70_166_U30 = SUB_70_U6 | SUB_70_U15; 
assign SUB_82_165_U19 = ~SUB_82_U6; 
assign SUB_82_165_U20 = ~SUB_82_U15; 
assign SUB_82_165_U30 = SUB_82_U6 | SUB_82_U15; 
assign R179_U19 = ~(R179_U46 & R179_U45); 
assign R179_U75 = ~(R179_U43 & R179_U73); 
assign SUB_70_U18 = ~R179_U23; 
assign SUB_70_U32 = ~(R179_U23 & SUB_70_U10); 
assign U337 = ~(U398 & U397); 
assign U338 = ~(U396 & U395); 
assign U339 = ~(U394 & U393); 
assign U340 = ~(U392 & U391); 
assign U341 = ~(U390 & U389); 
assign U342 = ~(U388 & U387); 
assign U343 = ~(U386 & U385); 
assign U344 = ~(U384 & U383); 
assign U401 = ~(U374 & U400); 
assign U404 = ~(DATA_IN_7_ & U403); 
assign U406 = ~(DATA_IN_6_ & U403); 
assign U408 = ~(DATA_IN_5_ & U403); 
assign U410 = ~(DATA_IN_4_ & U403); 
assign U412 = ~(DATA_IN_3_ & U403); 
assign U414 = ~(DATA_IN_2_ & U403); 
assign U416 = ~(DATA_IN_1_ & U403); 
assign U418 = ~(DATA_IN_0_ & U403); 
assign GTE_67_U6 = ~ADD_65_U5; 
assign SUB_82_U26 = ~(SUB_82_U22 & SUB_82_U18); 
assign SUB_82_U33 = ~(SUB_82_U22 & SUB_82_U18); 
assign SUB_70_166_U34 = ~(SUB_70_U6 & SUB_70_166_U20); 
assign SUB_70_166_U35 = ~(SUB_70_U15 & SUB_70_166_U19); 
assign SUB_82_165_U34 = ~(SUB_82_U6 & SUB_82_165_U20); 
assign SUB_82_165_U35 = ~(SUB_82_U15 & SUB_82_165_U19); 
assign GTE_79_U6 = ~ADD_77_U5; 
assign R179_U22 = ~(R179_U75 & R179_U74); 
assign R179_U47 = ~R179_U19; 
assign R179_U49 = ~(R179_U48 & R179_U19); 
assign R179_U67 = ~(R179_U63 & R179_U62 & R179_U19); 
assign SUB_70_U26 = ~(SUB_70_U22 & SUB_70_U18); 
assign SUB_70_U33 = ~(SUB_70_U22 & SUB_70_U18); 
assign U352 = ~GTE_79_U6; 
assign U373 = ~GTE_67_U6; 
assign U405 = ~(U401 & RMIN_REG_7__SCAN_IN); 
assign U407 = ~(U401 & RMIN_REG_6__SCAN_IN); 
assign U409 = ~(U401 & RMIN_REG_5__SCAN_IN); 
assign U411 = ~(U401 & RMIN_REG_4__SCAN_IN); 
assign U413 = ~(U401 & RMIN_REG_3__SCAN_IN); 
assign U415 = ~(U401 & RMIN_REG_2__SCAN_IN); 
assign U417 = ~(U401 & RMIN_REG_1__SCAN_IN); 
assign U419 = ~(U401 & RMIN_REG_0__SCAN_IN); 
assign U548 = ~(ENABLE & U349 & GTE_79_U6); 
assign SUB_82_U14 = ~R179_U22; 
assign SUB_82_U19 = SUB_82_U33 & SUB_82_U32; 
assign SUB_82_U27 = ~(R179_U22 & SUB_82_U26); 
assign SUB_70_166_U16 = ~(SUB_70_166_U35 & SUB_70_166_U34); 
assign SUB_82_165_U16 = ~(SUB_82_165_U35 & SUB_82_165_U34); 
assign R179_U51 = ~(R179_U58 & R179_U57 & R179_U50 & R179_U49); 
assign R179_U53 = ~(R179_U47 & R179_U52); 
assign R179_U68 = ~(R179_U66 & R179_U47); 
assign SUB_70_U14 = ~R179_U22; 
assign SUB_70_U19 = SUB_70_U33 & SUB_70_U32; 
assign SUB_70_U27 = ~(R179_U22 & SUB_70_U26); 
assign U273 = ENABLE & U272 & U349 & U352; 
assign U274 = U279 & RESTART & U373; 
assign U329 = ~(U419 & U418); 
assign U330 = ~(U417 & U416); 
assign U331 = ~(U415 & U414); 
assign U332 = ~(U413 & U412); 
assign U333 = ~(U411 & U410); 
assign U334 = ~(U409 & U408); 
assign U335 = ~(U407 & U406); 
assign U336 = ~(U405 & U404); 
assign U549 = ~(RESTART & U373); 
assign U550 = ~(U548 & U351); 
assign SUB_82_U11 = ~(SUB_82_U22 & SUB_82_U18 & SUB_82_U14); 
assign SUB_70_166_U10 = SUB_70_U6 | SUB_70_U15 | SUB_70_U19; 
assign SUB_70_166_U31 = ~(SUB_70_U19 & SUB_70_166_U30); 
assign SUB_82_165_U10 = SUB_82_U6 | SUB_82_U15 | SUB_82_U19; 
assign SUB_82_165_U31 = ~(SUB_82_U19 & SUB_82_165_U30); 
assign R179_U21 = ~(R179_U68 & R179_U67); 
assign R179_U55 = ~(R179_U54 & R179_U61 & R179_U53); 
assign SUB_70_U11 = ~(SUB_70_U22 & SUB_70_U18 & SUB_70_U14); 
assign U276 = U550 & U549 & U279; 
assign U539 = ~(SUB_70_166_U16 & U274); 
assign U540 = ~(SUB_82_165_U16 & U273); 
assign U545 = ~(SUB_70_U15 & U274); 
assign U546 = ~(SUB_82_U15 & U273); 
assign SUB_82_U7 = SUB_82_U27 & SUB_82_U11; 
assign SUB_82_U13 = ~R179_U21; 
assign SUB_82_U23 = ~SUB_82_U11; 
assign SUB_82_U25 = ~(R179_U21 & SUB_82_U11); 
assign SUB_70_166_U6 = SUB_70_166_U31 & SUB_70_166_U10; 
assign SUB_70_166_U23 = ~SUB_70_166_U10; 
assign SUB_82_165_U6 = SUB_82_165_U31 & SUB_82_165_U10; 
assign SUB_82_165_U23 = ~SUB_82_165_U10; 
assign R179_U4 = R179_U55 & R179_U51; 
assign SUB_70_U7 = SUB_70_U27 & SUB_70_U11; 
assign SUB_70_U13 = ~R179_U21; 
assign SUB_70_U23 = ~SUB_70_U11; 
assign SUB_70_U25 = ~(R179_U21 & SUB_70_U11); 
assign U513 = ~(R179_U4 & U276); 
assign U519 = ~(R179_U21 & U276); 
assign U525 = ~(R179_U22 & U276); 
assign U531 = ~(R179_U23 & U276); 
assign U533 = ~(SUB_70_166_U6 & U274); 
assign U534 = ~(SUB_82_165_U6 & U273); 
assign U537 = ~(R179_U24 & U276); 
assign U543 = ~(R179_U5 & U276); 
assign SUB_82_U12 = ~(SUB_82_U23 & SUB_82_U13); 
assign SUB_82_U16 = ~R179_U4; 
assign SUB_70_166_U17 = ~SUB_70_U7; 
assign SUB_70_166_U32 = ~(SUB_70_U7 & SUB_70_166_U10); 
assign SUB_82_165_U17 = ~SUB_82_U7; 
assign SUB_82_165_U32 = ~(SUB_82_U7 & SUB_82_165_U10); 
assign SUB_70_U12 = ~(SUB_70_U23 & SUB_70_U13); 
assign SUB_70_U16 = ~R179_U4; 
assign U281 = ~(U546 & U545 & U547 & U372 & U543); 
assign U282 = ~(U540 & U539 & U541 & U371 & U537); 
assign U283 = ~(U534 & U533 & U535 & U370 & U531); 
assign U367 = U514 & U512 & U513 & U517; 
assign U368 = U520 & U518 & U519 & U523; 
assign U369 = U526 & U524 & U525; 
assign SUB_82_U8 = SUB_82_U25 & SUB_82_U12; 
assign SUB_82_U24 = ~SUB_82_U12; 
assign SUB_82_U30 = ~(R179_U4 & SUB_82_U12); 
assign SUB_70_166_U28 = ~(SUB_70_166_U23 & SUB_70_166_U17); 
assign SUB_70_166_U33 = ~(SUB_70_166_U23 & SUB_70_166_U17); 
assign SUB_82_165_U28 = ~(SUB_82_165_U23 & SUB_82_165_U17); 
assign SUB_82_165_U33 = ~(SUB_82_165_U23 & SUB_82_165_U17); 
assign SUB_70_U8 = SUB_70_U25 & SUB_70_U12; 
assign SUB_70_U24 = ~SUB_70_U12; 
assign SUB_70_U30 = ~(R179_U4 & SUB_70_U12); 
assign SUB_82_U9 = ~(SUB_82_U24 & SUB_82_U16); 
assign SUB_82_U31 = ~(SUB_82_U24 & SUB_82_U16); 
assign SUB_70_166_U15 = ~SUB_70_U8; 
assign SUB_70_166_U18 = SUB_70_166_U33 & SUB_70_166_U32; 
assign SUB_70_166_U29 = ~(SUB_70_U8 & SUB_70_166_U28); 
assign SUB_82_165_U15 = ~SUB_82_U8; 
assign SUB_82_165_U18 = SUB_82_165_U33 & SUB_82_165_U32; 
assign SUB_82_165_U29 = ~(SUB_82_U8 & SUB_82_165_U28); 
assign SUB_70_U9 = ~(SUB_70_U24 & SUB_70_U16); 
assign SUB_70_U31 = ~(SUB_70_U24 & SUB_70_U16); 
assign U527 = ~(SUB_70_166_U18 & U274); 
assign U528 = ~(SUB_82_165_U18 & U273); 
assign SUB_82_U17 = SUB_82_U31 & SUB_82_U30; 
assign SUB_70_166_U11 = ~(SUB_70_166_U23 & SUB_70_166_U17 & SUB_70_166_U15); 
assign SUB_70_166_U13 = ~SUB_70_U9; 
assign SUB_82_165_U11 = ~(SUB_82_165_U23 & SUB_82_165_U17 & SUB_82_165_U15); 
assign SUB_82_165_U13 = ~SUB_82_U9; 
assign SUB_70_U17 = SUB_70_U31 & SUB_70_U30; 
assign U284 = ~(U528 & U527 & U529 & U369); 
assign SUB_70_166_U7 = SUB_70_166_U29 & SUB_70_166_U11; 
assign SUB_70_166_U14 = ~SUB_70_U17; 
assign SUB_70_166_U24 = ~SUB_70_166_U11; 
assign SUB_70_166_U27 = ~(SUB_70_U17 & SUB_70_166_U11); 
assign SUB_82_165_U7 = SUB_82_165_U29 & SUB_82_165_U11; 
assign SUB_82_165_U14 = ~SUB_82_U17; 
assign SUB_82_165_U24 = ~SUB_82_165_U11; 
assign SUB_82_165_U27 = ~(SUB_82_U17 & SUB_82_165_U11); 
assign U521 = ~(SUB_70_166_U7 & U274); 
assign U522 = ~(SUB_82_165_U7 & U273); 
assign SUB_70_166_U12 = ~(SUB_70_166_U24 & SUB_70_166_U14); 
assign SUB_82_165_U12 = ~(SUB_82_165_U24 & SUB_82_165_U14); 
assign U285 = ~(U522 & U521 & U368); 
assign SUB_70_166_U8 = SUB_70_166_U27 & SUB_70_166_U12; 
assign SUB_70_166_U21 = ~(SUB_70_166_U12 & SUB_70_166_U13); 
assign SUB_70_166_U25 = ~SUB_70_166_U12; 
assign SUB_82_165_U8 = SUB_82_165_U27 & SUB_82_165_U12; 
assign SUB_82_165_U21 = ~(SUB_82_165_U12 & SUB_82_165_U13); 
assign SUB_82_165_U25 = ~SUB_82_165_U12; 
assign U515 = ~(SUB_70_166_U8 & U274); 
assign U516 = ~(SUB_82_165_U8 & U273); 
assign SUB_70_166_U22 = ~SUB_70_166_U21; 
assign SUB_70_166_U26 = ~(SUB_70_U9 & SUB_70_166_U25); 
assign SUB_82_165_U22 = ~SUB_82_165_U21; 
assign SUB_82_165_U26 = ~(SUB_82_U9 & SUB_82_165_U25); 
assign U286 = ~(U516 & U515 & U367); 
assign U504 = ~(SUB_70_166_U22 & U274); 
assign U505 = ~(SUB_82_165_U22 & U273); 
assign SUB_70_166_U9 = ~(SUB_70_166_U21 & SUB_70_166_U26); 
assign SUB_82_165_U9 = ~(SUB_82_165_U21 & SUB_82_165_U26); 
assign U288 = ~(U503 & U502 & U504 & U506 & U505); 
assign U509 = ~(SUB_70_166_U9 & U274); 
assign U510 = ~(SUB_82_165_U9 & U273); 
assign U287 = ~(U508 & U507 & U509 & U511 & U510); 
endmodule 
