module b08_C( O_REG_0__SCAN_IN, START, I_7_, I_6_, I_5_, I_4_, I_3_, I_2_, I_1_, I_0_, STATO_REG_1__SCAN_IN, STATO_REG_0__SCAN_IN, MAR_REG_2__SCAN_IN, MAR_REG_1__SCAN_IN, MAR_REG_0__SCAN_IN, IN_R_REG_7__SCAN_IN, IN_R_REG_6__SCAN_IN, IN_R_REG_5__SCAN_IN, IN_R_REG_4__SCAN_IN, IN_R_REG_3__SCAN_IN, IN_R_REG_2__SCAN_IN, IN_R_REG_1__SCAN_IN, IN_R_REG_0__SCAN_IN, OUT_R_REG_3__SCAN_IN, OUT_R_REG_2__SCAN_IN, OUT_R_REG_1__SCAN_IN, OUT_R_REG_0__SCAN_IN, O_REG_3__SCAN_IN, O_REG_2__SCAN_IN, O_REG_1__SCAN_IN, U183, U184, U185, U186, U187, U188, U189, U206, U207, U208, U209, U210, U211, U212, U213, U214, U215, U216, U217, U218, U219); 
input O_REG_0__SCAN_IN, START, I_7_, I_6_, I_5_, I_4_, I_3_, I_2_, I_1_, I_0_, STATO_REG_1__SCAN_IN, STATO_REG_0__SCAN_IN, MAR_REG_2__SCAN_IN, MAR_REG_1__SCAN_IN, MAR_REG_0__SCAN_IN, IN_R_REG_7__SCAN_IN, IN_R_REG_6__SCAN_IN, IN_R_REG_5__SCAN_IN, IN_R_REG_4__SCAN_IN, IN_R_REG_3__SCAN_IN, IN_R_REG_2__SCAN_IN, IN_R_REG_1__SCAN_IN, IN_R_REG_0__SCAN_IN, OUT_R_REG_3__SCAN_IN, OUT_R_REG_2__SCAN_IN, OUT_R_REG_1__SCAN_IN, OUT_R_REG_0__SCAN_IN, O_REG_3__SCAN_IN, O_REG_2__SCAN_IN, O_REG_1__SCAN_IN; 
output U183, U184, U185, U186, U187, U188, U189, U206, U207, U208, U209, U210, U211, U212, U213, U214, U215, U216, U217, U218, U219; 
wire U176, U177, U178, U179, U180, U181, U182, U190, U191, U192, U193, U194, U195, U196, U197, U198, U199, U200, U201, U202, U203, U204, U205, U220, U221, U222, U223, U224, U225, U226, U227, U228, U229, U230, U231, U232, U233, U234, U235, U236, U237, U238, U239, U240, U241, U242, U243, U244, U245, U246, U247, U248, U249, U250, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, U280, U281, U282, U283, U284, U285, U286, U287, U288, U289, U290, U291, U292, U293, U294, U295, U296, U297, U298, U299, U300, U301, U302, U303, U304, U305, U306, U307, U308, U309, U310, U311, U312, U313, U314, U315, U316, U317, U318, U319, U320, U321, U322, U323, U324; 
assign U177 = STATO_REG_1__SCAN_IN & STATO_REG_0__SCAN_IN; 
assign U178 = MAR_REG_1__SCAN_IN & MAR_REG_0__SCAN_IN; 
assign U190 = ~STATO_REG_1__SCAN_IN; 
assign U191 = ~STATO_REG_0__SCAN_IN; 
assign U192 = ~MAR_REG_1__SCAN_IN; 
assign U193 = ~MAR_REG_0__SCAN_IN; 
assign U194 = ~MAR_REG_2__SCAN_IN; 
assign U196 = ~START; 
assign U222 = ~IN_R_REG_7__SCAN_IN; 
assign U224 = ~IN_R_REG_6__SCAN_IN; 
assign U225 = ~IN_R_REG_5__SCAN_IN; 
assign U226 = ~IN_R_REG_4__SCAN_IN; 
assign U227 = ~IN_R_REG_3__SCAN_IN; 
assign U228 = ~IN_R_REG_2__SCAN_IN; 
assign U229 = ~IN_R_REG_1__SCAN_IN; 
assign U230 = ~IN_R_REG_0__SCAN_IN; 
assign U247 = MAR_REG_2__SCAN_IN | MAR_REG_1__SCAN_IN | MAR_REG_0__SCAN_IN; 
assign U195 = ~(U178 & MAR_REG_2__SCAN_IN); 
assign U198 = ~(U178 & U194); 
assign U204 = ~(U191 & STATO_REG_1__SCAN_IN); 
assign U223 = ~(U190 & STATO_REG_0__SCAN_IN); 
assign U245 = ~(U193 & STATO_REG_1__SCAN_IN); 
assign U248 = ~(U192 & MAR_REG_2__SCAN_IN & MAR_REG_0__SCAN_IN); 
assign U249 = ~(U194 & U192 & MAR_REG_0__SCAN_IN); 
assign U250 = ~(U192 & U193 & MAR_REG_2__SCAN_IN); 
assign U251 = ~(U194 & U193 & MAR_REG_1__SCAN_IN); 
assign U254 = ~(U193 & MAR_REG_2__SCAN_IN & MAR_REG_1__SCAN_IN); 
assign U284 = ~(U177 & U192 & MAR_REG_0__SCAN_IN); 
assign U285 = ~(U177 & U193); 
assign U179 = U195 & U251; 
assign U181 = U248 & U250; 
assign U202 = ~(U251 & U254); 
assign U233 = ~U204; 
assign U234 = ~U223; 
assign U235 = ~U195; 
assign U241 = ~U198; 
assign U278 = ~(U250 & U249 & U247 & U198); 
assign U287 = ~(U223 & IN_R_REG_7__SCAN_IN); 
assign U289 = ~(U223 & IN_R_REG_6__SCAN_IN); 
assign U291 = ~(U223 & IN_R_REG_5__SCAN_IN); 
assign U293 = ~(U223 & IN_R_REG_4__SCAN_IN); 
assign U295 = ~(U223 & IN_R_REG_3__SCAN_IN); 
assign U297 = ~(U223 & IN_R_REG_2__SCAN_IN); 
assign U299 = ~(U223 & IN_R_REG_1__SCAN_IN); 
assign U301 = ~(U223 & IN_R_REG_0__SCAN_IN); 
assign U182 = U179 & U254; 
assign U199 = ~(U179 & U250); 
assign U200 = ~(U181 & U198); 
assign U205 = ~(U235 & U196); 
assign U238 = ~(U235 & STATO_REG_1__SCAN_IN); 
assign U244 = ~(U177 & U241); 
assign U255 = ~U202; 
assign U270 = ~(U179 & U248 & U198 & U227); 
assign U288 = ~(I_7_ & U234); 
assign U290 = ~(I_6_ & U234); 
assign U292 = ~(I_5_ & U234); 
assign U294 = ~(I_4_ & U234); 
assign U296 = ~(I_3_ & U234); 
assign U298 = ~(I_2_ & U234); 
assign U300 = ~(I_1_ & U234); 
assign U302 = ~(I_0_ & U234); 
assign U197 = ~(U238 & STATO_REG_0__SCAN_IN); 
assign U208 = ~(U288 & U287); 
assign U209 = ~(U290 & U289); 
assign U210 = ~(U292 & U291); 
assign U211 = ~(U294 & U293); 
assign U212 = ~(U296 & U295); 
assign U213 = ~(U298 & U297); 
assign U214 = ~(U300 & U299); 
assign U215 = ~(U302 & U301); 
assign U236 = ~U205; 
assign U237 = ~(U205 & STATO_REG_0__SCAN_IN); 
assign U252 = ~U199; 
assign U253 = ~U200; 
assign U260 = ~(U182 & U181); 
assign U268 = ~(U182 & U198); 
assign U315 = ~(U200 & IN_R_REG_4__SCAN_IN); 
assign U180 = U252 & U249; 
assign U189 = ~(U223 & U204 & U237); 
assign U201 = ~(U253 & U195); 
assign U203 = ~(U179 & U249 & U253); 
assign U231 = ~(U236 & STATO_REG_1__SCAN_IN & STATO_REG_0__SCAN_IN); 
assign U239 = ~U197; 
assign U240 = ~(START & U197); 
assign U256 = ~(U253 & U247); 
assign U286 = ~(U197 & MAR_REG_0__SCAN_IN); 
assign U304 = ~(U255 & U253 & IN_R_REG_7__SCAN_IN); 
assign U305 = ~(U182 & U253 & U225); 
assign U310 = ~(U268 & U230); 
assign U316 = ~(U260 & U226); 
assign U188 = ~(U204 & U240); 
assign U207 = ~(U286 & U285); 
assign U242 = ~(U239 & U190); 
assign U246 = ~(U239 & U245); 
assign U257 = ~(U180 & U198); 
assign U259 = ~U203; 
assign U261 = ~(U249 & U247 & U316 & U315); 
assign U262 = ~U201; 
assign U263 = ~(U180 & U254); 
assign U282 = ~U231; 
assign U303 = ~(U248 & U247 & U180 & U222); 
assign U307 = ~(U203 & U229); 
assign U311 = ~(U201 & IN_R_REG_2__SCAN_IN); 
assign U313 = ~(U256 & IN_R_REG_6__SCAN_IN); 
assign U317 = ~(U231 & O_REG_3__SCAN_IN); 
assign U319 = ~(U231 & O_REG_2__SCAN_IN); 
assign U321 = ~(U231 & O_REG_1__SCAN_IN); 
assign U323 = ~(U231 & O_REG_0__SCAN_IN); 
assign U243 = ~(U242 & MAR_REG_2__SCAN_IN); 
assign U265 = ~(U262 & U254); 
assign U267 = ~(U262 & U249); 
assign U283 = ~(U246 & MAR_REG_1__SCAN_IN); 
assign U306 = ~(U259 & U247 & IN_R_REG_5__SCAN_IN); 
assign U312 = ~(U263 & U228); 
assign U314 = ~(U257 & U224); 
assign U318 = ~(U282 & OUT_R_REG_3__SCAN_IN); 
assign U320 = ~(U282 & OUT_R_REG_2__SCAN_IN); 
assign U322 = ~(U282 & OUT_R_REG_1__SCAN_IN); 
assign U324 = ~(U282 & OUT_R_REG_0__SCAN_IN); 
assign U187 = ~(U244 & U243); 
assign U206 = ~(U284 & U283); 
assign U216 = ~(U318 & U317); 
assign U217 = ~(U320 & U319); 
assign U218 = ~(U322 & U321); 
assign U219 = ~(U324 & U323); 
assign U221 = U306 & U305 & U304 & U303; 
assign U258 = ~(U314 & U313 & U254); 
assign U264 = ~(U312 & U311 & U247); 
assign U308 = ~(U265 & IN_R_REG_1__SCAN_IN); 
assign U309 = ~(U267 & IN_R_REG_0__SCAN_IN); 
assign U266 = ~(U308 & U307 & U247); 
assign U269 = ~(U310 & U309 & U247); 
assign U220 = U233 & U270 & U221 & U269 & U266; 
assign U271 = ~(U261 & U258 & U264 & U220); 
assign U272 = ~(U223 & U271); 
assign U176 = U272 & STATO_REG_1__SCAN_IN; 
assign U273 = ~(U190 & U272); 
assign U232 = ~(U176 & U202); 
assign U274 = ~(U176 & U256); 
assign U275 = ~(U273 & OUT_R_REG_3__SCAN_IN); 
assign U276 = ~(U176 & U199); 
assign U277 = ~(U273 & OUT_R_REG_2__SCAN_IN); 
assign U279 = ~(U176 & U278); 
assign U280 = ~(U273 & OUT_R_REG_1__SCAN_IN); 
assign U281 = ~(U273 & OUT_R_REG_0__SCAN_IN); 
assign U183 = ~(U232 & U281); 
assign U184 = ~(U279 & U232 & U280); 
assign U185 = ~(U277 & U276); 
assign U186 = ~(U274 & U232 & U275); 
endmodule 
