module b05_C( STATO_REG_2__SCAN_IN, START, STATO_REG_1__SCAN_IN, STATO_REG_0__SCAN_IN, FLAG_REG_SCAN_IN, RES_DISP_REG_SCAN_IN, EN_DISP_REG_SCAN_IN, MAX_REG_0__SCAN_IN, MAX_REG_1__SCAN_IN, MAX_REG_2__SCAN_IN, MAX_REG_3__SCAN_IN, MAX_REG_4__SCAN_IN, MAX_REG_5__SCAN_IN, MAX_REG_6__SCAN_IN, MAX_REG_7__SCAN_IN, MAX_REG_8__SCAN_IN, TEMP_REG_0__SCAN_IN, TEMP_REG_1__SCAN_IN, TEMP_REG_2__SCAN_IN, TEMP_REG_3__SCAN_IN, TEMP_REG_4__SCAN_IN, TEMP_REG_5__SCAN_IN, TEMP_REG_6__SCAN_IN, TEMP_REG_7__SCAN_IN, TEMP_REG_8__SCAN_IN, MAR_REG_0__SCAN_IN, MAR_REG_1__SCAN_IN, MAR_REG_2__SCAN_IN, MAR_REG_3__SCAN_IN, MAR_REG_4__SCAN_IN, NUM_REG_0__SCAN_IN, NUM_REG_1__SCAN_IN, NUM_REG_2__SCAN_IN, NUM_REG_3__SCAN_IN, NUM_REG_4__SCAN_IN, U590, U591, U643, U644, U645, U646, U647, U648, U649, U650, U651, U652, U653, U654, U655, U656, U657, U658, U659, U660, U661, U662, U663, U664, U665, U666, U667, U668, U669, U670, U671, U672, U673, U674, U675, U676, U677, U678, U679, U680, U727, U728, U729, U730, U731, U732, U733, U734, U735, U736, U737, U738, U739, U740, U741, U742, U743, U744, U792); 
input STATO_REG_2__SCAN_IN, START, STATO_REG_1__SCAN_IN, STATO_REG_0__SCAN_IN, FLAG_REG_SCAN_IN, RES_DISP_REG_SCAN_IN, EN_DISP_REG_SCAN_IN, MAX_REG_0__SCAN_IN, MAX_REG_1__SCAN_IN, MAX_REG_2__SCAN_IN, MAX_REG_3__SCAN_IN, MAX_REG_4__SCAN_IN, MAX_REG_5__SCAN_IN, MAX_REG_6__SCAN_IN, MAX_REG_7__SCAN_IN, MAX_REG_8__SCAN_IN, TEMP_REG_0__SCAN_IN, TEMP_REG_1__SCAN_IN, TEMP_REG_2__SCAN_IN, TEMP_REG_3__SCAN_IN, TEMP_REG_4__SCAN_IN, TEMP_REG_5__SCAN_IN, TEMP_REG_6__SCAN_IN, TEMP_REG_7__SCAN_IN, TEMP_REG_8__SCAN_IN, MAR_REG_0__SCAN_IN, MAR_REG_1__SCAN_IN, MAR_REG_2__SCAN_IN, MAR_REG_3__SCAN_IN, MAR_REG_4__SCAN_IN, NUM_REG_0__SCAN_IN, NUM_REG_1__SCAN_IN, NUM_REG_2__SCAN_IN, NUM_REG_3__SCAN_IN, NUM_REG_4__SCAN_IN; 
output U590, U591, U643, U644, U645, U646, U647, U648, U649, U650, U651, U652, U653, U654, U655, U656, U657, U658, U659, U660, U661, U662, U663, U664, U665, U666, U667, U668, U669, U670, U671, U672, U673, U674, U675, U676, U677, U678, U679, U680, U727, U728, U729, U730, U731, U732, U733, U734, U735, U736, U737, U738, U739, U740, U741, U742, U743, U744, U792; 
wire U587, U588, U589, U592, U593, U594, U595, U596, U597, U598, U599, U600, U601, U602, U603, U604, U605, U606, U607, U608, U609, U610, U611, U612, U613, U614, U615, U616, U617, U618, U619, U620, U621, U622, U623, U624, U625, U626, U627, U628, U629, U630, U631, U632, U633, U634, U635, U636, U637, U638, U639, U640, U641, U642, U681, U682, U683, U684, U685, U686, U687, U688, U689, U690, U691, U692, U693, U694, U695, U696, U697, U698, U699, U700, U701, U702, U703, U704, U705, U706, U707, U708, U709, U710, U711, U712, U713, U714, U715, U716, U717, U718, U719, U720, U721, U722, U723, U724, U725, U726, U745, U746, U747, U748, U749, U750, U751, U752, U753, U754, U755, U756, U757, U758, U759, U760, U761, U762, U763, U764, U765, U766, U767, U768, U769, U770, U771, U772, U773, U774, U775, U776, U777, U778, U779, U780, U781, U782, U783, U784, U785, U786, U787, U788, U789, U790, U791, U793, U794, U795, U796, U797, U798, U799, U800, U801, U802, U803, U804, U805, U806, U807, U808, U809, U810, U811, U812, U813, U814, U815, U816, U817, U818, U819, U820, U821, U822, U823, U824, U825, U826, U827, U828, U829, U830, U831, U832, U833, U834, U835, U836, U837, U838, U839, U840, U841, U842, U843, U844, U845, U846, U847, U848, U849, U850, U851, U852, U853, U854, U855, U856, U857, U858, U859, U860, U861, U862, U863, U864, U865, U866, U867, U868, U869, U870, U871, U872, U873, U874, U875, U876, U877, U878, U879, U880, U881, U882, U883, U884, U885, U886, U887, U888, U889, U890, U891, U892, U893, U894, U895, U896, U897, U898, U899, U900, U901, U902, U903, U904, U905, U906, U907, U908, U909, U910, U911, U912, U913, U914, U915, U916, U917, U918, U919, U920, U921, U922, U923, U924, U925, U926, U927, U928, U929, U930, U931, U932, U933, U934, U935, U936, U937, U938, U939, U940, U941, U942, U943, U944, U945, U946, U947, U948, U949, U950, U951, U952, U953, U954, U955, U956, U957, U958, U959, U960, U961, U962, U963, U964, U965, U966, U967, U968, U969, U970, U971, U972, U973, U974, U975, U976, U977, U978, U979, U980, U981, U982, U983, U984, U985, U986, U987, U988, U989, U990, U991, U992, U993, U994, U995, U996, U997, U998, U999, U1000, U1001, U1002, U1003, U1004, U1005, U1006, U1007, U1008, U1009, U1010, U1011, U1012, U1013, U1014, U1015, U1016, U1017, U1018, U1019, U1020, U1021, U1022, U1023, U1024, U1025, U1026, U1027, U1028, U1029, U1030, U1031, U1032, U1033, U1034, U1035, U1036, U1037, U1038, U1039, U1040, U1041, GT_138_U8, GT_138_U7, GT_138_U6, GT_118_U9, GT_118_U8, GT_118_U7, GT_118_U6, GT_166_U9, SUB_103_U6, SUB_103_U7, SUB_103_U8, SUB_103_U9, SUB_103_U10, SUB_103_U11, SUB_103_U12, SUB_103_U13, SUB_103_U14, SUB_103_U15, SUB_103_U16, SUB_103_U17, SUB_103_U18, SUB_103_U19, SUB_103_U20, SUB_103_U21, SUB_103_U22, SUB_103_U23, SUB_103_U24, SUB_103_U25, GT_218_U6, GT_218_U7, GT_218_U8, GT_160_U6, GT_160_U7, GT_160_U8, GT_160_U9, GT_206_U6, GT_206_U7, SUB_110_U6, SUB_110_U7, SUB_110_U8, SUB_110_U9, SUB_110_U10, SUB_110_U11, SUB_110_U12, SUB_110_U13, SUB_110_U14, SUB_110_U15, SUB_110_U16, SUB_110_U17, SUB_110_U18, SUB_110_U19, SUB_110_U20, SUB_110_U21, SUB_110_U22, SUB_110_U23, SUB_110_U24, SUB_110_U25, SUB_110_U26, SUB_110_U27, SUB_110_U28, SUB_110_U29, SUB_110_U30, SUB_110_U31, SUB_110_U32, SUB_110_U33, SUB_110_U34, GT_146_U6, GT_146_U7, GT_146_U8, GT_146_U9, GT_126_U6, GT_126_U7, GT_126_U8, GT_163_U6, GT_163_U7, GT_184_U6, GT_184_U7, GT_184_U8, GT_221_U6, GT_221_U7, GT_221_U8, GT_221_U9, GT_227_U6, GT_227_U7, GT_227_U8, ADD_283_U5, ADD_283_U6, ADD_283_U7, ADD_283_U8, ADD_283_U9, ADD_283_U10, ADD_283_U11, ADD_283_U12, ADD_283_U13, ADD_283_U14, ADD_283_U15, ADD_283_U16, ADD_283_U17, ADD_283_U18, ADD_283_U19, ADD_283_U20, ADD_283_U21, ADD_283_U22, ADD_283_U23, ADD_283_U24, ADD_283_U25, ADD_283_U26, ADD_283_U27, GT_197_U6, GT_197_U7, GT_197_U8, GT_114_U6, GT_114_U7, GT_114_U8, GT_114_U9, GT_114_U10, GT_114_U11, GT_224_U6, GT_224_U7, GT_224_U8, ADD_304_U5, ADD_304_U6, ADD_304_U7, ADD_304_U8, ADD_304_U9, ADD_304_U10, ADD_304_U11, ADD_304_U12, ADD_304_U13, ADD_304_U14, ADD_304_U15, ADD_304_U16, ADD_304_U17, ADD_304_U18, ADD_304_U19, ADD_304_U20, ADD_304_U21, ADD_304_U22, ADD_304_U23, ADD_304_U24, ADD_304_U25, ADD_304_U26, ADD_304_U27, R794_U6, R794_U7, R794_U8, R794_U9, R794_U10, R794_U11, R794_U12, R794_U13, R794_U14, R794_U15, R794_U16, R794_U17, R794_U18, R794_U19, R794_U20, R794_U21, R794_U22, R794_U23, R794_U24, R794_U25, R794_U26, R794_U27, R794_U28, R794_U29, R794_U30, R794_U31, R794_U32, R794_U33, R794_U34, R794_U35, R794_U36, R794_U37, R794_U38, R794_U39, R794_U40, R794_U41, R794_U42, R794_U43, R794_U44, R794_U45, R794_U46, R794_U47, R794_U48, R794_U49, R794_U50, R794_U51, R794_U52, R794_U53, R794_U54, R794_U55, R794_U56, R794_U57, R794_U58, R794_U59, R794_U60, R794_U61, R794_U62, R794_U63, R794_U64, R794_U65, R794_U66, R794_U67, R794_U68, R794_U69, R794_U70, R794_U71, R794_U72, R794_U73, R794_U74, R794_U75, R794_U76, R794_U77, R794_U78, R794_U79, R794_U80, R794_U81, R794_U82, R794_U83, R794_U84, R794_U85, R794_U86, R794_U87, R794_U88, R794_U89, R794_U90, R794_U91, GT_130_U6, GT_130_U7, GT_130_U8, GT_130_U9, GT_175_U6, GT_175_U7, GT_175_U8, GT_142_U6, GT_142_U7, GT_142_U8, GT_142_U9, GT_172_U6, GT_172_U7, GT_172_U8, GT_172_U9, GT_172_U10, GT_203_U6, GT_203_U7, GT_203_U8, GT_203_U9, GT_134_U6, GT_134_U7, GT_134_U8, GT_134_U9, SUB_60_U6, SUB_60_U7, SUB_60_U8, SUB_60_U9, SUB_60_U10, SUB_60_U11, SUB_60_U12, SUB_60_U13, SUB_60_U14, SUB_60_U15, SUB_60_U16, SUB_60_U17, SUB_60_U18, SUB_60_U19, SUB_60_U20, SUB_60_U21, SUB_60_U22, SUB_60_U23, SUB_60_U24, SUB_60_U25, SUB_60_U26, SUB_60_U27, SUB_60_U28, SUB_60_U29, SUB_60_U30, SUB_60_U31, SUB_60_U32, SUB_60_U33, SUB_60_U34, SUB_60_U35, SUB_60_U36, SUB_60_U37, SUB_60_U38, SUB_60_U39, SUB_60_U40, SUB_60_U41, SUB_60_U42, SUB_60_U43, SUB_60_U44, SUB_60_U45, SUB_60_U46, SUB_60_U47, SUB_60_U48, SUB_60_U49, SUB_60_U50, SUB_60_U51, SUB_60_U52, SUB_60_U53, SUB_60_U54, SUB_60_U55, SUB_60_U56, SUB_60_U57, SUB_60_U58, SUB_60_U59, SUB_60_U60, SUB_60_U61, SUB_60_U62, SUB_60_U63, SUB_60_U64, SUB_60_U65, SUB_60_U66, SUB_60_U67, SUB_60_U68, SUB_60_U69, SUB_60_U70, SUB_60_U71, SUB_60_U72, SUB_60_U73, SUB_60_U74, SUB_60_U75, SUB_60_U76, SUB_60_U77, SUB_60_U78, SUB_60_U79, SUB_60_U80, SUB_60_U81, SUB_60_U82, SUB_60_U83, SUB_60_U84, SUB_60_U85, SUB_60_U86, SUB_60_U87, SUB_60_U88, SUB_60_U89, SUB_60_U90, SUB_60_U91, SUB_60_U92, SUB_60_U93, SUB_60_U94, SUB_60_U95, SUB_60_U96, SUB_60_U97, SUB_60_U98, SUB_60_U99, SUB_60_U100, SUB_60_U101, SUB_60_U102, SUB_60_U103, SUB_60_U104, SUB_60_U105, SUB_60_U106, SUB_60_U107, SUB_60_U108, SUB_60_U109, SUB_60_U110, SUB_60_U111, SUB_60_U112, SUB_60_U113, SUB_60_U114, SUB_60_U115, SUB_60_U116, SUB_60_U117, SUB_60_U118, SUB_60_U119, SUB_60_U120, GT_181_U6, GT_181_U7, GT_181_U8, SUB_73_U6, SUB_73_U7, SUB_73_U8, SUB_73_U9, SUB_73_U10, SUB_73_U11, SUB_73_U12, SUB_73_U13, SUB_73_U14, SUB_73_U15, SUB_73_U16, SUB_73_U17, SUB_73_U18, SUB_73_U19, SUB_73_U20, SUB_73_U21, SUB_73_U22, SUB_73_U23, SUB_73_U24, SUB_73_U25, SUB_73_U26, SUB_73_U27, SUB_73_U28, SUB_73_U29, SUB_73_U30, SUB_73_U31, SUB_73_U32, SUB_73_U33, SUB_73_U34, SUB_73_U35, SUB_73_U36, SUB_73_U37, SUB_73_U38, SUB_73_U39, SUB_73_U40, SUB_73_U41, SUB_73_U42, SUB_73_U43, SUB_73_U44, SUB_73_U45, SUB_73_U46, SUB_73_U47, SUB_73_U48, SUB_73_U49, SUB_73_U50, SUB_73_U51, SUB_73_U52, SUB_73_U53, SUB_73_U54, SUB_73_U55, SUB_73_U56, SUB_73_U57, SUB_73_U58, GT_212_U6, GT_212_U7, GT_212_U8, GT_212_U9, GT_108_U6, GT_108_U7, GT_108_U8, GT_108_U9, GT_122_U6, GT_122_U7, GT_122_U8, GT_122_U9, GT_122_U10, GT_169_U6, GT_169_U7, GT_169_U8, GT_169_U9, GT_178_U6, GT_178_U7, GT_178_U8, GT_178_U9, SUB_199_U6, SUB_199_U7, SUB_199_U8, SUB_199_U9, SUB_199_U10, SUB_199_U11, SUB_199_U12, SUB_199_U13, SUB_199_U14, SUB_199_U15, SUB_199_U16, SUB_199_U17, SUB_199_U18, SUB_199_U19, SUB_199_U20, GT_209_U6, GT_209_U7, GT_209_U8, GT_209_U9, GT_215_U6, GT_215_U7, GT_215_U8, GT_215_U9, GT_215_U10, GT_166_U6, GT_166_U7, GT_166_U8; 
assign U595 = ~(MAR_REG_3__SCAN_IN | MAR_REG_1__SCAN_IN); 
assign U596 = ~(MAR_REG_4__SCAN_IN | MAR_REG_0__SCAN_IN); 
assign U681 = ~STATO_REG_1__SCAN_IN; 
assign U682 = ~STATO_REG_0__SCAN_IN; 
assign U684 = ~FLAG_REG_SCAN_IN; 
assign U686 = ~STATO_REG_2__SCAN_IN; 
assign U687 = ~MAR_REG_2__SCAN_IN; 
assign U688 = ~MAR_REG_0__SCAN_IN; 
assign U689 = ~MAR_REG_4__SCAN_IN; 
assign U690 = ~MAR_REG_3__SCAN_IN; 
assign U691 = ~MAR_REG_1__SCAN_IN; 
assign U692 = ~(MAR_REG_3__SCAN_IN & MAR_REG_1__SCAN_IN); 
assign U693 = ~(MAR_REG_4__SCAN_IN & MAR_REG_2__SCAN_IN & MAR_REG_0__SCAN_IN); 
assign U694 = ~START; 
assign U705 = ~EN_DISP_REG_SCAN_IN; 
assign U708 = ~MAX_REG_8__SCAN_IN; 
assign U791 = EN_DISP_REG_SCAN_IN | RES_DISP_REG_SCAN_IN; 
assign U800 = START | STATO_REG_1__SCAN_IN; 
assign U869 = STATO_REG_0__SCAN_IN | STATO_REG_1__SCAN_IN | STATO_REG_2__SCAN_IN; 
assign U882 = ~(STATO_REG_0__SCAN_IN & STATO_REG_1__SCAN_IN); 
assign U885 = STATO_REG_0__SCAN_IN | STATO_REG_2__SCAN_IN; 
assign U1021 = ~(MAX_REG_8__SCAN_IN & MAX_REG_0__SCAN_IN); 
assign SUB_103_U9 = MAX_REG_2__SCAN_IN | MAX_REG_1__SCAN_IN | MAX_REG_0__SCAN_IN; 
assign SUB_103_U11 = ~MAX_REG_3__SCAN_IN; 
assign SUB_103_U13 = ~MAX_REG_4__SCAN_IN; 
assign SUB_103_U15 = ~MAX_REG_1__SCAN_IN; 
assign SUB_103_U16 = ~MAX_REG_0__SCAN_IN; 
assign SUB_103_U20 = MAX_REG_1__SCAN_IN | MAX_REG_0__SCAN_IN; 
assign ADD_283_U5 = ~NUM_REG_0__SCAN_IN; 
assign ADD_283_U6 = ~NUM_REG_1__SCAN_IN; 
assign ADD_283_U7 = ~(NUM_REG_1__SCAN_IN & NUM_REG_0__SCAN_IN); 
assign ADD_283_U8 = ~NUM_REG_2__SCAN_IN; 
assign ADD_283_U10 = ~NUM_REG_3__SCAN_IN; 
assign ADD_283_U15 = ~NUM_REG_4__SCAN_IN; 
assign GT_197_U8 = NUM_REG_2__SCAN_IN | NUM_REG_1__SCAN_IN; 
assign ADD_304_U5 = ~MAR_REG_0__SCAN_IN; 
assign ADD_304_U6 = ~MAR_REG_1__SCAN_IN; 
assign ADD_304_U7 = ~(MAR_REG_1__SCAN_IN & MAR_REG_0__SCAN_IN); 
assign ADD_304_U8 = ~MAR_REG_2__SCAN_IN; 
assign ADD_304_U10 = ~MAR_REG_3__SCAN_IN; 
assign ADD_304_U15 = ~MAR_REG_4__SCAN_IN; 
assign SUB_60_U8 = ~TEMP_REG_0__SCAN_IN; 
assign SUB_60_U11 = ~TEMP_REG_2__SCAN_IN; 
assign SUB_60_U13 = ~TEMP_REG_3__SCAN_IN; 
assign SUB_60_U15 = ~TEMP_REG_4__SCAN_IN; 
assign SUB_60_U17 = ~TEMP_REG_5__SCAN_IN; 
assign SUB_60_U19 = ~TEMP_REG_6__SCAN_IN; 
assign SUB_60_U21 = ~TEMP_REG_7__SCAN_IN; 
assign SUB_60_U39 = ~TEMP_REG_8__SCAN_IN; 
assign SUB_60_U46 = ~TEMP_REG_1__SCAN_IN; 
assign SUB_73_U7 = ~MAX_REG_6__SCAN_IN; 
assign SUB_73_U9 = ~MAX_REG_1__SCAN_IN; 
assign SUB_73_U12 = ~MAX_REG_2__SCAN_IN; 
assign SUB_73_U13 = ~MAX_REG_3__SCAN_IN; 
assign SUB_73_U16 = ~MAX_REG_4__SCAN_IN; 
assign SUB_73_U17 = ~MAX_REG_5__SCAN_IN; 
assign SUB_73_U19 = ~MAX_REG_7__SCAN_IN; 
assign SUB_73_U22 = ~MAX_REG_8__SCAN_IN; 
assign SUB_199_U7 = ~NUM_REG_1__SCAN_IN; 
assign SUB_199_U10 = ~NUM_REG_4__SCAN_IN; 
assign SUB_199_U11 = ~NUM_REG_2__SCAN_IN; 
assign SUB_199_U15 = NUM_REG_2__SCAN_IN | NUM_REG_1__SCAN_IN; 
assign SUB_199_U18 = NUM_REG_3__SCAN_IN | NUM_REG_2__SCAN_IN | NUM_REG_1__SCAN_IN; 
assign U589 = U705 & RES_DISP_REG_SCAN_IN; 
assign U597 = U688 & MAR_REG_4__SCAN_IN; 
assign U599 = U690 & MAR_REG_1__SCAN_IN; 
assign U601 = U596 & U687; 
assign U695 = ~(U687 & U689 & MAR_REG_0__SCAN_IN); 
assign U696 = ~(U596 & MAR_REG_2__SCAN_IN); 
assign U697 = ~(U687 & MAR_REG_4__SCAN_IN & MAR_REG_0__SCAN_IN); 
assign U698 = ~(U691 & MAR_REG_3__SCAN_IN); 
assign U700 = ~(U689 & MAR_REG_2__SCAN_IN & MAR_REG_0__SCAN_IN); 
assign U792 = ~U791; 
assign U793 = ~(U681 & START & STATO_REG_0__SCAN_IN); 
assign U799 = ~(U682 & STATO_REG_1__SCAN_IN); 
assign U802 = ~(U684 & STATO_REG_1__SCAN_IN); 
assign U814 = ~U693; 
assign U815 = ~U692; 
assign U825 = ~(ADD_304_U5 & STATO_REG_2__SCAN_IN); 
assign U865 = ~(U686 & STATO_REG_1__SCAN_IN); 
assign U870 = ~(U869 & RES_DISP_REG_SCAN_IN); 
assign U886 = ~(U705 & MAX_REG_8__SCAN_IN); 
assign U958 = ~(U681 & TEMP_REG_8__SCAN_IN); 
assign U960 = ~(U681 & TEMP_REG_7__SCAN_IN); 
assign U962 = ~(U681 & TEMP_REG_6__SCAN_IN); 
assign U964 = ~(U681 & TEMP_REG_5__SCAN_IN); 
assign U966 = ~(U681 & TEMP_REG_4__SCAN_IN); 
assign U968 = ~(U681 & TEMP_REG_3__SCAN_IN); 
assign U970 = ~(U681 & TEMP_REG_2__SCAN_IN); 
assign U972 = ~(U681 & TEMP_REG_1__SCAN_IN); 
assign U974 = ~(U681 & TEMP_REG_0__SCAN_IN); 
assign U1004 = ~(U708 & MAX_REG_4__SCAN_IN); 
assign U1008 = ~(U708 & MAX_REG_3__SCAN_IN); 
assign U1012 = ~(U708 & MAX_REG_2__SCAN_IN); 
assign U1016 = ~(U708 & MAX_REG_1__SCAN_IN); 
assign U1020 = ~(U708 & MAX_REG_0__SCAN_IN); 
assign SUB_103_U17 = ~SUB_103_U9; 
assign SUB_103_U19 = ~(SUB_103_U9 & MAX_REG_3__SCAN_IN); 
assign SUB_103_U21 = ~(SUB_103_U20 & MAX_REG_2__SCAN_IN); 
assign SUB_103_U24 = ~(SUB_103_U16 & MAX_REG_1__SCAN_IN); 
assign SUB_103_U25 = ~(SUB_103_U15 & MAX_REG_0__SCAN_IN); 
assign ADD_283_U17 = ~ADD_283_U7; 
assign ADD_283_U24 = ~(ADD_283_U7 & NUM_REG_2__SCAN_IN); 
assign ADD_283_U26 = ~(ADD_283_U5 & NUM_REG_1__SCAN_IN); 
assign ADD_283_U27 = ~(ADD_283_U6 & NUM_REG_0__SCAN_IN); 
assign GT_197_U7 = GT_197_U8 & NUM_REG_3__SCAN_IN; 
assign ADD_304_U17 = ~ADD_304_U7; 
assign ADD_304_U24 = ~(ADD_304_U7 & MAR_REG_2__SCAN_IN); 
assign ADD_304_U26 = ~(ADD_304_U5 & MAR_REG_1__SCAN_IN); 
assign ADD_304_U27 = ~(ADD_304_U6 & MAR_REG_0__SCAN_IN); 
assign SUB_199_U9 = ~(SUB_199_U15 & NUM_REG_3__SCAN_IN); 
assign SUB_199_U19 = ~(SUB_199_U7 & NUM_REG_2__SCAN_IN); 
assign SUB_199_U20 = ~(SUB_199_U11 & NUM_REG_1__SCAN_IN); 
assign U646 = ~(U791 & U886); 
assign U669 = ~(U793 & U870); 
assign U699 = ~(U597 & U687); 
assign U701 = ~(U597 & MAR_REG_2__SCAN_IN); 
assign U703 = ~(U814 & U815); 
assign U758 = ~(U1021 & U1020); 
assign U827 = ~U695; 
assign U829 = ~U696; 
assign U831 = ~U697; 
assign U833 = ~U698; 
assign U837 = ~U700; 
assign U848 = ~(U692 & U698); 
assign U852 = ~(U595 & U814); 
assign U854 = ~(U700 & U693); 
assign U858 = ~(U601 & U595); 
assign U860 = ~(U599 & U814); 
assign SUB_103_U6 = SUB_103_U21 & SUB_103_U9; 
assign SUB_103_U10 = ~(SUB_103_U17 & SUB_103_U11); 
assign SUB_103_U12 = ~(SUB_103_U25 & SUB_103_U24); 
assign ADD_283_U9 = ~(ADD_283_U17 & NUM_REG_2__SCAN_IN); 
assign ADD_283_U14 = ~(ADD_283_U27 & ADD_283_U26); 
assign ADD_283_U25 = ~(ADD_283_U17 & ADD_283_U8); 
assign GT_197_U6 = GT_197_U7 | NUM_REG_4__SCAN_IN; 
assign ADD_304_U9 = ~(ADD_304_U17 & MAR_REG_2__SCAN_IN); 
assign ADD_304_U14 = ~(ADD_304_U27 & ADD_304_U26); 
assign ADD_304_U25 = ~(ADD_304_U17 & ADD_304_U8); 
assign SUB_199_U6 = SUB_199_U18 & SUB_199_U9; 
assign SUB_199_U12 = SUB_199_U20 & SUB_199_U19; 
assign SUB_199_U13 = ~(SUB_199_U9 & SUB_199_U10); 
assign SUB_199_U16 = ~SUB_199_U9; 
assign U706 = ~GT_197_U6; 
assign U795 = ~(U601 & U848); 
assign U796 = ~(U703 & STATO_REG_2__SCAN_IN); 
assign U816 = ~U703; 
assign U823 = ~(ADD_304_U14 & STATO_REG_2__SCAN_IN); 
assign U828 = ~(U827 & U815); 
assign U830 = ~(U595 & U829); 
assign U832 = ~(U831 & U815); 
assign U834 = ~(U833 & U831); 
assign U835 = ~U699; 
assign U838 = ~(U837 & U815); 
assign U840 = ~(U696 & U695 & U699); 
assign U841 = ~U701; 
assign U842 = ~(U697 & U701); 
assign U845 = ~(U833 & U827); 
assign U846 = ~(U599 & U831); 
assign U847 = ~(U599 & U837); 
assign U851 = ~(U837 & U595); 
assign U853 = ~(U595 & U827); 
assign U855 = ~(U833 & U854); 
assign U856 = ~(U701 & U696); 
assign U873 = ~(U833 & MAR_REG_2__SCAN_IN & MAR_REG_0__SCAN_IN); 
assign U997 = ~(SUB_199_U6 & GT_197_U6); 
assign U999 = ~(SUB_199_U12 & GT_197_U6); 
assign U1001 = ~(SUB_199_U7 & GT_197_U6); 
assign U1003 = ~(GT_197_U6 & NUM_REG_0__SCAN_IN); 
assign U1013 = ~(SUB_103_U6 & MAX_REG_8__SCAN_IN); 
assign U1017 = ~(SUB_103_U12 & MAX_REG_8__SCAN_IN); 
assign SUB_103_U7 = SUB_103_U19 & SUB_103_U10; 
assign SUB_103_U18 = ~SUB_103_U10; 
assign SUB_103_U22 = ~(SUB_103_U10 & MAX_REG_4__SCAN_IN); 
assign ADD_283_U13 = ~(ADD_283_U25 & ADD_283_U24); 
assign ADD_283_U18 = ~ADD_283_U9; 
assign ADD_283_U22 = ~(ADD_283_U9 & NUM_REG_3__SCAN_IN); 
assign ADD_304_U13 = ~(ADD_304_U25 & ADD_304_U24); 
assign ADD_304_U18 = ~ADD_304_U9; 
assign ADD_304_U22 = ~(ADD_304_U9 & MAR_REG_3__SCAN_IN); 
assign SUB_199_U14 = ~SUB_199_U13; 
assign SUB_199_U17 = ~(SUB_199_U16 & NUM_REG_4__SCAN_IN); 
assign U588 = GT_197_U6 & SUB_199_U14; 
assign U591 = U589 & U706; 
assign U594 = U793 & U796; 
assign U704 = ~(U816 & STATO_REG_2__SCAN_IN); 
assign U754 = ~(U1013 & U1012); 
assign U756 = ~(U1017 & U1016); 
assign U821 = ~(ADD_304_U13 & STATO_REG_2__SCAN_IN); 
assign U836 = ~(U835 & U595); 
assign U843 = ~(U595 & U842); 
assign U844 = ~(U599 & U840); 
assign U849 = ~(U841 & U599); 
assign U850 = ~(U835 & U833); 
assign U857 = ~(U815 & U856); 
assign U866 = ~(U865 & U682 & U796); 
assign U994 = ~(U706 & NUM_REG_4__SCAN_IN); 
assign U996 = ~(U706 & NUM_REG_3__SCAN_IN); 
assign U998 = ~(U706 & NUM_REG_2__SCAN_IN); 
assign U1000 = ~(U706 & NUM_REG_1__SCAN_IN); 
assign U1002 = ~(U706 & NUM_REG_0__SCAN_IN); 
assign U1009 = ~(SUB_103_U7 & MAX_REG_8__SCAN_IN); 
assign SUB_103_U8 = ~(SUB_103_U18 & SUB_103_U13); 
assign SUB_103_U23 = ~(SUB_103_U18 & SUB_103_U13); 
assign ADD_283_U16 = ~(ADD_283_U18 & NUM_REG_3__SCAN_IN); 
assign ADD_283_U23 = ~(ADD_283_U18 & ADD_283_U10); 
assign ADD_304_U16 = ~(ADD_304_U18 & MAR_REG_3__SCAN_IN); 
assign ADD_304_U23 = ~(ADD_304_U18 & ADD_304_U10); 
assign SUB_199_U8 = ~(SUB_199_U13 & SUB_199_U17); 
assign U587 = SUB_103_U8 & MAX_REG_8__SCAN_IN; 
assign U598 = U838 & U836 & U834 & U832; 
assign U600 = U845 & U843 & U844; 
assign U602 = U851 & U850; 
assign U604 = U853 & U849 & U836 & U832; 
assign U606 = U830 & U795 & U703 & U858 & U857; 
assign U608 = U849 & U847 & U846 & U828; 
assign U644 = ~(U594 & U799); 
assign U746 = ~(U997 & U996); 
assign U747 = ~(U999 & U998); 
assign U748 = ~(U1001 & U1000); 
assign U749 = ~(U1003 & U1002); 
assign U752 = ~(U1009 & U1008); 
assign U797 = ~U704; 
assign U818 = ~(U594 & MAR_REG_4__SCAN_IN); 
assign U820 = ~(U594 & MAR_REG_3__SCAN_IN); 
assign U822 = ~(U594 & MAR_REG_2__SCAN_IN); 
assign U824 = ~(U594 & MAR_REG_1__SCAN_IN); 
assign U826 = ~(U594 & MAR_REG_0__SCAN_IN); 
assign U868 = ~(U866 & EN_DISP_REG_SCAN_IN); 
assign U883 = ~(U704 & STATO_REG_1__SCAN_IN); 
assign U995 = ~(SUB_199_U8 & GT_197_U6); 
assign SUB_103_U14 = SUB_103_U23 & SUB_103_U22; 
assign SUB_110_U7 = ~U754; 
assign ADD_283_U12 = ~(ADD_283_U23 & ADD_283_U22); 
assign ADD_283_U19 = ~ADD_283_U16; 
assign ADD_283_U20 = ~(ADD_283_U16 & NUM_REG_4__SCAN_IN); 
assign ADD_304_U12 = ~(ADD_304_U23 & ADD_304_U22); 
assign ADD_304_U19 = ~ADD_304_U16; 
assign ADD_304_U20 = ~(ADD_304_U16 & MAR_REG_4__SCAN_IN); 
assign U603 = U600 & U852; 
assign U605 = U604 & U855; 
assign U609 = U602 & U860 & U834 & U795; 
assign U610 = U604 & U873; 
assign U624 = ~(U830 & U828 & U598); 
assign U625 = ~(U608 & U602 & U600 & U838); 
assign U626 = ~(U860 & U846 & U598 & U606 & U602); 
assign U629 = ~(U608 & U606); 
assign U671 = ~(U826 & U825); 
assign U672 = ~(U824 & U823); 
assign U673 = ~(U822 & U821); 
assign U745 = ~(U995 & U994); 
assign U819 = ~(ADD_304_U12 & STATO_REG_2__SCAN_IN); 
assign U867 = ~(U797 & STATO_REG_0__SCAN_IN); 
assign U881 = ~(U797 & START); 
assign U884 = ~(U883 & U694); 
assign U1005 = ~(SUB_103_U14 & MAX_REG_8__SCAN_IN); 
assign SUB_110_U9 = U754 | U752; 
assign SUB_110_U10 = ~U587; 
assign SUB_110_U26 = ~(U752 & U754); 
assign GT_221_U7 = U749 & U748; 
assign GT_227_U8 = U748 | U588 | U588 | U749; 
assign ADD_283_U21 = ~(ADD_283_U19 & ADD_283_U15); 
assign GT_224_U8 = U748 | U588 | U588 | U588; 
assign ADD_304_U21 = ~(ADD_304_U19 & ADD_304_U15); 
assign GT_203_U9 = U747 | U749 | U748; 
assign GT_212_U7 = U747 & U748; 
assign GT_209_U7 = U748 & U747 & U749; 
assign GT_215_U10 = U749 | U748; 
assign U607 = U838 & U828 & U847 & U606 & U603; 
assign U627 = ~(U834 & U830 & U836 & U608 & U603); 
assign U628 = ~(U610 & U609); 
assign U643 = ~(U882 & U881); 
assign U645 = ~(U799 & U885 & U796 & U884); 
assign U670 = ~(U868 & U793 & U867); 
assign U674 = ~(U820 & U819); 
assign U750 = ~(U1005 & U1004); 
assign U839 = ~U624; 
assign U861 = ~(U609 & U605); 
assign U959 = ~(U624 & STATO_REG_1__SCAN_IN); 
assign U967 = ~(U629 & STATO_REG_1__SCAN_IN); 
assign U973 = ~(U626 & STATO_REG_1__SCAN_IN); 
assign U975 = ~(U625 & STATO_REG_1__SCAN_IN); 
assign GT_218_U8 = U588 | U588 | U745; 
assign GT_206_U7 = ~(U588 | U746 | U745 | U588 | U588); 
assign SUB_110_U6 = ~(SUB_110_U9 & SUB_110_U26); 
assign SUB_110_U20 = ~SUB_110_U9; 
assign GT_221_U9 = U746 | U745 | U588 | U588; 
assign GT_227_U6 = ~(GT_227_U8 | U588 | U747 | U746 | U745); 
assign ADD_283_U11 = ~(ADD_283_U21 & ADD_283_U20); 
assign GT_224_U7 = ~(GT_224_U8 | U745 | U747 | U746); 
assign ADD_304_U11 = ~(ADD_304_U21 & ADD_304_U20); 
assign GT_203_U7 = U746 & GT_203_U9; 
assign SUB_60_U10 = ~U626; 
assign SUB_60_U16 = ~U629; 
assign SUB_60_U24 = ~U625; 
assign SUB_60_U40 = ~U624; 
assign SUB_60_U62 = ~(U629 & SUB_60_U15); 
assign SUB_60_U80 = ~(U625 & SUB_60_U8); 
assign SUB_60_U82 = ~(U624 & SUB_60_U39); 
assign SUB_60_U84 = ~(U624 & SUB_60_U39); 
assign SUB_60_U102 = ~(U629 & SUB_60_U15); 
assign SUB_60_U117 = ~(U626 & SUB_60_U46); 
assign SUB_73_U10 = ~U626; 
assign SUB_73_U14 = ~U629; 
assign SUB_73_U23 = ~U624; 
assign SUB_73_U24 = ~U625; 
assign SUB_73_U29 = ~(U626 & SUB_73_U9); 
assign SUB_73_U35 = ~(U629 & SUB_73_U16); 
assign SUB_73_U55 = ~(U624 & SUB_73_U22); 
assign SUB_73_U57 = ~(U624 & SUB_73_U22); 
assign GT_212_U9 = U588 | U588 | U745; 
assign GT_209_U9 = U588 | U746 | U745; 
assign GT_215_U7 = U747 & GT_215_U10; 
assign GT_215_U9 = U588 | U746 | U745; 
assign U630 = ~(U610 & U607); 
assign U631 = ~(U602 & U603 & U849 & U839); 
assign U632 = ~(U795 & U846 & U839 & U600 & U847); 
assign U727 = ~(U959 & U958); 
assign U731 = ~(U967 & U966); 
assign U734 = ~(U973 & U972); 
assign U735 = ~(U975 & U974); 
assign U817 = ~(ADD_304_U11 & STATO_REG_2__SCAN_IN); 
assign U859 = ~(U605 & U607); 
assign U969 = ~(U861 & STATO_REG_1__SCAN_IN); 
assign U971 = ~(U627 & STATO_REG_1__SCAN_IN); 
assign GT_218_U7 = ~(GT_218_U8 | U747 | U746 | U588); 
assign GT_206_U6 = ~(U588 | GT_206_U7); 
assign SUB_110_U12 = ~U750; 
assign SUB_110_U25 = ~(U750 & SUB_110_U9); 
assign GT_221_U8 = ~(GT_221_U9 | GT_221_U7 | U588 | U747); 
assign GT_227_U7 = ~(GT_227_U6 | U588); 
assign GT_224_U6 = ~(U588 | GT_224_U7); 
assign GT_203_U8 = ~(U588 | GT_203_U7 | U745 | U588 | U588); 
assign SUB_60_U9 = ~(SUB_60_U24 & TEMP_REG_0__SCAN_IN); 
assign SUB_60_U12 = ~U627; 
assign SUB_60_U14 = ~U628; 
assign SUB_60_U54 = ~(U627 & SUB_60_U11); 
assign SUB_60_U58 = ~(U628 & SUB_60_U13); 
assign SUB_60_U60 = ~(SUB_60_U16 & TEMP_REG_4__SCAN_IN); 
assign SUB_60_U81 = ~(SUB_60_U40 & TEMP_REG_8__SCAN_IN); 
assign SUB_60_U83 = ~(SUB_60_U40 & TEMP_REG_8__SCAN_IN); 
assign SUB_60_U101 = ~(SUB_60_U16 & TEMP_REG_4__SCAN_IN); 
assign SUB_60_U107 = ~(U628 & SUB_60_U13); 
assign SUB_60_U112 = ~(U627 & SUB_60_U11); 
assign SUB_60_U116 = ~(SUB_60_U10 & TEMP_REG_1__SCAN_IN); 
assign SUB_73_U11 = ~U627; 
assign SUB_73_U15 = ~U628; 
assign SUB_73_U26 = ~(SUB_73_U10 & MAX_REG_1__SCAN_IN); 
assign SUB_73_U27 = ~(SUB_73_U24 & MAX_REG_0__SCAN_IN); 
assign SUB_73_U30 = ~(U627 & SUB_73_U12); 
assign SUB_73_U36 = ~(U628 & SUB_73_U13); 
assign SUB_73_U38 = ~(SUB_73_U14 & MAX_REG_4__SCAN_IN); 
assign SUB_73_U54 = ~(SUB_73_U23 & MAX_REG_8__SCAN_IN); 
assign SUB_73_U56 = ~(SUB_73_U23 & MAX_REG_8__SCAN_IN); 
assign GT_212_U8 = ~(GT_212_U9 | GT_212_U7 | U588 | U746); 
assign GT_108_U9 = U754 | U752 | U750; 
assign GT_209_U8 = ~(GT_209_U9 | GT_209_U7 | U588 | U588); 
assign GT_215_U8 = ~(GT_215_U9 | GT_215_U7 | U588 | U588); 
assign U675 = ~(U818 & U817); 
assign U714 = ~GT_224_U6; 
assign U732 = ~(U969 & U968); 
assign U733 = ~(U971 & U970); 
assign U789 = ~GT_206_U6; 
assign U903 = GT_224_U6 | GT_227_U7; 
assign U961 = ~(U632 & STATO_REG_1__SCAN_IN); 
assign U963 = ~(U631 & STATO_REG_1__SCAN_IN); 
assign U965 = ~(U859 & STATO_REG_1__SCAN_IN); 
assign GT_218_U6 = ~(U588 | GT_218_U7); 
assign SUB_110_U18 = ~(SUB_110_U20 & SUB_110_U12); 
assign GT_221_U6 = ~(U588 | GT_221_U8); 
assign GT_203_U6 = ~(U588 | GT_203_U8); 
assign SUB_60_U7 = ~(SUB_60_U9 & SUB_60_U80); 
assign SUB_60_U18 = ~U630; 
assign SUB_60_U20 = ~U631; 
assign SUB_60_U22 = ~U632; 
assign SUB_60_U35 = ~(SUB_60_U102 & SUB_60_U101); 
assign SUB_60_U38 = ~(SUB_60_U117 & SUB_60_U116); 
assign SUB_60_U47 = ~SUB_60_U9; 
assign SUB_60_U50 = ~(U626 & SUB_60_U9); 
assign SUB_60_U52 = ~(SUB_60_U12 & TEMP_REG_2__SCAN_IN); 
assign SUB_60_U56 = ~(SUB_60_U14 & TEMP_REG_3__SCAN_IN); 
assign SUB_60_U66 = ~(U630 & SUB_60_U17); 
assign SUB_60_U70 = ~(U631 & SUB_60_U19); 
assign SUB_60_U72 = ~(U632 & SUB_60_U21); 
assign SUB_60_U78 = ~(U632 & SUB_60_U21); 
assign SUB_60_U85 = ~(SUB_60_U84 & SUB_60_U83); 
assign SUB_60_U87 = ~(U632 & SUB_60_U21); 
assign SUB_60_U92 = ~(U631 & SUB_60_U19); 
assign SUB_60_U97 = ~(U630 & SUB_60_U17); 
assign SUB_60_U106 = ~(SUB_60_U14 & TEMP_REG_3__SCAN_IN); 
assign SUB_60_U111 = ~(SUB_60_U12 & TEMP_REG_2__SCAN_IN); 
assign SUB_73_U8 = ~U630; 
assign SUB_73_U18 = ~U631; 
assign SUB_73_U20 = ~U632; 
assign SUB_73_U28 = ~(SUB_73_U27 & SUB_73_U26); 
assign SUB_73_U32 = ~(SUB_73_U11 & MAX_REG_2__SCAN_IN); 
assign SUB_73_U33 = ~(SUB_73_U15 & MAX_REG_3__SCAN_IN); 
assign SUB_73_U41 = ~(U630 & SUB_73_U17); 
assign SUB_73_U44 = ~(U631 & SUB_73_U7); 
assign SUB_73_U46 = ~(U632 & SUB_73_U19); 
assign SUB_73_U52 = ~(U632 & SUB_73_U19); 
assign SUB_73_U58 = ~(SUB_73_U57 & SUB_73_U56); 
assign GT_212_U6 = ~(U588 | GT_212_U8); 
assign GT_108_U7 = U587 & U587 & GT_108_U9; 
assign GT_209_U6 = ~(U588 | GT_209_U8); 
assign GT_215_U6 = ~(U588 | GT_215_U8); 
assign U613 = ~(GT_206_U6 | GT_203_U6); 
assign U711 = ~GT_218_U6; 
assign U712 = ~(GT_227_U7 & U714); 
assign U713 = GT_212_U6 | GT_215_U6; 
assign U728 = ~(U961 & U960); 
assign U729 = ~(U963 & U962); 
assign U730 = ~(U965 & U964); 
assign U776 = ~GT_203_U6; 
assign U780 = ~GT_215_U6; 
assign U782 = ~GT_209_U6; 
assign U783 = ~GT_212_U6; 
assign U790 = ~GT_221_U6; 
assign U890 = GT_221_U6 | GT_224_U6; 
assign U901 = GT_221_U6 | GT_227_U7 | GT_224_U6 | GT_209_U6; 
assign SUB_110_U8 = ~(SUB_110_U18 & SUB_110_U25); 
assign SUB_110_U11 = ~(U587 & SUB_110_U18); 
assign SUB_110_U21 = ~SUB_110_U18; 
assign SUB_110_U33 = ~(U587 & SUB_110_U18); 
assign SUB_60_U36 = ~(SUB_60_U107 & SUB_60_U106); 
assign SUB_60_U37 = ~(SUB_60_U112 & SUB_60_U111); 
assign SUB_60_U48 = ~(SUB_60_U47 & SUB_60_U10); 
assign SUB_60_U64 = ~(SUB_60_U18 & TEMP_REG_5__SCAN_IN); 
assign SUB_60_U68 = ~(SUB_60_U20 & TEMP_REG_6__SCAN_IN); 
assign SUB_60_U74 = ~(SUB_60_U22 & TEMP_REG_7__SCAN_IN); 
assign SUB_60_U76 = ~(SUB_60_U22 & TEMP_REG_7__SCAN_IN); 
assign SUB_60_U86 = ~(SUB_60_U22 & TEMP_REG_7__SCAN_IN); 
assign SUB_60_U91 = ~(SUB_60_U20 & TEMP_REG_6__SCAN_IN); 
assign SUB_60_U96 = ~(SUB_60_U18 & TEMP_REG_5__SCAN_IN); 
assign SUB_60_U103 = ~SUB_60_U35; 
assign SUB_60_U118 = ~SUB_60_U38; 
assign SUB_60_U120 = ~(SUB_60_U38 & SUB_60_U9); 
assign SUB_73_U25 = ~(SUB_73_U18 & MAX_REG_6__SCAN_IN); 
assign SUB_73_U31 = ~(SUB_73_U29 & SUB_73_U28 & SUB_73_U30); 
assign SUB_73_U39 = ~(SUB_73_U8 & MAX_REG_5__SCAN_IN); 
assign SUB_73_U48 = ~(SUB_73_U20 & MAX_REG_7__SCAN_IN); 
assign SUB_73_U50 = ~(SUB_73_U20 & MAX_REG_7__SCAN_IN); 
assign GT_108_U8 = ~(GT_108_U7 | U587); 
assign U887 = ~U713; 
assign U888 = ~(U713 & U782); 
assign U889 = ~(GT_218_U6 & U782); 
assign U891 = ~(U890 & U782); 
assign U893 = ~U712; 
assign U898 = ~(U613 & U782 & U713); 
assign U899 = ~(U790 & U711 & U712); 
assign U904 = ~(U790 & U903); 
assign SUB_110_U22 = ~SUB_110_U11; 
assign SUB_110_U31 = ~(U587 & SUB_110_U11); 
assign SUB_110_U34 = ~(SUB_110_U21 & SUB_110_U10); 
assign SUB_60_U32 = ~(SUB_60_U87 & SUB_60_U86); 
assign SUB_60_U33 = ~(SUB_60_U92 & SUB_60_U91); 
assign SUB_60_U34 = ~(SUB_60_U97 & SUB_60_U96); 
assign SUB_60_U49 = ~(SUB_60_U48 & SUB_60_U46); 
assign SUB_60_U108 = ~SUB_60_U36; 
assign SUB_60_U113 = ~SUB_60_U37; 
assign SUB_60_U119 = ~(SUB_60_U118 & SUB_60_U47); 
assign SUB_73_U34 = ~(SUB_73_U32 & SUB_73_U33 & SUB_73_U31); 
assign GT_108_U6 = ~(U587 | GT_108_U8); 
assign U614 = U613 & U888; 
assign U616 = U613 & U782 & U887; 
assign U657 = U589 & U898; 
assign U707 = ~GT_108_U6; 
assign U894 = ~(U893 & U790); 
assign U905 = ~(U780 & U711 & U904); 
assign U1007 = ~(SUB_110_U8 & GT_108_U6); 
assign U1011 = ~(SUB_110_U6 & GT_108_U6); 
assign U1015 = ~(SUB_110_U7 & GT_108_U6); 
assign U1019 = ~(U756 & GT_108_U6); 
assign U1023 = ~(U758 & GT_108_U6); 
assign SUB_110_U16 = ~(U587 & SUB_110_U22); 
assign SUB_110_U19 = SUB_110_U34 & SUB_110_U33; 
assign SUB_110_U32 = ~(SUB_110_U22 & SUB_110_U10); 
assign SUB_60_U31 = ~(SUB_60_U120 & SUB_60_U119); 
assign SUB_60_U45 = ~(SUB_60_U50 & SUB_60_U49); 
assign SUB_60_U88 = ~SUB_60_U32; 
assign SUB_60_U93 = ~SUB_60_U33; 
assign SUB_60_U98 = ~SUB_60_U34; 
assign SUB_73_U37 = ~(SUB_73_U35 & SUB_73_U36 & SUB_73_U34); 
assign U590 = U589 & U707; 
assign U615 = U614 & U889; 
assign U794 = ~(U587 & U707); 
assign U877 = ~(SUB_110_U19 & GT_108_U6); 
assign U895 = ~(U782 & U711 & U894); 
assign U897 = ~(GT_224_U6 & U711 & U790 & U616); 
assign U900 = ~(U616 & U899); 
assign U906 = ~(U783 & U905); 
assign U1006 = ~(U750 & U707); 
assign U1010 = ~(U752 & U707); 
assign U1014 = ~(U754 & U707); 
assign U1018 = ~(U756 & U707); 
assign U1022 = ~(U758 & U707); 
assign SUB_110_U14 = ~(SUB_110_U32 & SUB_110_U31); 
assign SUB_110_U15 = ~(SUB_110_U10 & SUB_110_U16); 
assign SUB_110_U23 = ~SUB_110_U16; 
assign SUB_110_U29 = ~(U587 & SUB_110_U16); 
assign SUB_60_U51 = ~SUB_60_U45; 
assign SUB_60_U53 = ~(SUB_60_U52 & SUB_60_U45); 
assign SUB_60_U115 = ~(SUB_60_U37 & SUB_60_U45); 
assign SUB_73_U40 = ~(SUB_73_U38 & SUB_73_U39 & SUB_73_U37); 
assign U636 = ~(U794 & U877); 
assign U656 = U589 & U897; 
assign U658 = U589 & U900; 
assign U751 = ~(U1007 & U1006); 
assign U753 = ~(U1011 & U1010); 
assign U755 = ~(U1015 & U1014); 
assign U757 = ~(U1019 & U1018); 
assign U759 = ~(U1023 & U1022); 
assign U876 = ~(SUB_110_U14 & GT_108_U6); 
assign U892 = ~(U891 & U615 & RES_DISP_REG_SCAN_IN); 
assign U896 = ~(U614 & U895); 
assign U902 = ~(U615 & U901); 
assign U907 = ~(U906 & U782); 
assign SUB_110_U24 = ~SUB_110_U15; 
assign SUB_110_U27 = ~(U587 & SUB_110_U15); 
assign SUB_110_U30 = ~(SUB_110_U23 & SUB_110_U10); 
assign SUB_60_U44 = ~(SUB_60_U54 & SUB_60_U53); 
assign SUB_60_U114 = ~(SUB_60_U51 & SUB_60_U113); 
assign SUB_73_U42 = ~(SUB_73_U40 & SUB_73_U41); 
assign U635 = ~(U794 & U876); 
assign U654 = U892 & U705; 
assign U655 = U589 & U896; 
assign U659 = U589 & U902; 
assign U908 = ~(U789 & U907); 
assign GT_138_U7 = U755 & U753 & U751 & U757; 
assign GT_118_U9 = U636 | U751; 
assign SUB_110_U17 = SUB_110_U30 & SUB_110_U29; 
assign SUB_110_U28 = ~(SUB_110_U24 & SUB_110_U10); 
assign GT_146_U9 = U755 | U757; 
assign GT_126_U7 = U636 & U755 & U753 & U751; 
assign GT_114_U10 = U755 | U757; 
assign R794_U9 = ~U755; 
assign R794_U11 = ~U753; 
assign R794_U13 = ~U751; 
assign R794_U15 = ~U636; 
assign R794_U19 = ~U757; 
assign GT_130_U9 = U755 | U753 | U757; 
assign GT_142_U9 = U755 | U753; 
assign GT_134_U9 = U753 | U751; 
assign SUB_60_U30 = ~(SUB_60_U115 & SUB_60_U114); 
assign SUB_60_U55 = ~SUB_60_U44; 
assign SUB_60_U57 = ~(SUB_60_U56 & SUB_60_U44); 
assign SUB_60_U110 = ~(SUB_60_U36 & SUB_60_U44); 
assign SUB_73_U43 = ~(SUB_73_U42 & SUB_73_U25); 
assign GT_122_U7 = U755 & U757; 
assign U660 = U589 & U776 & U908; 
assign U875 = ~(SUB_110_U17 & GT_108_U6); 
assign GT_118_U7 = U635 & GT_118_U9; 
assign SUB_110_U13 = ~(SUB_110_U28 & SUB_110_U27); 
assign GT_146_U7 = U753 & GT_146_U9; 
assign GT_114_U7 = U753 & U751 & GT_114_U10; 
assign R794_U17 = ~U635; 
assign GT_130_U7 = U636 & U751 & GT_130_U9; 
assign GT_142_U7 = U751 & GT_142_U9; 
assign GT_134_U7 = U636 & GT_134_U9; 
assign SUB_60_U43 = ~(SUB_60_U58 & SUB_60_U57); 
assign SUB_60_U109 = ~(SUB_60_U55 & SUB_60_U108); 
assign SUB_73_U21 = ~(SUB_73_U44 & SUB_73_U43); 
assign GT_122_U10 = U753 | GT_122_U7 | U751 | U636; 
assign U634 = ~(U794 & U875); 
assign U874 = ~(GT_108_U6 & SUB_110_U13); 
assign GT_114_U11 = GT_114_U7 | U636; 
assign SUB_60_U29 = ~(SUB_60_U110 & SUB_60_U109); 
assign SUB_60_U59 = ~SUB_60_U43; 
assign SUB_60_U61 = ~(SUB_60_U60 & SUB_60_U43); 
assign SUB_60_U105 = ~(SUB_60_U35 & SUB_60_U43); 
assign SUB_73_U45 = ~SUB_73_U21; 
assign SUB_73_U51 = ~(SUB_73_U50 & SUB_73_U21); 
assign GT_122_U8 = U635 & GT_122_U10; 
assign U633 = ~(U794 & U874); 
assign GT_138_U8 = ~(U634 | U636 | U635 | GT_138_U7); 
assign GT_118_U8 = ~(GT_118_U7 | U634); 
assign GT_146_U8 = ~(U634 | U635 | GT_146_U7 | U636 | U751); 
assign GT_126_U8 = ~(U634 | GT_126_U7 | U635); 
assign GT_114_U8 = U635 & GT_114_U11; 
assign R794_U34 = ~U634; 
assign GT_130_U8 = ~(U634 | GT_130_U7 | U635); 
assign GT_142_U8 = ~(U634 | U635 | U636 | GT_142_U7); 
assign GT_134_U8 = ~(U634 | GT_134_U7 | U635); 
assign SUB_60_U42 = ~(SUB_60_U62 & SUB_60_U61); 
assign SUB_60_U104 = ~(SUB_60_U59 & SUB_60_U103); 
assign SUB_73_U47 = ~(SUB_73_U45 & SUB_73_U46); 
assign SUB_73_U53 = ~(SUB_73_U55 & SUB_73_U54 & SUB_73_U52 & SUB_73_U51); 
assign GT_122_U9 = ~(GT_122_U8 | U634); 
assign GT_138_U6 = ~(U633 | GT_138_U8); 
assign GT_118_U6 = ~(U633 | GT_118_U8); 
assign GT_146_U6 = ~(U633 | GT_146_U8); 
assign GT_126_U6 = ~(U633 | GT_126_U8); 
assign GT_114_U9 = ~(GT_114_U8 | U634); 
assign R794_U32 = ~U633; 
assign GT_130_U6 = ~(U633 | GT_130_U8); 
assign GT_142_U6 = ~(U633 | GT_142_U8); 
assign GT_134_U6 = ~(U633 | GT_134_U8); 
assign SUB_60_U28 = ~(SUB_60_U105 & SUB_60_U104); 
assign SUB_60_U63 = ~SUB_60_U42; 
assign SUB_60_U65 = ~(SUB_60_U64 & SUB_60_U42); 
assign SUB_60_U100 = ~(SUB_60_U34 & SUB_60_U42); 
assign SUB_73_U49 = ~(SUB_73_U48 & SUB_73_U58 & SUB_73_U47); 
assign GT_122_U6 = ~(U633 | GT_122_U9); 
assign U709 = GT_130_U6 | GT_126_U6; 
assign U710 = GT_138_U6 | GT_142_U6 | GT_134_U6; 
assign U719 = ~GT_146_U6; 
assign U721 = ~GT_142_U6; 
assign U722 = ~GT_130_U6; 
assign U723 = ~GT_126_U6; 
assign U724 = ~GT_134_U6; 
assign U725 = ~GT_138_U6; 
assign U726 = ~GT_122_U6; 
assign U774 = ~GT_118_U6; 
assign U941 = GT_138_U6 | GT_142_U6 | GT_146_U6; 
assign U945 = GT_146_U6 | GT_142_U6; 
assign GT_114_U6 = ~(U633 | GT_114_U9); 
assign SUB_60_U41 = ~(SUB_60_U66 & SUB_60_U65); 
assign SUB_60_U99 = ~(SUB_60_U63 & SUB_60_U98); 
assign SUB_73_U6 = ~(SUB_73_U49 & SUB_73_U53); 
assign U611 = ~(GT_114_U6 | GT_118_U6); 
assign U720 = ~(GT_146_U6 & U721); 
assign U778 = ~GT_114_U6; 
assign U879 = ~U710; 
assign U880 = ~U709; 
assign U931 = ~(U709 & U726); 
assign U932 = ~(U710 & U726); 
assign U942 = ~(U724 & U941); 
assign U946 = ~(U725 & U945); 
assign U955 = ~(GT_122_U6 & U774); 
assign SUB_60_U27 = ~(SUB_60_U100 & SUB_60_U99); 
assign SUB_60_U67 = ~SUB_60_U41; 
assign SUB_60_U69 = ~(SUB_60_U68 & SUB_60_U41); 
assign SUB_60_U95 = ~(SUB_60_U33 & SUB_60_U41); 
assign U612 = U880 & U719 & U879; 
assign U621 = U611 & U931; 
assign U637 = ~(U611 & U726); 
assign U934 = ~U720; 
assign U939 = ~(U724 & U725 & U720); 
assign U943 = ~(U942 & U726); 
assign U947 = ~(U724 & U722 & U946); 
assign U953 = ~(U726 & U774 & GT_134_U6 & U880); 
assign U954 = ~(GT_122_U6 & U611); 
assign SUB_60_U23 = ~(SUB_60_U70 & SUB_60_U69); 
assign SUB_60_U94 = ~(SUB_60_U67 & SUB_60_U93); 
assign U772 = ~(U611 & U726 & U612); 
assign U878 = ~U637; 
assign U933 = ~(U621 & U932 & RES_DISP_REG_SCAN_IN); 
assign U935 = ~(U934 & U725); 
assign U944 = ~(U621 & U943); 
assign U948 = ~(U723 & U947); 
assign R794_U16 = ~U637; 
assign R794_U57 = ~(U637 & R794_U17); 
assign R794_U67 = ~(U637 & R794_U17); 
assign SUB_60_U26 = ~(SUB_60_U95 & SUB_60_U94); 
assign SUB_60_U71 = ~SUB_60_U23; 
assign SUB_60_U77 = ~(SUB_60_U76 & SUB_60_U23); 
assign SUB_60_U90 = ~(SUB_60_U32 & SUB_60_U23); 
assign U593 = U880 & U878; 
assign U661 = U933 & U705; 
assign U666 = U589 & U944; 
assign U769 = SUB_60_U31 | SUB_60_U7 | SUB_60_U30 | SUB_60_U29 | SUB_60_U26; 
assign U771 = ~(U612 & U878); 
assign U784 = ~(GT_130_U6 & U723 & U878); 
assign U786 = ~(GT_126_U6 & U878); 
assign U936 = ~(U724 & U726 & U935); 
assign U938 = ~(U709 & U878); 
assign U949 = ~(U948 & U726); 
assign U956 = ~U772; 
assign U1040 = ~(U759 & U772); 
assign R794_U59 = ~(U635 & R794_U16); 
assign R794_U68 = ~(U635 & R794_U16); 
assign SUB_60_U73 = ~(SUB_60_U71 & SUB_60_U72); 
assign SUB_60_U79 = ~(SUB_60_U82 & SUB_60_U81 & SUB_60_U78 & SUB_60_U77); 
assign SUB_60_U89 = ~(SUB_60_U88 & SUB_60_U71); 
assign U664 = U589 & U938; 
assign U785 = ~(U724 & U725 & GT_142_U6 & U593); 
assign U787 = ~(GT_138_U6 & U724 & U593); 
assign U937 = ~(U621 & U936); 
assign U940 = ~(U593 & U939); 
assign U950 = ~(U774 & U949); 
assign U951 = ~(GT_134_U6 & U593); 
assign U952 = ~(U593 & U879); 
assign U957 = ~U771; 
assign U1033 = ~(U956 & U751); 
assign U1035 = ~(U956 & U753); 
assign U1037 = ~(U956 & U755); 
assign U1039 = ~(U956 & U757); 
assign U1041 = ~(U956 & U759); 
assign R794_U27 = ~(R794_U68 & R794_U67); 
assign SUB_60_U25 = ~(SUB_60_U90 & SUB_60_U89); 
assign SUB_60_U75 = ~(SUB_60_U74 & SUB_60_U85 & SUB_60_U73); 
assign U622 = U786 & U785 & U787; 
assign U623 = U787 & U778 & U952; 
assign U638 = ~(U786 & U784 & U951); 
assign U662 = U589 & U937; 
assign U663 = U589 & U785; 
assign U665 = U589 & U940; 
assign U667 = U589 & U778 & U950; 
assign U768 = ~(U1041 & U1040); 
assign U1024 = ~(U957 & U633); 
assign U1026 = ~(U957 & U634); 
assign U1028 = ~(U957 & U635); 
assign U1030 = ~(U957 & U636); 
assign R794_U69 = ~R794_U27; 
assign SUB_60_U6 = ~(SUB_60_U75 & SUB_60_U79); 
assign U592 = SUB_60_U6 & FLAG_REG_SCAN_IN & STATO_REG_0__SCAN_IN & STATO_REG_1__SCAN_IN; 
assign U639 = ~(U611 & U784 & U622); 
assign U640 = ~(U953 & U786 & U623); 
assign U641 = ~(U622 & U954); 
assign U642 = ~(U955 & U784 & U623); 
assign U683 = ~SUB_60_U6; 
assign U862 = SUB_60_U27 | SUB_60_U28 | SUB_60_U6 | SUB_60_U25 | U769; 
assign R794_U14 = ~U638; 
assign R794_U53 = ~(U638 & R794_U15); 
assign R794_U72 = ~(U638 & R794_U15); 
assign U702 = ~(U683 & STATO_REG_1__SCAN_IN); 
assign U804 = ~(ADD_283_U11 & U592); 
assign U806 = ~(ADD_283_U12 & U592); 
assign U808 = ~(ADD_283_U13 & U592); 
assign U810 = ~(ADD_283_U14 & U592); 
assign U812 = ~(ADD_283_U5 & U592); 
assign R794_U7 = ~U642; 
assign R794_U8 = ~U641; 
assign R794_U10 = ~U640; 
assign R794_U12 = ~U639; 
assign R794_U39 = ~(U642 & R794_U19); 
assign R794_U41 = ~(U641 & R794_U9); 
assign R794_U45 = ~(U640 & R794_U11); 
assign R794_U49 = ~(U639 & R794_U13); 
assign R794_U55 = ~(U636 & R794_U14); 
assign R794_U73 = ~(U636 & R794_U14); 
assign R794_U77 = ~(U639 & R794_U13); 
assign R794_U82 = ~(U640 & R794_U11); 
assign R794_U87 = ~(U641 & R794_U9); 
assign U685 = ~(U800 & U702 & STATO_REG_0__SCAN_IN); 
assign U798 = ~U702; 
assign R794_U28 = ~(R794_U73 & R794_U72); 
assign R794_U40 = ~R794_U39; 
assign R794_U42 = ~(R794_U41 & R794_U39); 
assign R794_U43 = ~(U755 & R794_U8); 
assign R794_U47 = ~(U753 & R794_U10); 
assign R794_U51 = ~(U751 & R794_U12); 
assign R794_U62 = ~(U757 & R794_U7); 
assign R794_U78 = ~(U751 & R794_U12); 
assign R794_U83 = ~(U753 & R794_U10); 
assign R794_U88 = ~(U755 & R794_U8); 
assign U801 = ~U685; 
assign U863 = ~(U798 & SUB_73_U6 & U862); 
assign U871 = ~(U798 & U862 & STATO_REG_0__SCAN_IN); 
assign U872 = ~(U685 & FLAG_REG_SCAN_IN); 
assign R794_U6 = ~(R794_U39 & R794_U62); 
assign R794_U29 = ~(R794_U78 & R794_U77); 
assign R794_U30 = ~(R794_U83 & R794_U82); 
assign R794_U31 = ~(R794_U88 & R794_U87); 
assign R794_U38 = ~(R794_U43 & R794_U42); 
assign R794_U74 = ~R794_U28; 
assign U668 = ~(U872 & U871); 
assign U770 = ~(U799 & U863); 
assign U803 = ~(U801 & U802); 
assign U1038 = ~(R794_U6 & U772); 
assign R794_U44 = ~R794_U38; 
assign R794_U46 = ~(R794_U45 & R794_U38); 
assign R794_U79 = ~R794_U29; 
assign R794_U84 = ~R794_U30; 
assign R794_U86 = ~(R794_U30 & R794_U38); 
assign R794_U89 = ~R794_U31; 
assign R794_U91 = ~(R794_U31 & R794_U39); 
assign U767 = ~(U1039 & U1038); 
assign U805 = ~(U803 & NUM_REG_4__SCAN_IN); 
assign U807 = ~(U803 & NUM_REG_3__SCAN_IN); 
assign U809 = ~(U803 & NUM_REG_2__SCAN_IN); 
assign U811 = ~(U803 & NUM_REG_1__SCAN_IN); 
assign U813 = ~(U803 & NUM_REG_0__SCAN_IN); 
assign U864 = ~U770; 
assign U977 = ~(U770 & U624); 
assign U979 = ~(U770 & U632); 
assign U981 = ~(U770 & U631); 
assign U983 = ~(U770 & U859); 
assign U985 = ~(U770 & U629); 
assign U987 = ~(U770 & U861); 
assign U989 = ~(U770 & U627); 
assign U991 = ~(U770 & U626); 
assign U993 = ~(U770 & U625); 
assign R794_U37 = ~(R794_U47 & R794_U46); 
assign R794_U85 = ~(R794_U44 & R794_U84); 
assign R794_U90 = ~(R794_U40 & R794_U89); 
assign U676 = ~(U813 & U812); 
assign U677 = ~(U811 & U810); 
assign U678 = ~(U809 & U808); 
assign U679 = ~(U807 & U806); 
assign U680 = ~(U805 & U804); 
assign U976 = ~(U864 & MAX_REG_8__SCAN_IN); 
assign U978 = ~(U864 & MAX_REG_7__SCAN_IN); 
assign U980 = ~(U864 & MAX_REG_6__SCAN_IN); 
assign U982 = ~(U864 & MAX_REG_5__SCAN_IN); 
assign U984 = ~(U864 & MAX_REG_4__SCAN_IN); 
assign U986 = ~(U864 & MAX_REG_3__SCAN_IN); 
assign U988 = ~(U864 & MAX_REG_2__SCAN_IN); 
assign U990 = ~(U864 & MAX_REG_1__SCAN_IN); 
assign U992 = ~(U864 & MAX_REG_0__SCAN_IN); 
assign R794_U25 = ~(R794_U86 & R794_U85); 
assign R794_U26 = ~(R794_U91 & R794_U90); 
assign R794_U48 = ~R794_U37; 
assign R794_U50 = ~(R794_U49 & R794_U37); 
assign R794_U81 = ~(R794_U29 & R794_U37); 
assign GT_172_U10 = U768 | U767; 
assign GT_178_U7 = U768 & U767; 
assign U736 = ~(U977 & U976); 
assign U737 = ~(U979 & U978); 
assign U738 = ~(U981 & U980); 
assign U739 = ~(U983 & U982); 
assign U740 = ~(U985 & U984); 
assign U741 = ~(U987 & U986); 
assign U742 = ~(U989 & U988); 
assign U743 = ~(U991 & U990); 
assign U744 = ~(U993 & U992); 
assign U1034 = ~(R794_U25 & U772); 
assign U1036 = ~(R794_U26 & U772); 
assign R794_U36 = ~(R794_U51 & R794_U50); 
assign R794_U80 = ~(R794_U48 & R794_U79); 
assign U765 = ~(U1035 & U1034); 
assign U766 = ~(U1037 & U1036); 
assign R794_U24 = ~(R794_U81 & R794_U80); 
assign R794_U52 = ~R794_U36; 
assign R794_U54 = ~(R794_U53 & R794_U36); 
assign R794_U76 = ~(R794_U28 & R794_U36); 
assign U1032 = ~(R794_U24 & U772); 
assign GT_160_U9 = U767 | U768 | U766; 
assign GT_184_U8 = U767 | U768 | U766 | U765; 
assign R794_U35 = ~(R794_U55 & R794_U54); 
assign R794_U75 = ~(R794_U52 & R794_U74); 
assign GT_172_U7 = U766 & GT_172_U10; 
assign GT_169_U7 = U766 & U767; 
assign GT_166_U7 = U767 & U768 & U766; 
assign U764 = ~(U1033 & U1032); 
assign GT_160_U7 = U765 & GT_160_U9; 
assign R794_U23 = ~(R794_U76 & R794_U75); 
assign R794_U56 = ~R794_U35; 
assign R794_U58 = ~(R794_U57 & R794_U35); 
assign R794_U71 = ~(R794_U27 & R794_U35); 
assign U1031 = ~(R794_U23 & U771); 
assign R794_U18 = ~(R794_U59 & R794_U58); 
assign R794_U70 = ~(R794_U56 & R794_U69); 
assign U763 = ~(U1031 & U1030); 
assign R794_U22 = ~(R794_U71 & R794_U70); 
assign R794_U60 = ~R794_U18; 
assign R794_U65 = ~(U634 & R794_U18); 
assign U1029 = ~(R794_U22 & U771); 
assign GT_166_U9 = U764 | U765 | U763; 
assign R794_U33 = ~(R794_U60 & R794_U34); 
assign R794_U66 = ~(R794_U60 & R794_U34); 
assign GT_172_U9 = U764 | U765 | U763; 
assign GT_181_U8 = U765 | U767 | U764 | U766 | U763; 
assign GT_169_U9 = U764 | U765 | U763; 
assign GT_178_U9 = U765 | U766 | U764 | U763; 
assign U762 = ~(U1029 & U1028); 
assign R794_U21 = ~(R794_U66 & R794_U65); 
assign R794_U61 = ~R794_U33; 
assign R794_U63 = ~(U633 & R794_U33); 
assign U1027 = ~(R794_U21 & U771); 
assign R794_U64 = ~(R794_U61 & R794_U32); 
assign GT_175_U8 = U764 | U765 | U766 | U763 | U762; 
assign U761 = ~(U1027 & U1026); 
assign R794_U20 = ~(R794_U64 & R794_U63); 
assign U1025 = ~(R794_U20 & U771); 
assign GT_160_U8 = ~(U761 | U762 | GT_160_U7 | U763 | U764); 
assign GT_163_U7 = ~(U761 | U762 | U763 | U764 | U765); 
assign GT_184_U6 = ~(U761 | U762 | GT_184_U8 | U764 | U763); 
assign GT_175_U7 = ~(U761 | GT_175_U8); 
assign GT_172_U8 = ~(U761 | U762 | GT_172_U7 | GT_172_U9); 
assign GT_181_U7 = ~(U761 | GT_181_U8 | U762); 
assign GT_169_U8 = ~(U761 | U762 | GT_169_U7 | GT_169_U9); 
assign GT_178_U8 = ~(U761 | U762 | GT_178_U7 | GT_178_U9); 
assign GT_166_U8 = ~(U761 | U762 | GT_166_U7 | GT_166_U9); 
assign U760 = ~(U1025 & U1024); 
assign GT_160_U6 = ~(U760 | GT_160_U8); 
assign GT_163_U6 = ~(U760 | GT_163_U7); 
assign GT_184_U7 = ~(GT_184_U6 | U760); 
assign GT_175_U6 = ~(U760 | GT_175_U7); 
assign GT_172_U6 = ~(U760 | GT_172_U8); 
assign GT_181_U6 = ~(U760 | GT_181_U7); 
assign GT_169_U6 = ~(U760 | GT_169_U8); 
assign GT_178_U6 = ~(U760 | GT_178_U8); 
assign GT_166_U6 = ~(U760 | GT_166_U8); 
assign U619 = ~(GT_160_U6 | GT_163_U6 | GT_166_U6); 
assign U715 = ~GT_175_U6; 
assign U717 = GT_169_U6 | GT_172_U6; 
assign U718 = ~GT_181_U6; 
assign U773 = ~GT_160_U6; 
assign U775 = ~GT_163_U6; 
assign U777 = ~GT_178_U6; 
assign U779 = ~GT_166_U6; 
assign U781 = ~GT_172_U6; 
assign U788 = ~GT_169_U6; 
assign U912 = GT_178_U6 | GT_181_U6; 
assign U923 = GT_166_U6 | GT_184_U7 | GT_181_U6 | GT_178_U6; 
assign U925 = GT_181_U6 | GT_184_U7; 
assign U716 = ~(GT_184_U7 & U718); 
assign U909 = ~U717; 
assign U910 = ~(U717 & U779); 
assign U911 = ~(GT_175_U6 & U779); 
assign U913 = ~(U912 & U779); 
assign U920 = ~(U619 & U717); 
assign U926 = ~(U777 & U925); 
assign U617 = U775 & U773 & U910; 
assign U620 = U909 & U619; 
assign U650 = U589 & U920; 
assign U915 = ~U716; 
assign U921 = ~(U715 & U777 & U716); 
assign U927 = ~(U715 & U781 & U926); 
assign U618 = U617 & U911; 
assign U916 = ~(U915 & U777); 
assign U919 = ~(U715 & U777 & GT_181_U6 & U620); 
assign U922 = ~(U620 & U921); 
assign U928 = ~(U788 & U927); 
assign U649 = U589 & U919; 
assign U651 = U589 & U922; 
assign U914 = ~(U913 & U618 & RES_DISP_REG_SCAN_IN); 
assign U917 = ~(U715 & U779 & U916); 
assign U924 = ~(U618 & U923); 
assign U929 = ~(U928 & U779); 
assign U647 = U914 & U705; 
assign U652 = U589 & U924; 
assign U918 = ~(U617 & U917); 
assign U930 = ~(U775 & U929); 
assign U648 = U589 & U918; 
assign U653 = U589 & U773 & U930; 
endmodule 
