module b01_C( LINE1, LINE2, STATO_REG_2__SCAN_IN, STATO_REG_1__SCAN_IN, STATO_REG_0__SCAN_IN, U35, U36, U44, U45); 
input LINE1, LINE2, STATO_REG_2__SCAN_IN, STATO_REG_1__SCAN_IN, STATO_REG_0__SCAN_IN; 
output U35, U36, U44, U45; 
wire U34, U37, U38, U39, U40, U41, U42, U43, U46, U47, U48, U49, U50, U51, U52, U53, U54, U55, U56, U57, U58, U59, U60, U61, U62, U63, U64, U65, U66, U67, U68, U69, U70, U71, U72, U73; 
assign U37 = LINE2 | LINE1; 
assign U38 = ~STATO_REG_2__SCAN_IN; 
assign U39 = ~STATO_REG_1__SCAN_IN; 
assign U40 = ~LINE2; 
assign U41 = ~LINE1; 
assign U42 = ~STATO_REG_0__SCAN_IN; 
assign U47 = ~(LINE1 & LINE2); 
assign U34 = U38 & STATO_REG_1__SCAN_IN & STATO_REG_0__SCAN_IN; 
assign U43 = ~(U42 & STATO_REG_1__SCAN_IN); 
assign U49 = ~U37; 
assign U51 = ~U47; 
assign U54 = ~(U47 & STATO_REG_2__SCAN_IN); 
assign U55 = ~(U39 & U47 & STATO_REG_0__SCAN_IN); 
assign U62 = ~(U37 & U42); 
assign U63 = ~(U47 & STATO_REG_0__SCAN_IN); 
assign U69 = ~(LINE1 & U40); 
assign U70 = ~(LINE2 & U41); 
assign U46 = ~(U70 & U69); 
assign U48 = ~(U43 & STATO_REG_2__SCAN_IN); 
assign U50 = ~(U49 & U42); 
assign U52 = ~U43; 
assign U53 = ~(U47 & U43); 
assign U61 = ~(U49 & STATO_REG_1__SCAN_IN); 
assign U64 = ~(U51 & U42); 
assign U66 = ~(U43 & U37 & STATO_REG_2__SCAN_IN); 
assign U67 = ~(U34 & U47); 
assign U56 = ~(U52 & U54); 
assign U57 = ~(U62 & U61 & STATO_REG_2__SCAN_IN); 
assign U58 = ~U48; 
assign U59 = ~(U53 & U38); 
assign U60 = ~(U50 & U39 & STATO_REG_2__SCAN_IN); 
assign U65 = ~(U64 & U63 & U39 & U38); 
assign U68 = ~(U51 & U52); 
assign U71 = ~U46; 
assign U73 = ~(U46 & U48); 
assign U35 = ~(U68 & U67 & U66 & U65); 
assign U36 = ~(U57 & U55 & U56); 
assign U45 = ~(U60 & U59); 
assign U72 = ~(U58 & U71); 
assign U44 = ~(U73 & U72); 
endmodule 
