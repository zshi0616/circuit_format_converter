module b12_C( GAMMA_REG_0__SCAN_IN, START, K_3_, K_2_, K_1_, K_0_, COUNT_REG_0__SCAN_IN, MEMORY_REG_31__1__SCAN_IN, MEMORY_REG_31__0__SCAN_IN, MEMORY_REG_30__1__SCAN_IN, MEMORY_REG_30__0__SCAN_IN, MEMORY_REG_29__1__SCAN_IN, MEMORY_REG_29__0__SCAN_IN, MEMORY_REG_28__1__SCAN_IN, MEMORY_REG_28__0__SCAN_IN, MEMORY_REG_27__1__SCAN_IN, MEMORY_REG_27__0__SCAN_IN, MEMORY_REG_26__1__SCAN_IN, MEMORY_REG_26__0__SCAN_IN, MEMORY_REG_25__1__SCAN_IN, MEMORY_REG_25__0__SCAN_IN, MEMORY_REG_24__1__SCAN_IN, MEMORY_REG_24__0__SCAN_IN, MEMORY_REG_23__1__SCAN_IN, MEMORY_REG_23__0__SCAN_IN, MEMORY_REG_22__1__SCAN_IN, MEMORY_REG_22__0__SCAN_IN, MEMORY_REG_21__1__SCAN_IN, MEMORY_REG_21__0__SCAN_IN, MEMORY_REG_20__1__SCAN_IN, MEMORY_REG_20__0__SCAN_IN, MEMORY_REG_19__1__SCAN_IN, MEMORY_REG_19__0__SCAN_IN, MEMORY_REG_18__1__SCAN_IN, MEMORY_REG_18__0__SCAN_IN, MEMORY_REG_17__1__SCAN_IN, MEMORY_REG_17__0__SCAN_IN, MEMORY_REG_16__1__SCAN_IN, MEMORY_REG_16__0__SCAN_IN, MEMORY_REG_15__1__SCAN_IN, MEMORY_REG_15__0__SCAN_IN, MEMORY_REG_14__1__SCAN_IN, MEMORY_REG_14__0__SCAN_IN, MEMORY_REG_13__1__SCAN_IN, MEMORY_REG_13__0__SCAN_IN, MEMORY_REG_12__1__SCAN_IN, MEMORY_REG_12__0__SCAN_IN, MEMORY_REG_11__1__SCAN_IN, MEMORY_REG_11__0__SCAN_IN, MEMORY_REG_10__1__SCAN_IN, MEMORY_REG_10__0__SCAN_IN, MEMORY_REG_9__1__SCAN_IN, MEMORY_REG_9__0__SCAN_IN, MEMORY_REG_8__1__SCAN_IN, MEMORY_REG_8__0__SCAN_IN, MEMORY_REG_7__1__SCAN_IN, MEMORY_REG_7__0__SCAN_IN, MEMORY_REG_6__1__SCAN_IN, MEMORY_REG_6__0__SCAN_IN, MEMORY_REG_5__1__SCAN_IN, MEMORY_REG_5__0__SCAN_IN, MEMORY_REG_4__1__SCAN_IN, MEMORY_REG_4__0__SCAN_IN, MEMORY_REG_3__1__SCAN_IN, MEMORY_REG_3__0__SCAN_IN, MEMORY_REG_2__1__SCAN_IN, MEMORY_REG_2__0__SCAN_IN, MEMORY_REG_1__1__SCAN_IN, MEMORY_REG_1__0__SCAN_IN, MEMORY_REG_0__1__SCAN_IN, MEMORY_REG_0__0__SCAN_IN, NL_REG_3__SCAN_IN, NL_REG_2__SCAN_IN, NL_REG_1__SCAN_IN, NL_REG_0__SCAN_IN, SCAN_REG_4__SCAN_IN, SCAN_REG_3__SCAN_IN, SCAN_REG_2__SCAN_IN, SCAN_REG_1__SCAN_IN, SCAN_REG_0__SCAN_IN, MAX_REG_4__SCAN_IN, MAX_REG_3__SCAN_IN, MAX_REG_2__SCAN_IN, MAX_REG_1__SCAN_IN, MAX_REG_0__SCAN_IN, IND_REG_1__SCAN_IN, IND_REG_0__SCAN_IN, TIMEBASE_REG_5__SCAN_IN, TIMEBASE_REG_4__SCAN_IN, TIMEBASE_REG_3__SCAN_IN, TIMEBASE_REG_2__SCAN_IN, TIMEBASE_REG_1__SCAN_IN, TIMEBASE_REG_0__SCAN_IN, COUNT_REG2_5__SCAN_IN, COUNT_REG2_4__SCAN_IN, COUNT_REG2_3__SCAN_IN, COUNT_REG2_2__SCAN_IN, COUNT_REG2_1__SCAN_IN, COUNT_REG2_0__SCAN_IN, SOUND_REG_2__SCAN_IN, SOUND_REG_1__SCAN_IN, SOUND_REG_0__SCAN_IN, ADDRESS_REG_4__SCAN_IN, ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, DATA_IN_REG_1__SCAN_IN, DATA_IN_REG_0__SCAN_IN, S_REG_SCAN_IN, PLAY_REG_SCAN_IN, NLOSS_REG_SCAN_IN, SPEAKER_REG_SCAN_IN, WR_REG_SCAN_IN, COUNTER_REG_2__SCAN_IN, COUNTER_REG_1__SCAN_IN, COUNTER_REG_0__SCAN_IN, COUNT_REG_1__SCAN_IN, NUM_REG_1__SCAN_IN, NUM_REG_0__SCAN_IN, DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN, GAMMA_REG_4__SCAN_IN, GAMMA_REG_3__SCAN_IN, GAMMA_REG_2__SCAN_IN, GAMMA_REG_1__SCAN_IN, U1381, U1382, U1383, U1384, U1385, U1386, U1387, U1388, U1389, U1390, U1392, U1393, U1394, U1395, U1396, U1397, U1398, U1399, U1400, U1401, U1402, U1403, U1404, U1405, U1406, U1407, U1408, U1409, U1410, U1411, U1412, U1413, U1414, U1415, U1416, U1417, U1418, U1419, U1420, U1421, U1422, U1423, U1424, U1425, U1426, U1427, U1428, U1429, U1430, U1431, U1432, U1433, U1434, U1435, U1436, U1437, U1438, U1439, U1440, U1441, U1442, U1443, U1444, U1445, U1446, U1447, U1448, U1449, U1450, U1451, U1452, U1453, U1454, U1455, U1456, U1457, U1458, U1459, U1460, U1461, U1462, U1463, U1464, U1465, U1466, U1467, U1468, U1469, U1470, U1471, U1472, U1473, U1474, U1475, U1476, U1477, U1478, U1479, U1480, U1481, U1482, U1483, U1484, U1485, U1486, U1563, U1564, U1565, U1566, U1567, U1568, U1569, U1570, U1571, U1572, U1573, U1574, U1575); 
input GAMMA_REG_0__SCAN_IN, START, K_3_, K_2_, K_1_, K_0_, COUNT_REG_0__SCAN_IN, MEMORY_REG_31__1__SCAN_IN, MEMORY_REG_31__0__SCAN_IN, MEMORY_REG_30__1__SCAN_IN, MEMORY_REG_30__0__SCAN_IN, MEMORY_REG_29__1__SCAN_IN, MEMORY_REG_29__0__SCAN_IN, MEMORY_REG_28__1__SCAN_IN, MEMORY_REG_28__0__SCAN_IN, MEMORY_REG_27__1__SCAN_IN, MEMORY_REG_27__0__SCAN_IN, MEMORY_REG_26__1__SCAN_IN, MEMORY_REG_26__0__SCAN_IN, MEMORY_REG_25__1__SCAN_IN, MEMORY_REG_25__0__SCAN_IN, MEMORY_REG_24__1__SCAN_IN, MEMORY_REG_24__0__SCAN_IN, MEMORY_REG_23__1__SCAN_IN, MEMORY_REG_23__0__SCAN_IN, MEMORY_REG_22__1__SCAN_IN, MEMORY_REG_22__0__SCAN_IN, MEMORY_REG_21__1__SCAN_IN, MEMORY_REG_21__0__SCAN_IN, MEMORY_REG_20__1__SCAN_IN, MEMORY_REG_20__0__SCAN_IN, MEMORY_REG_19__1__SCAN_IN, MEMORY_REG_19__0__SCAN_IN, MEMORY_REG_18__1__SCAN_IN, MEMORY_REG_18__0__SCAN_IN, MEMORY_REG_17__1__SCAN_IN, MEMORY_REG_17__0__SCAN_IN, MEMORY_REG_16__1__SCAN_IN, MEMORY_REG_16__0__SCAN_IN, MEMORY_REG_15__1__SCAN_IN, MEMORY_REG_15__0__SCAN_IN, MEMORY_REG_14__1__SCAN_IN, MEMORY_REG_14__0__SCAN_IN, MEMORY_REG_13__1__SCAN_IN, MEMORY_REG_13__0__SCAN_IN, MEMORY_REG_12__1__SCAN_IN, MEMORY_REG_12__0__SCAN_IN, MEMORY_REG_11__1__SCAN_IN, MEMORY_REG_11__0__SCAN_IN, MEMORY_REG_10__1__SCAN_IN, MEMORY_REG_10__0__SCAN_IN, MEMORY_REG_9__1__SCAN_IN, MEMORY_REG_9__0__SCAN_IN, MEMORY_REG_8__1__SCAN_IN, MEMORY_REG_8__0__SCAN_IN, MEMORY_REG_7__1__SCAN_IN, MEMORY_REG_7__0__SCAN_IN, MEMORY_REG_6__1__SCAN_IN, MEMORY_REG_6__0__SCAN_IN, MEMORY_REG_5__1__SCAN_IN, MEMORY_REG_5__0__SCAN_IN, MEMORY_REG_4__1__SCAN_IN, MEMORY_REG_4__0__SCAN_IN, MEMORY_REG_3__1__SCAN_IN, MEMORY_REG_3__0__SCAN_IN, MEMORY_REG_2__1__SCAN_IN, MEMORY_REG_2__0__SCAN_IN, MEMORY_REG_1__1__SCAN_IN, MEMORY_REG_1__0__SCAN_IN, MEMORY_REG_0__1__SCAN_IN, MEMORY_REG_0__0__SCAN_IN, NL_REG_3__SCAN_IN, NL_REG_2__SCAN_IN, NL_REG_1__SCAN_IN, NL_REG_0__SCAN_IN, SCAN_REG_4__SCAN_IN, SCAN_REG_3__SCAN_IN, SCAN_REG_2__SCAN_IN, SCAN_REG_1__SCAN_IN, SCAN_REG_0__SCAN_IN, MAX_REG_4__SCAN_IN, MAX_REG_3__SCAN_IN, MAX_REG_2__SCAN_IN, MAX_REG_1__SCAN_IN, MAX_REG_0__SCAN_IN, IND_REG_1__SCAN_IN, IND_REG_0__SCAN_IN, TIMEBASE_REG_5__SCAN_IN, TIMEBASE_REG_4__SCAN_IN, TIMEBASE_REG_3__SCAN_IN, TIMEBASE_REG_2__SCAN_IN, TIMEBASE_REG_1__SCAN_IN, TIMEBASE_REG_0__SCAN_IN, COUNT_REG2_5__SCAN_IN, COUNT_REG2_4__SCAN_IN, COUNT_REG2_3__SCAN_IN, COUNT_REG2_2__SCAN_IN, COUNT_REG2_1__SCAN_IN, COUNT_REG2_0__SCAN_IN, SOUND_REG_2__SCAN_IN, SOUND_REG_1__SCAN_IN, SOUND_REG_0__SCAN_IN, ADDRESS_REG_4__SCAN_IN, ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, DATA_IN_REG_1__SCAN_IN, DATA_IN_REG_0__SCAN_IN, S_REG_SCAN_IN, PLAY_REG_SCAN_IN, NLOSS_REG_SCAN_IN, SPEAKER_REG_SCAN_IN, WR_REG_SCAN_IN, COUNTER_REG_2__SCAN_IN, COUNTER_REG_1__SCAN_IN, COUNTER_REG_0__SCAN_IN, COUNT_REG_1__SCAN_IN, NUM_REG_1__SCAN_IN, NUM_REG_0__SCAN_IN, DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN, GAMMA_REG_4__SCAN_IN, GAMMA_REG_3__SCAN_IN, GAMMA_REG_2__SCAN_IN, GAMMA_REG_1__SCAN_IN; 
output U1381, U1382, U1383, U1384, U1385, U1386, U1387, U1388, U1389, U1390, U1392, U1393, U1394, U1395, U1396, U1397, U1398, U1399, U1400, U1401, U1402, U1403, U1404, U1405, U1406, U1407, U1408, U1409, U1410, U1411, U1412, U1413, U1414, U1415, U1416, U1417, U1418, U1419, U1420, U1421, U1422, U1423, U1424, U1425, U1426, U1427, U1428, U1429, U1430, U1431, U1432, U1433, U1434, U1435, U1436, U1437, U1438, U1439, U1440, U1441, U1442, U1443, U1444, U1445, U1446, U1447, U1448, U1449, U1450, U1451, U1452, U1453, U1454, U1455, U1456, U1457, U1458, U1459, U1460, U1461, U1462, U1463, U1464, U1465, U1466, U1467, U1468, U1469, U1470, U1471, U1472, U1473, U1474, U1475, U1476, U1477, U1478, U1479, U1480, U1481, U1482, U1483, U1484, U1485, U1486, U1563, U1564, U1565, U1566, U1567, U1568, U1569, U1570, U1571, U1572, U1573, U1574, U1575; 
wire U1305, U1306, U1307, U1308, U1309, U1310, U1311, U1312, U1313, U1314, U1315, U1316, U1317, U1318, U1319, U1320, U1321, U1322, U1323, U1324, U1325, U1326, U1327, U1328, U1329, U1330, U1331, U1332, U1333, U1334, U1335, U1336, U1337, U1338, U1339, U1340, U1341, U1342, U1343, U1344, U1345, U1346, U1347, U1348, U1349, U1350, U1351, U1352, U1353, U1354, U1355, U1356, U1357, U1358, U1359, U1360, U1361, U1362, U1363, U1364, U1365, U1366, U1367, U1368, U1369, U1370, U1371, U1372, U1373, U1374, U1375, U1376, U1377, U1378, U1379, U1380, U1391, U1487, U1488, U1489, U1490, U1491, U1492, U1493, U1494, U1495, U1496, U1497, U1498, U1499, U1500, U1501, U1502, U1503, U1504, U1505, U1506, U1507, U1508, U1509, U1510, U1511, U1512, U1513, U1514, U1515, U1516, U1517, U1518, U1519, U1520, U1521, U1522, U1523, U1524, U1525, U1526, U1527, U1528, U1529, U1530, U1531, U1532, U1533, U1534, U1535, U1536, U1537, U1538, U1539, U1540, U1541, U1542, U1543, U1544, U1545, U1546, U1547, U1548, U1549, U1550, U1551, U1552, U1553, U1554, U1555, U1556, U1557, U1558, U1559, U1560, U1561, U1562, U1576, U1577, U1578, U1579, U1580, U1581, U1582, U1583, U1584, U1585, U1586, U1587, U1588, U1589, U1590, U1591, U1592, U1593, U1594, U1595, U1596, U1597, U1598, U1599, U1600, U1601, U1602, U1603, U1604, U1605, U1606, U1607, U1608, U1609, U1610, U1611, U1612, U1613, U1614, U1615, U1616, U1617, U1618, U1619, U1620, U1621, U1622, U1623, U1624, U1625, U1626, U1627, U1628, U1629, U1630, U1631, U1632, U1633, U1634, U1635, U1636, U1637, U1638, U1639, U1640, U1641, U1642, U1643, U1644, U1645, U1646, U1647, U1648, U1649, U1650, U1651, U1652, U1653, U1654, U1655, U1656, U1657, U1658, U1659, U1660, U1661, U1662, U1663, U1664, U1665, U1666, U1667, U1668, U1669, U1670, U1671, U1672, U1673, U1674, U1675, U1676, U1677, U1678, U1679, U1680, U1681, U1682, U1683, U1684, U1685, U1686, U1687, U1688, U1689, U1690, U1691, U1692, U1693, U1694, U1695, U1696, U1697, U1698, U1699, U1700, U1701, U1702, U1703, U1704, U1705, U1706, U1707, U1708, U1709, U1710, U1711, U1712, U1713, U1714, U1715, U1716, U1717, U1718, U1719, U1720, U1721, U1722, U1723, U1724, U1725, U1726, U1727, U1728, U1729, U1730, U1731, U1732, U1733, U1734, U1735, U1736, U1737, U1738, U1739, U1740, U1741, U1742, U1743, U1744, U1745, U1746, U1747, U1748, U1749, U1750, U1751, U1752, U1753, U1754, U1755, U1756, U1757, U1758, U1759, U1760, U1761, U1762, U1763, U1764, U1765, U1766, U1767, U1768, U1769, U1770, U1771, U1772, U1773, U1774, U1775, U1776, U1777, U1778, U1779, U1780, U1781, U1782, U1783, U1784, U1785, U1786, U1787, U1788, U1789, U1790, U1791, U1792, U1793, U1794, U1795, U1796, U1797, U1798, U1799, U1800, U1801, U1802, U1803, U1804, U1805, U1806, U1807, U1808, U1809, U1810, U1811, U1812, U1813, U1814, U1815, U1816, U1817, U1818, U1819, U1820, U1821, U1822, U1823, U1824, U1825, U1826, U1827, U1828, U1829, U1830, U1831, U1832, U1833, U1834, U1835, U1836, U1837, U1838, U1839, U1840, U1841, U1842, U1843, U1844, U1845, U1846, U1847, U1848, U1849, U1850, U1851, U1852, U1853, U1854, U1855, U1856, U1857, U1858, U1859, U1860, U1861, U1862, U1863, U1864, U1865, U1866, U1867, U1868, U1869, U1870, U1871, U1872, U1873, U1874, U1875, U1876, U1877, U1878, U1879, U1880, U1881, U1882, U1883, U1884, U1885, U1886, U1887, U1888, U1889, U1890, U1891, U1892, U1893, U1894, U1895, U1896, U1897, U1898, U1899, U1900, U1901, U1902, U1903, U1904, U1905, U1906, U1907, U1908, U1909, U1910, U1911, U1912, U1913, U1914, U1915, U1916, U1917, U1918, U1919, U1920, U1921, U1922, U1923, U1924, U1925, U1926, U1927, U1928, U1929, U1930, U1931, U1932, U1933, U1934, U1935, U1936, U1937, U1938, U1939, U1940, U1941, U1942, U1943, U1944, U1945, U1946, U1947, U1948, U1949, U1950, U1951, U1952, U1953, U1954, U1955, U1956, U1957, U1958, U1959, U1960, U1961, U1962, U1963, U1964, U1965, U1966, U1967, U1968, U1969, U1970, U1971, U1972, U1973, U1974, U1975, U1976, U1977, U1978, U1979, U1980, U1981, U1982, U1983, U1984, U1985, U1986, U1987, U1988, U1989, U1990, U1991, U1992, U1993, U1994, U1995, U1996, U1997, U1998, U1999, U2000, U2001, U2002, U2003, U2004, U2005, U2006, U2007, U2008, U2009, U2010, U2011, U2012, U2013, U2014, U2015, U2016, U2017, U2018, U2019, U2020, U2021, U2022, U2023, U2024, U2025, U2026, U2027, U2028, U2029, U2030, U2031, U2032, U2033, U2034, U2035, U2036, U2037, U2038, U2039, U2040, U2041, U2042, U2043, U2044, U2045, U2046, U2047, U2048, U2049, U2050, U2051, U2052, U2053, U2054, U2055, U2056, U2057, U2058, U2059, U2060, U2061, U2062, U2063, U2064, U2065, U2066, U2067, U2068, U2069, U2070, U2071, U2072, U2073, U2074, U2075, U2076, U2077, U2078, U2079, U2080, U2081, U2082, U2083, U2084, U2085, U2086, U2087, U2088, U2089, U2090, U2091, U2092, U2093, U2094, U2095, U2096, U2097, U2098, U2099, U2100, U2101, U2102, U2103, U2104, U2105, U2106, U2107, U2108, U2109, U2110, U2111, U2112, U2113, U2114, U2115, U2116, U2117, U2118, U2119, U2120, U2121, U2122, U2123, U2124, U2125, U2126, U2127, U2128, U2129, U2130, U2131, U2132, U2133, U2134, U2135, U2136, U2137, U2138, U2139, U2140, U2141, U2142, U2143, U2144, U2145, U2146, U2147, U2148, U2149, U2150, U2151, U2152, U2153, U2154, U2155, U2156, U2157, U2158, U2159, U2160, U2161, U2162, U2163, U2164, U2165, U2166, U2167, U2168, U2169, U2170, U2171, U2172, U2173, U2174, U2175, U2176, U2177, R745_U6, R745_U7, R745_U8, R745_U9, R745_U10, R745_U11, R745_U12, R745_U13, R745_U14, R745_U15, R745_U16, R745_U17, R745_U18, R745_U19, R745_U20, R745_U21, R745_U22, R745_U23, R745_U24, R745_U25, R745_U26, R745_U27, R745_U28, R745_U29, R745_U30, R730_U5, R730_U6, R730_U7, R730_U8, R730_U9, R730_U10, R730_U11, R730_U12, R730_U13, R730_U14, R730_U15, R730_U16, R730_U17, R730_U18, R730_U19, R730_U20, R730_U21, R730_U22, R730_U23, R730_U24, R730_U25, R730_U26, R730_U27, R785_U5, R785_U6, R785_U7, R785_U8, R785_U9, R785_U10, R785_U11, R785_U12, R785_U13, R785_U14, R785_U15, R785_U16, R785_U17, R785_U18, R785_U19, R785_U20, R785_U21, R785_U22, R785_U23, R785_U24, R785_U25, R785_U26, R785_U27; 
assign U1307 = DATA_IN_REG_0__SCAN_IN & WR_REG_SCAN_IN; 
assign U1308 = DATA_IN_REG_1__SCAN_IN & WR_REG_SCAN_IN; 
assign U1318 = ~(K_0_ | K_1_); 
assign U1324 = ADDRESS_REG_4__SCAN_IN & ADDRESS_REG_3__SCAN_IN & ADDRESS_REG_1__SCAN_IN; 
assign U1325 = ADDRESS_REG_2__SCAN_IN & ADDRESS_REG_0__SCAN_IN; 
assign U1334 = ~(ADDRESS_REG_2__SCAN_IN | ADDRESS_REG_0__SCAN_IN); 
assign U1361 = ~(ADDRESS_REG_4__SCAN_IN | ADDRESS_REG_3__SCAN_IN | ADDRESS_REG_1__SCAN_IN); 
assign U1391 = ~COUNT_REG_0__SCAN_IN; 
assign U1487 = ~ADDRESS_REG_4__SCAN_IN; 
assign U1488 = ~ADDRESS_REG_3__SCAN_IN; 
assign U1489 = ~ADDRESS_REG_1__SCAN_IN; 
assign U1490 = ~ADDRESS_REG_2__SCAN_IN; 
assign U1491 = ~ADDRESS_REG_0__SCAN_IN; 
assign U1494 = START | GAMMA_REG_0__SCAN_IN; 
assign U1505 = ~SCAN_REG_0__SCAN_IN; 
assign U1506 = ~MAX_REG_0__SCAN_IN; 
assign U1507 = ~SCAN_REG_1__SCAN_IN; 
assign U1508 = ~MAX_REG_1__SCAN_IN; 
assign U1509 = ~SCAN_REG_2__SCAN_IN; 
assign U1510 = ~MAX_REG_2__SCAN_IN; 
assign U1511 = ~SCAN_REG_3__SCAN_IN; 
assign U1512 = ~MAX_REG_3__SCAN_IN; 
assign U1513 = ~SCAN_REG_4__SCAN_IN; 
assign U1514 = ~MAX_REG_4__SCAN_IN; 
assign U1517 = ~IND_REG_0__SCAN_IN; 
assign U1518 = ~IND_REG_1__SCAN_IN; 
assign U1519 = ~DATA_OUT_REG_1__SCAN_IN; 
assign U1520 = ~DATA_OUT_REG_0__SCAN_IN; 
assign U1521 = ~(DATA_OUT_REG_1__SCAN_IN & DATA_OUT_REG_0__SCAN_IN); 
assign U1535 = ~K_2_; 
assign U1536 = ~(MAX_REG_4__SCAN_IN & MAX_REG_3__SCAN_IN & MAX_REG_2__SCAN_IN & MAX_REG_1__SCAN_IN & MAX_REG_0__SCAN_IN); 
assign U1544 = ~COUNT_REG2_4__SCAN_IN; 
assign U1546 = ~COUNT_REG2_2__SCAN_IN; 
assign U1547 = ~COUNT_REG2_1__SCAN_IN; 
assign U1550 = ~SOUND_REG_1__SCAN_IN; 
assign U1552 = ~COUNTER_REG_2__SCAN_IN; 
assign U1553 = ~COUNTER_REG_0__SCAN_IN; 
assign U1554 = ~COUNTER_REG_1__SCAN_IN; 
assign U1556 = ~S_REG_SCAN_IN; 
assign U1557 = ~K_3_; 
assign U1558 = ~K_1_; 
assign U1559 = ~K_0_; 
assign U1578 = ~(COUNT_REG2_5__SCAN_IN | COUNT_REG2_4__SCAN_IN | COUNT_REG2_3__SCAN_IN); 
assign U1601 = ~COUNT_REG2_5__SCAN_IN; 
assign U1602 = ~COUNT_REG2_3__SCAN_IN; 
assign U1603 = ~COUNT_REG2_0__SCAN_IN; 
assign U1605 = ~SOUND_REG_0__SCAN_IN; 
assign U1609 = ~COUNT_REG_1__SCAN_IN; 
assign U1625 = ~START; 
assign U1993 = ~(SOUND_REG_2__SCAN_IN & SOUND_REG_1__SCAN_IN); 
assign U2007 = DATA_OUT_REG_1__SCAN_IN | DATA_OUT_REG_0__SCAN_IN; 
assign U2099 = ~(COUNTER_REG_1__SCAN_IN & COUNTER_REG_0__SCAN_IN); 
assign U2153 = ~(SOUND_REG_2__SCAN_IN & SOUND_REG_0__SCAN_IN); 
assign U2164 = K_0_ | DATA_OUT_REG_0__SCAN_IN; 
assign U2167 = K_2_ | DATA_OUT_REG_0__SCAN_IN; 
assign R730_U5 = ~MAX_REG_0__SCAN_IN; 
assign R730_U6 = ~MAX_REG_1__SCAN_IN; 
assign R730_U7 = ~(MAX_REG_1__SCAN_IN & MAX_REG_0__SCAN_IN); 
assign R730_U8 = ~MAX_REG_2__SCAN_IN; 
assign R730_U10 = ~MAX_REG_3__SCAN_IN; 
assign R730_U15 = ~MAX_REG_4__SCAN_IN; 
assign R785_U5 = ~SCAN_REG_0__SCAN_IN; 
assign R785_U6 = ~SCAN_REG_1__SCAN_IN; 
assign R785_U7 = ~(SCAN_REG_1__SCAN_IN & SCAN_REG_0__SCAN_IN); 
assign R785_U8 = ~SCAN_REG_2__SCAN_IN; 
assign R785_U10 = ~SCAN_REG_3__SCAN_IN; 
assign R785_U15 = ~SCAN_REG_4__SCAN_IN; 
assign U1326 = U1324 & U1325; 
assign U1327 = U1491 & ADDRESS_REG_2__SCAN_IN; 
assign U1329 = U1489 & ADDRESS_REG_4__SCAN_IN & ADDRESS_REG_3__SCAN_IN; 
assign U1332 = U1490 & ADDRESS_REG_0__SCAN_IN; 
assign U1335 = U1334 & U1324; 
assign U1338 = U1488 & ADDRESS_REG_4__SCAN_IN & ADDRESS_REG_1__SCAN_IN; 
assign U1341 = U1488 & U1489 & ADDRESS_REG_4__SCAN_IN; 
assign U1348 = U1487 & ADDRESS_REG_3__SCAN_IN & ADDRESS_REG_1__SCAN_IN; 
assign U1351 = U1487 & U1489 & ADDRESS_REG_3__SCAN_IN; 
assign U1358 = U1487 & U1488 & ADDRESS_REG_1__SCAN_IN; 
assign U1362 = U1361 & U1325; 
assign U1367 = U1361 & U1334; 
assign U1492 = ~(U1625 & GAMMA_REG_4__SCAN_IN); 
assign U1493 = ~(U1625 & GAMMA_REG_3__SCAN_IN); 
assign U1496 = ~(U1625 & GAMMA_REG_1__SCAN_IN); 
assign U1500 = ~(U1625 & GAMMA_REG_2__SCAN_IN); 
assign U1501 = ~(U1547 & U1546 & U1603 & U1578); 
assign U1523 = ~(U1519 & DATA_OUT_REG_0__SCAN_IN); 
assign U1539 = ~(U1557 & U1535 & U1318); 
assign U1819 = ~U1494; 
assign U1837 = ~U1521; 
assign U1864 = ~U1536; 
assign U1884 = ~(K_2_ & U1558); 
assign U1983 = ~(U1605 & SOUND_REG_2__SCAN_IN); 
assign U1987 = ~(U1605 & SOUND_REG_1__SCAN_IN & COUNTER_REG_0__SCAN_IN); 
assign U2106 = ~(K_3_ & U1521); 
assign U2107 = ~(K_3_ & U1535); 
assign U2108 = ~(K_1_ & U1559); 
assign U2113 = ~(U2099 & U1552); 
assign U2114 = ~(U1510 & SCAN_REG_2__SCAN_IN); 
assign U2115 = ~(U1509 & MAX_REG_2__SCAN_IN); 
assign U2116 = ~(U1506 & SCAN_REG_0__SCAN_IN); 
assign U2117 = ~(U1505 & MAX_REG_0__SCAN_IN); 
assign U2118 = ~(U1508 & SCAN_REG_1__SCAN_IN); 
assign U2119 = ~(U1507 & MAX_REG_1__SCAN_IN); 
assign U2120 = ~(U1512 & SCAN_REG_3__SCAN_IN); 
assign U2121 = ~(U1511 & MAX_REG_3__SCAN_IN); 
assign U2122 = ~(U1514 & SCAN_REG_4__SCAN_IN); 
assign U2123 = ~(U1513 & MAX_REG_4__SCAN_IN); 
assign U2152 = ~(U1605 & COUNTER_REG_0__SCAN_IN); 
assign U2159 = ~(U1520 & K_2_ & DATA_OUT_REG_1__SCAN_IN); 
assign U2160 = ~(K_0_ & U2007); 
assign U2173 = ~(U1553 & COUNTER_REG_1__SCAN_IN); 
assign U2174 = ~(U1554 & COUNTER_REG_0__SCAN_IN); 
assign U2176 = ~(U1391 & COUNT_REG_1__SCAN_IN); 
assign U2177 = ~(U1609 & COUNT_REG_0__SCAN_IN); 
assign R730_U17 = ~R730_U7; 
assign R730_U24 = ~(R730_U7 & MAX_REG_2__SCAN_IN); 
assign R730_U26 = ~(R730_U5 & MAX_REG_1__SCAN_IN); 
assign R730_U27 = ~(R730_U6 & MAX_REG_0__SCAN_IN); 
assign R785_U17 = ~R785_U7; 
assign R785_U24 = ~(R785_U7 & SCAN_REG_2__SCAN_IN); 
assign R785_U26 = ~(R785_U5 & SCAN_REG_1__SCAN_IN); 
assign R785_U27 = ~(R785_U6 & SCAN_REG_0__SCAN_IN); 
assign U1312 = U1492 & U1493; 
assign U1328 = U1327 & U1324; 
assign U1330 = U1329 & U1325; 
assign U1331 = U1329 & U1327; 
assign U1333 = U1332 & U1324; 
assign U1336 = U1332 & U1329; 
assign U1337 = U1334 & U1329; 
assign U1339 = U1338 & U1325; 
assign U1340 = U1338 & U1327; 
assign U1342 = U1341 & U1325; 
assign U1343 = U1341 & U1327; 
assign U1344 = U1338 & U1332; 
assign U1345 = U1338 & U1334; 
assign U1346 = U1341 & U1332; 
assign U1347 = U1341 & U1334; 
assign U1349 = U1348 & U1325; 
assign U1350 = U1348 & U1327; 
assign U1352 = U1351 & U1325; 
assign U1353 = U1351 & U1327; 
assign U1354 = U1348 & U1332; 
assign U1355 = U1348 & U1334; 
assign U1356 = U1351 & U1332; 
assign U1357 = U1351 & U1334; 
assign U1359 = U1358 & U1325; 
assign U1360 = U1358 & U1327; 
assign U1363 = U1361 & U1327; 
assign U1364 = U1358 & U1332; 
assign U1365 = U1358 & U1334; 
assign U1366 = U1361 & U1332; 
assign U1499 = ~(U1500 & U1493); 
assign U1502 = ~(U1494 & U1496); 
assign U1504 = ~(U1500 & U1492); 
assign U1531 = ~(U1819 & U1496); 
assign U1563 = ~(U2177 & U2176); 
assign U1576 = U2119 & U2118 & U2117 & U2116; 
assign U1577 = U2123 & U2122 & U2121 & U2120; 
assign U1611 = ~U1493; 
assign U1614 = ~U1492; 
assign U1616 = ~U1500; 
assign U1618 = ~U1496; 
assign U1622 = ~U1501; 
assign U1659 = ~(U1326 & WR_REG_SCAN_IN); 
assign U1661 = ~(U1308 & U1326); 
assign U1663 = ~(U1307 & U1326); 
assign U1684 = ~(U1335 & WR_REG_SCAN_IN); 
assign U1686 = ~(U1335 & U1308); 
assign U1688 = ~(U1335 & U1307); 
assign U1789 = ~(U1362 & WR_REG_SCAN_IN); 
assign U1791 = ~(U1362 & U1308); 
assign U1793 = ~(U1362 & U1307); 
assign U1814 = ~(U1367 & WR_REG_SCAN_IN); 
assign U1816 = ~(U1367 & U1308); 
assign U1818 = ~(U1367 & U1307); 
assign U1844 = ~U1523; 
assign U1882 = ~U1539; 
assign U1898 = ~(U1819 & U1500 & U1501); 
assign U1913 = ~(U1819 & U1493); 
assign U1960 = ~(U1493 & DATA_OUT_REG_0__SCAN_IN); 
assign U1984 = ~(U1983 & U1550); 
assign U1986 = ~(U2153 & U2152 & U1550); 
assign U1990 = ~(U1550 & U1983 & COUNTER_REG_2__SCAN_IN); 
assign U2035 = ~(U1367 & MEMORY_REG_0__1__SCAN_IN); 
assign U2040 = ~(U1362 & MEMORY_REG_5__1__SCAN_IN); 
assign U2061 = ~(U1335 & MEMORY_REG_26__1__SCAN_IN); 
assign U2066 = ~(U1326 & MEMORY_REG_31__1__SCAN_IN); 
assign U2067 = ~(U1367 & MEMORY_REG_0__0__SCAN_IN); 
assign U2072 = ~(U1362 & MEMORY_REG_5__0__SCAN_IN); 
assign U2093 = ~(U1335 & MEMORY_REG_26__0__SCAN_IN); 
assign U2098 = ~(U1326 & MEMORY_REG_31__0__SCAN_IN); 
assign U2158 = ~(U2106 & U1535); 
assign U2161 = ~(K_1_ & U1523 & U1559); 
assign U2165 = ~(U2108 & DATA_OUT_REG_0__SCAN_IN); 
assign U2168 = ~(U2107 & DATA_OUT_REG_0__SCAN_IN); 
assign U2175 = ~(U2174 & U2173); 
assign R730_U9 = ~(R730_U17 & MAX_REG_2__SCAN_IN); 
assign R730_U14 = ~(R730_U27 & R730_U26); 
assign R730_U25 = ~(R730_U17 & R730_U8); 
assign R785_U9 = ~(R785_U17 & SCAN_REG_2__SCAN_IN); 
assign R785_U14 = ~(R785_U27 & R785_U26); 
assign R785_U25 = ~(R785_U17 & R785_U8); 
assign U1306 = U1312 & U1494; 
assign U1320 = U1614 & U1500; 
assign U1321 = U1616 & U1496; 
assign U1495 = ~(U1611 & U1614); 
assign U1497 = ~(U1618 & U1494); 
assign U1515 = ~(U2115 & U2114 & U1576 & U1577); 
assign U1516 = ~(U1616 & U1611); 
assign U1525 = ~(U1312 & U1819); 
assign U1530 = ~(U1618 & U1819); 
assign U1545 = ~(U1616 & U1614); 
assign U1612 = ~U1502; 
assign U1615 = ~U1499; 
assign U1621 = ~U1504; 
assign U1635 = ~U1531; 
assign U1660 = ~(U1659 & MEMORY_REG_31__1__SCAN_IN); 
assign U1662 = ~(U1659 & MEMORY_REG_31__0__SCAN_IN); 
assign U1664 = ~(U1328 & WR_REG_SCAN_IN); 
assign U1666 = ~(U1328 & U1308); 
assign U1668 = ~(U1328 & U1307); 
assign U1669 = ~(U1330 & WR_REG_SCAN_IN); 
assign U1671 = ~(U1330 & U1308); 
assign U1673 = ~(U1330 & U1307); 
assign U1674 = ~(U1331 & WR_REG_SCAN_IN); 
assign U1676 = ~(U1331 & U1308); 
assign U1678 = ~(U1331 & U1307); 
assign U1679 = ~(U1333 & WR_REG_SCAN_IN); 
assign U1681 = ~(U1333 & U1308); 
assign U1683 = ~(U1333 & U1307); 
assign U1685 = ~(U1684 & MEMORY_REG_26__1__SCAN_IN); 
assign U1687 = ~(U1684 & MEMORY_REG_26__0__SCAN_IN); 
assign U1689 = ~(U1336 & WR_REG_SCAN_IN); 
assign U1691 = ~(U1336 & U1308); 
assign U1693 = ~(U1336 & U1307); 
assign U1694 = ~(U1337 & WR_REG_SCAN_IN); 
assign U1696 = ~(U1337 & U1308); 
assign U1698 = ~(U1337 & U1307); 
assign U1699 = ~(U1339 & WR_REG_SCAN_IN); 
assign U1701 = ~(U1339 & U1308); 
assign U1703 = ~(U1339 & U1307); 
assign U1704 = ~(U1340 & WR_REG_SCAN_IN); 
assign U1706 = ~(U1340 & U1308); 
assign U1708 = ~(U1340 & U1307); 
assign U1709 = ~(U1342 & WR_REG_SCAN_IN); 
assign U1711 = ~(U1342 & U1308); 
assign U1713 = ~(U1342 & U1307); 
assign U1714 = ~(U1343 & WR_REG_SCAN_IN); 
assign U1716 = ~(U1343 & U1308); 
assign U1718 = ~(U1343 & U1307); 
assign U1719 = ~(U1344 & WR_REG_SCAN_IN); 
assign U1721 = ~(U1344 & U1308); 
assign U1723 = ~(U1344 & U1307); 
assign U1724 = ~(U1345 & WR_REG_SCAN_IN); 
assign U1726 = ~(U1345 & U1308); 
assign U1728 = ~(U1345 & U1307); 
assign U1729 = ~(U1346 & WR_REG_SCAN_IN); 
assign U1731 = ~(U1346 & U1308); 
assign U1733 = ~(U1346 & U1307); 
assign U1734 = ~(U1347 & WR_REG_SCAN_IN); 
assign U1736 = ~(U1347 & U1308); 
assign U1738 = ~(U1347 & U1307); 
assign U1739 = ~(U1349 & WR_REG_SCAN_IN); 
assign U1741 = ~(U1349 & U1308); 
assign U1743 = ~(U1349 & U1307); 
assign U1744 = ~(U1350 & WR_REG_SCAN_IN); 
assign U1746 = ~(U1350 & U1308); 
assign U1748 = ~(U1350 & U1307); 
assign U1749 = ~(U1352 & WR_REG_SCAN_IN); 
assign U1751 = ~(U1352 & U1308); 
assign U1753 = ~(U1352 & U1307); 
assign U1754 = ~(U1353 & WR_REG_SCAN_IN); 
assign U1756 = ~(U1353 & U1308); 
assign U1758 = ~(U1353 & U1307); 
assign U1759 = ~(U1354 & WR_REG_SCAN_IN); 
assign U1761 = ~(U1354 & U1308); 
assign U1763 = ~(U1354 & U1307); 
assign U1764 = ~(U1355 & WR_REG_SCAN_IN); 
assign U1766 = ~(U1355 & U1308); 
assign U1768 = ~(U1355 & U1307); 
assign U1769 = ~(U1356 & WR_REG_SCAN_IN); 
assign U1771 = ~(U1356 & U1308); 
assign U1773 = ~(U1356 & U1307); 
assign U1774 = ~(U1357 & WR_REG_SCAN_IN); 
assign U1776 = ~(U1357 & U1308); 
assign U1778 = ~(U1357 & U1307); 
assign U1779 = ~(U1359 & WR_REG_SCAN_IN); 
assign U1781 = ~(U1359 & U1308); 
assign U1783 = ~(U1359 & U1307); 
assign U1784 = ~(U1360 & WR_REG_SCAN_IN); 
assign U1786 = ~(U1360 & U1308); 
assign U1788 = ~(U1360 & U1307); 
assign U1790 = ~(U1789 & MEMORY_REG_5__1__SCAN_IN); 
assign U1792 = ~(U1789 & MEMORY_REG_5__0__SCAN_IN); 
assign U1794 = ~(U1363 & WR_REG_SCAN_IN); 
assign U1796 = ~(U1363 & U1308); 
assign U1798 = ~(U1363 & U1307); 
assign U1799 = ~(U1364 & WR_REG_SCAN_IN); 
assign U1801 = ~(U1364 & U1308); 
assign U1803 = ~(U1364 & U1307); 
assign U1804 = ~(U1365 & WR_REG_SCAN_IN); 
assign U1806 = ~(U1365 & U1308); 
assign U1808 = ~(U1365 & U1307); 
assign U1809 = ~(U1366 & WR_REG_SCAN_IN); 
assign U1811 = ~(U1366 & U1308); 
assign U1813 = ~(U1366 & U1307); 
assign U1815 = ~(U1814 & MEMORY_REG_0__1__SCAN_IN); 
assign U1817 = ~(U1814 & MEMORY_REG_0__0__SCAN_IN); 
assign U1820 = ~(U1616 & U1502); 
assign U1824 = ~(U1611 & U1502); 
assign U1908 = ~(U1312 & U1496); 
assign U1916 = ~(U1616 & U1618); 
assign U1925 = ~(U1616 & U1502 & U1501); 
assign U1935 = ~(U1616 & TIMEBASE_REG_3__SCAN_IN); 
assign U1955 = ~(U1614 & U1499); 
assign U1963 = ~(U1618 & U1492); 
assign U1985 = ~(U1552 & U1984); 
assign U1988 = ~(U1986 & COUNTER_REG_1__SCAN_IN); 
assign U2008 = ~(U2159 & U2158 & U1318); 
assign U2016 = ~(U1502 & U1531); 
assign U2036 = ~(U1366 & MEMORY_REG_1__1__SCAN_IN); 
assign U2037 = ~(U1365 & MEMORY_REG_2__1__SCAN_IN); 
assign U2038 = ~(U1364 & MEMORY_REG_3__1__SCAN_IN); 
assign U2039 = ~(U1363 & MEMORY_REG_4__1__SCAN_IN); 
assign U2041 = ~(U1360 & MEMORY_REG_6__1__SCAN_IN); 
assign U2042 = ~(U1359 & MEMORY_REG_7__1__SCAN_IN); 
assign U2043 = ~(U1357 & MEMORY_REG_8__1__SCAN_IN); 
assign U2044 = ~(U1356 & MEMORY_REG_9__1__SCAN_IN); 
assign U2045 = ~(U1355 & MEMORY_REG_10__1__SCAN_IN); 
assign U2046 = ~(U1354 & MEMORY_REG_11__1__SCAN_IN); 
assign U2047 = ~(U1353 & MEMORY_REG_12__1__SCAN_IN); 
assign U2048 = ~(U1352 & MEMORY_REG_13__1__SCAN_IN); 
assign U2049 = ~(U1350 & MEMORY_REG_14__1__SCAN_IN); 
assign U2050 = ~(U1349 & MEMORY_REG_15__1__SCAN_IN); 
assign U2051 = ~(U1347 & MEMORY_REG_16__1__SCAN_IN); 
assign U2052 = ~(U1346 & MEMORY_REG_17__1__SCAN_IN); 
assign U2053 = ~(U1345 & MEMORY_REG_18__1__SCAN_IN); 
assign U2054 = ~(U1344 & MEMORY_REG_19__1__SCAN_IN); 
assign U2055 = ~(U1343 & MEMORY_REG_20__1__SCAN_IN); 
assign U2056 = ~(U1342 & MEMORY_REG_21__1__SCAN_IN); 
assign U2057 = ~(U1340 & MEMORY_REG_22__1__SCAN_IN); 
assign U2058 = ~(U1339 & MEMORY_REG_23__1__SCAN_IN); 
assign U2059 = ~(U1337 & MEMORY_REG_24__1__SCAN_IN); 
assign U2060 = ~(U1336 & MEMORY_REG_25__1__SCAN_IN); 
assign U2062 = ~(U1333 & MEMORY_REG_27__1__SCAN_IN); 
assign U2063 = ~(U1331 & MEMORY_REG_28__1__SCAN_IN); 
assign U2064 = ~(U1330 & MEMORY_REG_29__1__SCAN_IN); 
assign U2065 = ~(U1328 & MEMORY_REG_30__1__SCAN_IN); 
assign U2068 = ~(U1366 & MEMORY_REG_1__0__SCAN_IN); 
assign U2069 = ~(U1365 & MEMORY_REG_2__0__SCAN_IN); 
assign U2070 = ~(U1364 & MEMORY_REG_3__0__SCAN_IN); 
assign U2071 = ~(U1363 & MEMORY_REG_4__0__SCAN_IN); 
assign U2073 = ~(U1360 & MEMORY_REG_6__0__SCAN_IN); 
assign U2074 = ~(U1359 & MEMORY_REG_7__0__SCAN_IN); 
assign U2075 = ~(U1357 & MEMORY_REG_8__0__SCAN_IN); 
assign U2076 = ~(U1356 & MEMORY_REG_9__0__SCAN_IN); 
assign U2077 = ~(U1355 & MEMORY_REG_10__0__SCAN_IN); 
assign U2078 = ~(U1354 & MEMORY_REG_11__0__SCAN_IN); 
assign U2079 = ~(U1353 & MEMORY_REG_12__0__SCAN_IN); 
assign U2080 = ~(U1352 & MEMORY_REG_13__0__SCAN_IN); 
assign U2081 = ~(U1350 & MEMORY_REG_14__0__SCAN_IN); 
assign U2082 = ~(U1349 & MEMORY_REG_15__0__SCAN_IN); 
assign U2083 = ~(U1347 & MEMORY_REG_16__0__SCAN_IN); 
assign U2084 = ~(U1346 & MEMORY_REG_17__0__SCAN_IN); 
assign U2085 = ~(U1345 & MEMORY_REG_18__0__SCAN_IN); 
assign U2086 = ~(U1344 & MEMORY_REG_19__0__SCAN_IN); 
assign U2087 = ~(U1343 & MEMORY_REG_20__0__SCAN_IN); 
assign U2088 = ~(U1342 & MEMORY_REG_21__0__SCAN_IN); 
assign U2089 = ~(U1340 & MEMORY_REG_22__0__SCAN_IN); 
assign U2090 = ~(U1339 & MEMORY_REG_23__0__SCAN_IN); 
assign U2091 = ~(U1337 & MEMORY_REG_24__0__SCAN_IN); 
assign U2092 = ~(U1336 & MEMORY_REG_25__0__SCAN_IN); 
assign U2094 = ~(U1333 & MEMORY_REG_27__0__SCAN_IN); 
assign U2095 = ~(U1331 & MEMORY_REG_28__0__SCAN_IN); 
assign U2096 = ~(U1330 & MEMORY_REG_29__0__SCAN_IN); 
assign U2097 = ~(U1328 & MEMORY_REG_30__0__SCAN_IN); 
assign U2100 = ~(U1622 & TIMEBASE_REG_5__SCAN_IN); 
assign U2101 = ~(U1622 & TIMEBASE_REG_4__SCAN_IN); 
assign U2102 = ~(U1622 & TIMEBASE_REG_3__SCAN_IN); 
assign U2103 = ~(U1622 & TIMEBASE_REG_2__SCAN_IN); 
assign U2104 = ~(U1622 & TIMEBASE_REG_1__SCAN_IN); 
assign U2105 = ~(U1622 & TIMEBASE_REG_0__SCAN_IN); 
assign U2109 = ~(U2168 & U2167 & U1318); 
assign U2133 = ~(U1502 & U1493 & U1614); 
assign U2154 = ~(U1616 & U1614); 
assign U2166 = ~(U2165 & U2164); 
assign R730_U13 = ~(R730_U25 & R730_U24); 
assign R730_U18 = ~R730_U9; 
assign R730_U22 = ~(R730_U9 & MAX_REG_3__SCAN_IN); 
assign R785_U13 = ~(R785_U25 & R785_U24); 
assign R785_U18 = ~R785_U9; 
assign R785_U22 = ~(R785_U9 & SCAN_REG_3__SCAN_IN); 
assign U1375 = ~(U2100 & U1601); 
assign U1376 = ~(U2101 & U1544); 
assign U1377 = ~(U2102 & U1602); 
assign U1378 = ~(U2103 & U1546); 
assign U1379 = ~(U2104 & U1547); 
assign U1380 = ~(U2105 & U1603); 
assign U1423 = ~(U1818 & U1817); 
assign U1424 = ~(U1816 & U1815); 
assign U1433 = ~(U1793 & U1792); 
assign U1434 = ~(U1791 & U1790); 
assign U1475 = ~(U1688 & U1687); 
assign U1476 = ~(U1686 & U1685); 
assign U1485 = ~(U1663 & U1662); 
assign U1486 = ~(U1661 & U1660); 
assign U1503 = ~(U1612 & U1493); 
assign U1526 = ~(U1616 & U1618 & U1306); 
assign U1528 = ~(U1612 & U1614); 
assign U1584 = U2038 & U2037 & U2036 & U2035; 
assign U1586 = U2046 & U2045 & U2044 & U2043; 
assign U1588 = U2054 & U2053 & U2052 & U2051; 
assign U1590 = U2062 & U2061 & U2060 & U2059; 
assign U1592 = U2070 & U2069 & U2068 & U2067; 
assign U1594 = U2078 & U2077 & U2076 & U2075; 
assign U1596 = U2086 & U2085 & U2084 & U2083; 
assign U1598 = U2094 & U2093 & U2092 & U2091; 
assign U1613 = ~U1525; 
assign U1619 = ~U1530; 
assign U1636 = ~(U2016 & U1500); 
assign U1646 = ~(U1621 & U1611 & U1635); 
assign U1649 = ~(U1635 & U1616 & U1622); 
assign U1650 = ~(U1312 & U1321); 
assign U1651 = ~U1495; 
assign U1653 = ~(U1615 & U1618); 
assign U1654 = ~U1516; 
assign U1655 = ~U1497; 
assign U1656 = ~U1545; 
assign U1665 = ~(U1664 & MEMORY_REG_30__1__SCAN_IN); 
assign U1667 = ~(U1664 & MEMORY_REG_30__0__SCAN_IN); 
assign U1670 = ~(U1669 & MEMORY_REG_29__1__SCAN_IN); 
assign U1672 = ~(U1669 & MEMORY_REG_29__0__SCAN_IN); 
assign U1675 = ~(U1674 & MEMORY_REG_28__1__SCAN_IN); 
assign U1677 = ~(U1674 & MEMORY_REG_28__0__SCAN_IN); 
assign U1680 = ~(U1679 & MEMORY_REG_27__1__SCAN_IN); 
assign U1682 = ~(U1679 & MEMORY_REG_27__0__SCAN_IN); 
assign U1690 = ~(U1689 & MEMORY_REG_25__1__SCAN_IN); 
assign U1692 = ~(U1689 & MEMORY_REG_25__0__SCAN_IN); 
assign U1695 = ~(U1694 & MEMORY_REG_24__1__SCAN_IN); 
assign U1697 = ~(U1694 & MEMORY_REG_24__0__SCAN_IN); 
assign U1700 = ~(U1699 & MEMORY_REG_23__1__SCAN_IN); 
assign U1702 = ~(U1699 & MEMORY_REG_23__0__SCAN_IN); 
assign U1705 = ~(U1704 & MEMORY_REG_22__1__SCAN_IN); 
assign U1707 = ~(U1704 & MEMORY_REG_22__0__SCAN_IN); 
assign U1710 = ~(U1709 & MEMORY_REG_21__1__SCAN_IN); 
assign U1712 = ~(U1709 & MEMORY_REG_21__0__SCAN_IN); 
assign U1715 = ~(U1714 & MEMORY_REG_20__1__SCAN_IN); 
assign U1717 = ~(U1714 & MEMORY_REG_20__0__SCAN_IN); 
assign U1720 = ~(U1719 & MEMORY_REG_19__1__SCAN_IN); 
assign U1722 = ~(U1719 & MEMORY_REG_19__0__SCAN_IN); 
assign U1725 = ~(U1724 & MEMORY_REG_18__1__SCAN_IN); 
assign U1727 = ~(U1724 & MEMORY_REG_18__0__SCAN_IN); 
assign U1730 = ~(U1729 & MEMORY_REG_17__1__SCAN_IN); 
assign U1732 = ~(U1729 & MEMORY_REG_17__0__SCAN_IN); 
assign U1735 = ~(U1734 & MEMORY_REG_16__1__SCAN_IN); 
assign U1737 = ~(U1734 & MEMORY_REG_16__0__SCAN_IN); 
assign U1740 = ~(U1739 & MEMORY_REG_15__1__SCAN_IN); 
assign U1742 = ~(U1739 & MEMORY_REG_15__0__SCAN_IN); 
assign U1745 = ~(U1744 & MEMORY_REG_14__1__SCAN_IN); 
assign U1747 = ~(U1744 & MEMORY_REG_14__0__SCAN_IN); 
assign U1750 = ~(U1749 & MEMORY_REG_13__1__SCAN_IN); 
assign U1752 = ~(U1749 & MEMORY_REG_13__0__SCAN_IN); 
assign U1755 = ~(U1754 & MEMORY_REG_12__1__SCAN_IN); 
assign U1757 = ~(U1754 & MEMORY_REG_12__0__SCAN_IN); 
assign U1760 = ~(U1759 & MEMORY_REG_11__1__SCAN_IN); 
assign U1762 = ~(U1759 & MEMORY_REG_11__0__SCAN_IN); 
assign U1765 = ~(U1764 & MEMORY_REG_10__1__SCAN_IN); 
assign U1767 = ~(U1764 & MEMORY_REG_10__0__SCAN_IN); 
assign U1770 = ~(U1769 & MEMORY_REG_9__1__SCAN_IN); 
assign U1772 = ~(U1769 & MEMORY_REG_9__0__SCAN_IN); 
assign U1775 = ~(U1774 & MEMORY_REG_8__1__SCAN_IN); 
assign U1777 = ~(U1774 & MEMORY_REG_8__0__SCAN_IN); 
assign U1780 = ~(U1779 & MEMORY_REG_7__1__SCAN_IN); 
assign U1782 = ~(U1779 & MEMORY_REG_7__0__SCAN_IN); 
assign U1785 = ~(U1784 & MEMORY_REG_6__1__SCAN_IN); 
assign U1787 = ~(U1784 & MEMORY_REG_6__0__SCAN_IN); 
assign U1795 = ~(U1794 & MEMORY_REG_4__1__SCAN_IN); 
assign U1797 = ~(U1794 & MEMORY_REG_4__0__SCAN_IN); 
assign U1800 = ~(U1799 & MEMORY_REG_3__1__SCAN_IN); 
assign U1802 = ~(U1799 & MEMORY_REG_3__0__SCAN_IN); 
assign U1805 = ~(U1804 & MEMORY_REG_2__1__SCAN_IN); 
assign U1807 = ~(U1804 & MEMORY_REG_2__0__SCAN_IN); 
assign U1810 = ~(U1809 & MEMORY_REG_1__1__SCAN_IN); 
assign U1812 = ~(U1809 & MEMORY_REG_1__0__SCAN_IN); 
assign U1821 = ~(U1493 & U1820); 
assign U1823 = ~U1515; 
assign U1834 = ~(U1530 & U1504); 
assign U1868 = ~(U1615 & U1614 & U1635); 
assign U1899 = ~(U1320 & U1496); 
assign U1900 = ~(U1635 & U1492); 
assign U1902 = ~(U1320 & U1635); 
assign U1910 = ~(U1621 & U1539); 
assign U1912 = ~(U1612 & U1611); 
assign U1917 = ~(U1531 & U1916); 
assign U1919 = ~(U1882 & U1621); 
assign U1924 = ~(U1621 & U1618 & U1882); 
assign U1928 = ~(U1618 & U1539 & U1621); 
assign U1956 = ~(U1516 & U1955); 
assign U1957 = ~(U1318 & U1621); 
assign U1961 = ~(U1884 & U1559 & U1621); 
assign U1989 = ~(U1988 & U1987); 
assign U2009 = ~(U2161 & U2160 & U2008); 
assign U2014 = ~(U1306 & U1500); 
assign U2029 = ~(U1621 & U1612); 
assign U2031 = ~(U1320 & U1635); 
assign U2110 = ~(U1497 & U1493); 
assign U2134 = ~(U1306 & U1496); 
assign U2155 = ~(U1495 & U1500); 
assign U2169 = ~(U2109 & DATA_OUT_REG_1__SCAN_IN); 
assign U2170 = ~(U2166 & U1519); 
assign R730_U16 = ~(R730_U18 & MAX_REG_3__SCAN_IN); 
assign R730_U23 = ~(R730_U18 & R730_U10); 
assign R785_U16 = ~(R785_U18 & SCAN_REG_3__SCAN_IN); 
assign R785_U23 = ~(R785_U18 & R785_U10); 
assign U1305 = U1654 & U1819; 
assign U1310 = U1823 & U1622; 
assign U1371 = U1528 & U1495 & U1912; 
assign U1425 = ~(U1813 & U1812); 
assign U1426 = ~(U1811 & U1810); 
assign U1427 = ~(U1808 & U1807); 
assign U1428 = ~(U1806 & U1805); 
assign U1429 = ~(U1803 & U1802); 
assign U1430 = ~(U1801 & U1800); 
assign U1431 = ~(U1798 & U1797); 
assign U1432 = ~(U1796 & U1795); 
assign U1435 = ~(U1788 & U1787); 
assign U1436 = ~(U1786 & U1785); 
assign U1437 = ~(U1783 & U1782); 
assign U1438 = ~(U1781 & U1780); 
assign U1439 = ~(U1778 & U1777); 
assign U1440 = ~(U1776 & U1775); 
assign U1441 = ~(U1773 & U1772); 
assign U1442 = ~(U1771 & U1770); 
assign U1443 = ~(U1768 & U1767); 
assign U1444 = ~(U1766 & U1765); 
assign U1445 = ~(U1763 & U1762); 
assign U1446 = ~(U1761 & U1760); 
assign U1447 = ~(U1758 & U1757); 
assign U1448 = ~(U1756 & U1755); 
assign U1449 = ~(U1753 & U1752); 
assign U1450 = ~(U1751 & U1750); 
assign U1451 = ~(U1748 & U1747); 
assign U1452 = ~(U1746 & U1745); 
assign U1453 = ~(U1743 & U1742); 
assign U1454 = ~(U1741 & U1740); 
assign U1455 = ~(U1738 & U1737); 
assign U1456 = ~(U1736 & U1735); 
assign U1457 = ~(U1733 & U1732); 
assign U1458 = ~(U1731 & U1730); 
assign U1459 = ~(U1728 & U1727); 
assign U1460 = ~(U1726 & U1725); 
assign U1461 = ~(U1723 & U1722); 
assign U1462 = ~(U1721 & U1720); 
assign U1463 = ~(U1718 & U1717); 
assign U1464 = ~(U1716 & U1715); 
assign U1465 = ~(U1713 & U1712); 
assign U1466 = ~(U1711 & U1710); 
assign U1467 = ~(U1708 & U1707); 
assign U1468 = ~(U1706 & U1705); 
assign U1469 = ~(U1703 & U1702); 
assign U1470 = ~(U1701 & U1700); 
assign U1471 = ~(U1698 & U1697); 
assign U1472 = ~(U1696 & U1695); 
assign U1473 = ~(U1693 & U1692); 
assign U1474 = ~(U1691 & U1690); 
assign U1477 = ~(U1683 & U1682); 
assign U1478 = ~(U1681 & U1680); 
assign U1479 = ~(U1678 & U1677); 
assign U1480 = ~(U1676 & U1675); 
assign U1481 = ~(U1673 & U1672); 
assign U1482 = ~(U1671 & U1670); 
assign U1483 = ~(U1668 & U1667); 
assign U1484 = ~(U1666 & U1665); 
assign U1498 = ~(U1655 & U1614); 
assign U1524 = ~(U1654 & U1612); 
assign U1534 = ~(U1611 & U1500 & U1619); 
assign U1537 = ~(U1654 & U1618); 
assign U1542 = ~(U1650 & U1653); 
assign U1585 = U2042 & U2041 & U2040 & U2039 & U1584; 
assign U1587 = U2050 & U2049 & U2048 & U2047 & U1586; 
assign U1589 = U2058 & U2057 & U2056 & U2055 & U1588; 
assign U1591 = U2066 & U2065 & U2064 & U2063 & U1590; 
assign U1593 = U2074 & U2073 & U2072 & U2071 & U1592; 
assign U1595 = U2082 & U2081 & U2080 & U2079 & U1594; 
assign U1597 = U2090 & U2089 & U2088 & U2087 & U1596; 
assign U1599 = U2098 & U2097 & U2096 & U2095 & U1598; 
assign U1606 = ~(U1618 & U1500 & U1613); 
assign U1610 = ~U1503; 
assign U1623 = ~(U1651 & U1494); 
assign U1624 = ~(U1656 & U1635); 
assign U1626 = ~(U1619 & U1616); 
assign U1627 = ~U1526; 
assign U1631 = ~(U1619 & U1654); 
assign U1640 = ~(U1655 & U1500); 
assign U1643 = ~(U1613 & U1321); 
assign U1652 = ~U1528; 
assign U1822 = ~(U1614 & U1821 & U1622); 
assign U1827 = ~(U1621 & U1611 & U1655); 
assign U1831 = ~(U1503 & U1499); 
assign U1835 = ~(U1611 & U1834); 
assign U1901 = ~(U1899 & U1900 & U1898); 
assign U1918 = ~(U1917 & U1501); 
assign U1936 = ~(U1656 & U1618); 
assign U1962 = ~(U1960 & U1545 & U1961); 
assign U1964 = ~(U1528 & U1963); 
assign U1967 = ~(U1528 & U1530); 
assign U1991 = ~(U1989 & U1985); 
assign U1997 = ~(U1616 & U1493 & U1619); 
assign U2001 = ~(U1656 & U1494); 
assign U2003 = ~(U2155 & U2154 & U1612); 
assign U2015 = ~(U2014 & WR_REG_SCAN_IN); 
assign U2026 = ~(U1619 & U1615); 
assign U2027 = ~(U1614 & U1500 & U1619); 
assign U2132 = ~(U1655 & U1501 & U1492); 
assign U2135 = ~(U1613 & U1618); 
assign R745_U7 = ~U1380; 
assign R745_U10 = U1380 | U1379; 
assign R745_U13 = ~U1377; 
assign R745_U14 = ~U1378; 
assign R745_U17 = ~U1375; 
assign R745_U19 = ~U1376; 
assign R745_U26 = ~(U1379 & U1380); 
assign R730_U12 = ~(R730_U23 & R730_U22); 
assign R730_U19 = ~R730_U16; 
assign R730_U20 = ~(R730_U16 & MAX_REG_4__SCAN_IN); 
assign R785_U12 = ~(R785_U23 & R785_U22); 
assign R785_U19 = ~R785_U16; 
assign R785_U20 = ~(R785_U16 & SCAN_REG_4__SCAN_IN); 
assign U1389 = ~(U1599 & U1597 & U1595 & U1593); 
assign U1390 = ~(U1591 & U1589 & U1587 & U1585); 
assign U1392 = ~(U1606 & U2015); 
assign U1529 = ~(U1652 & U1616); 
assign U1548 = ~R745_U7; 
assign U1549 = ~(U1610 & U1492); 
assign U1562 = ~(U1991 & U1990); 
assign U1617 = ~U1498; 
assign U1620 = ~U1537; 
assign U1628 = ~U1534; 
assign U1629 = ~(U1305 & U1496); 
assign U1630 = ~U1524; 
assign U1825 = ~(U1823 & U1610); 
assign U1829 = ~(U1618 & U1492 & U1305); 
assign U1832 = ~(U1614 & U1831); 
assign U1851 = ~U1606; 
assign U1852 = ~(U1627 & U1622); 
assign U1865 = ~(U1621 & U1610); 
assign U1897 = ~(U2135 & U2134 & U2133 & U2132); 
assign U1903 = ~(U1611 & U1901); 
assign U1907 = ~(U1525 & U1537); 
assign U1914 = ~(U1371 & U1913); 
assign U1927 = ~U1542; 
assign U1937 = ~(U1936 & U1935 & U1371); 
assign U1951 = ~(U1612 & U1616 & U1864 & U1310); 
assign U1952 = ~(U1498 & U1623); 
assign U1958 = ~(U1542 & DATA_OUT_REG_1__SCAN_IN); 
assign U1965 = ~(U1615 & U1964); 
assign U2002 = ~(U1498 & U2001); 
assign U2011 = ~(U1621 & U1610); 
assign U2019 = ~(U1636 & U1640); 
assign U2022 = ~(U1310 & U1627); 
assign U2025 = ~(U1627 & U1515); 
assign U2030 = ~(U1610 & U1500); 
assign U2148 = ~(U1606 & DATA_IN_REG_1__SCAN_IN); 
assign U2150 = ~(U1606 & DATA_IN_REG_0__SCAN_IN); 
assign R745_U9 = ~(R745_U10 & R745_U26); 
assign R745_U20 = ~R745_U10; 
assign R745_U25 = ~(U1378 & R745_U10); 
assign R730_U21 = ~(R730_U19 & R730_U15); 
assign R785_U21 = ~(R785_U19 & R785_U15); 
assign U1368 = U1549 & U1822; 
assign U1538 = ~(U1620 & U1494); 
assign U1551 = ~(U1646 & U1965); 
assign U1555 = ~(U1562 & U1993); 
assign U1561 = ~(U1524 & U1529); 
assign U1600 = ~(U1539 & U1501 & U1628); 
assign U1633 = ~U1529; 
assign U1634 = ~(U1616 & U1617); 
assign U1637 = ~(U1864 & U1630 & U1310); 
assign U1638 = ~(U1630 & U1536 & U1310); 
assign U1641 = ~(U1622 & U1515 & U1630); 
assign U1645 = ~(U1628 & U1501 & U2009); 
assign U1648 = ~(U1615 & U1617); 
assign U1657 = ~U1549; 
assign U1826 = ~(U1824 & U1530 & U1825); 
assign U1894 = ~(U1611 & U1548); 
assign U1904 = ~(U1616 & U1897); 
assign U1909 = ~(U1622 & U1907); 
assign U1915 = ~(U1914 & U1501); 
assign U1929 = ~(U1622 & U1907); 
assign U1938 = ~(U1622 & U1937); 
assign U1953 = ~(U1622 & U1952); 
assign U1959 = ~(U1958 & U1957); 
assign U1992 = ~U1562; 
assign U2004 = ~(U2002 & U1493); 
assign U2005 = ~(U1628 & U1492); 
assign U2010 = ~(U1628 & U1622); 
assign U2021 = ~(U1611 & U2019); 
assign U2028 = ~(U1628 & U1501); 
assign U2033 = ~(U2170 & U2169 & U1628); 
assign U2111 = ~(U1864 & U1630); 
assign U2149 = ~(U1851 & NUM_REG_1__SCAN_IN); 
assign U2151 = ~(U1851 & NUM_REG_0__SCAN_IN); 
assign R745_U11 = ~(R745_U20 & R745_U14); 
assign R730_U11 = ~(R730_U21 & R730_U20); 
assign R785_U11 = ~(R785_U21 & R785_U20); 
assign U1311 = U1993 & U1992 & PLAY_REG_SCAN_IN; 
assign U1314 = U2110 & U1551; 
assign U1315 = U1967 & U1551; 
assign U1522 = ~(U1650 & U1832 & U1634); 
assign U1527 = ~(U1606 & U1852 & U1641); 
assign U1532 = ~(U1638 & U1865); 
assign U1543 = ~(U1927 & U1928 & U1929); 
assign U1560 = ~(U1534 & U1538); 
assign U1572 = ~(U2149 & U2148); 
assign U1573 = ~(U2151 & U2150); 
assign U1579 = U1903 & U1902 & U1648 & U1637; 
assign U1580 = U1495 & U1641 & U1631 & U1629; 
assign U1581 = U1626 & U1624 & U1629 & U1640 & U1634; 
assign U1608 = ~(U2010 & U2011 & U1645); 
assign U1632 = ~U1538; 
assign U1642 = ~(U1657 & U1616); 
assign U1644 = ~(U1633 & U1310); 
assign U1828 = ~(U1616 & U1622 & U1826); 
assign U1867 = ~(U1633 & U1515); 
assign U1883 = ~U1600; 
assign U1895 = ~U1561; 
assign U1896 = ~(U1561 & U1501); 
assign U1911 = ~(U1653 & U1908 & U1649 & U1910 & U1909); 
assign U1920 = ~(U1918 & U1919 & U1915); 
assign U1926 = ~(U1924 & U1925 & U1915); 
assign U1966 = ~U1551; 
assign U1994 = ~U1555; 
assign U1998 = ~(U1538 & U1629 & U1997); 
assign U2006 = ~(U2005 & U2003 & U2004); 
assign U2013 = ~(U1555 & PLAY_REG_SCAN_IN & SPEAKER_REG_SCAN_IN); 
assign U2023 = ~(U1526 & U1538); 
assign U2124 = ~(U1600 & IND_REG_1__SCAN_IN); 
assign U2126 = ~(U1600 & IND_REG_0__SCAN_IN); 
assign R745_U6 = ~(R745_U11 & R745_U25); 
assign R745_U21 = ~R745_U11; 
assign R745_U24 = ~(U1377 & R745_U11); 
assign U1316 = U1616 & U1515 & U1527; 
assign U1317 = U1611 & U1532; 
assign U1369 = U1534 & U1867; 
assign U1370 = U1644 & U1896; 
assign U1372 = U1951 & U1600 & U1648 & U1644; 
assign U1381 = U1311 & U2113; 
assign U1382 = U1311 & U2175; 
assign U1383 = U1311 & U1553; 
assign U1582 = U1643 & U1642 & U1645 & U1581; 
assign U1583 = U1634 & U1626 & U1638 & U1549 & U1644; 
assign U1658 = ~(U1556 & U1994 & PLAY_REG_SCAN_IN); 
assign U1830 = ~(U1827 & U1648 & U1828 & U1368 & U1829); 
assign U1833 = ~U1522; 
assign U1853 = ~U1527; 
assign U1866 = ~U1532; 
assign U1905 = ~(U1632 & U1492); 
assign U1922 = ~(U1911 & TIMEBASE_REG_5__SCAN_IN); 
assign U1930 = ~U1543; 
assign U1940 = ~(U1543 & TIMEBASE_REG_3__SCAN_IN); 
assign U1948 = ~(R745_U7 & U1920); 
assign U1949 = ~(U1911 & TIMEBASE_REG_0__SCAN_IN); 
assign U1968 = ~(U1315 & MAX_REG_4__SCAN_IN); 
assign U1969 = ~(U1314 & SCAN_REG_4__SCAN_IN); 
assign U1970 = ~(U1966 & ADDRESS_REG_4__SCAN_IN); 
assign U1971 = ~(U1315 & MAX_REG_3__SCAN_IN); 
assign U1972 = ~(U1314 & SCAN_REG_3__SCAN_IN); 
assign U1973 = ~(U1966 & ADDRESS_REG_3__SCAN_IN); 
assign U1974 = ~(U1315 & MAX_REG_2__SCAN_IN); 
assign U1975 = ~(U1314 & SCAN_REG_2__SCAN_IN); 
assign U1976 = ~(U1966 & ADDRESS_REG_2__SCAN_IN); 
assign U1977 = ~(U1315 & MAX_REG_1__SCAN_IN); 
assign U1978 = ~(U1314 & SCAN_REG_1__SCAN_IN); 
assign U1979 = ~(U1966 & ADDRESS_REG_1__SCAN_IN); 
assign U1980 = ~(U1315 & MAX_REG_0__SCAN_IN); 
assign U1981 = ~(U1314 & SCAN_REG_0__SCAN_IN); 
assign U1982 = ~(U1966 & ADDRESS_REG_0__SCAN_IN); 
assign U1995 = ~(U1994 & PLAY_REG_SCAN_IN); 
assign U1999 = ~(U1622 & U1998); 
assign U2012 = ~U1608; 
assign U2017 = ~U1560; 
assign U2018 = ~(U1622 & U1560); 
assign U2024 = ~(U2023 & U1501); 
assign U2034 = ~(U1895 & U2033 & U1634 & U1623); 
assign U2125 = ~(U1883 & U1318); 
assign U2127 = ~(U1884 & U1559 & U1883); 
assign U2131 = ~(U1894 & U1532); 
assign U2163 = ~(U1611 & U1608); 
assign R745_U12 = ~(R745_U21 & R745_U13); 
assign U1309 = U1834 & U1611 & U1830; 
assign U1319 = U1522 & U1830; 
assign U1373 = U1631 & U2024; 
assign U1384 = ~(U2018 & U1637 & U1492); 
assign U1393 = ~(U1658 & U2013); 
assign U1395 = ~(U1981 & U1980 & U1982); 
assign U1396 = ~(U1978 & U1977 & U1979); 
assign U1397 = ~(U1975 & U1974 & U1976); 
assign U1398 = ~(U1972 & U1971 & U1973); 
assign U1399 = ~(U1969 & U1968 & U1970); 
assign U1541 = ~(U1905 & U1904 & U1370 & U1579); 
assign U1564 = ~(U2125 & U2124); 
assign U1565 = ~(U2127 & U2126); 
assign U1604 = ~(U1953 & U1642 & U1372); 
assign U1607 = ~(U1368 & U1999 & U1372); 
assign U1639 = ~(U1819 & U1651 & U1830); 
assign U1836 = ~(U1835 & U1833 & U1830); 
assign U1854 = ~(R785_U11 & U1316); 
assign U1855 = ~(U1853 & SCAN_REG_4__SCAN_IN); 
assign U1856 = ~(R785_U12 & U1316); 
assign U1857 = ~(U1853 & SCAN_REG_3__SCAN_IN); 
assign U1858 = ~(R785_U13 & U1316); 
assign U1859 = ~(U1853 & SCAN_REG_2__SCAN_IN); 
assign U1860 = ~(R785_U14 & U1316); 
assign U1861 = ~(U1853 & SCAN_REG_1__SCAN_IN); 
assign U1862 = ~(R785_U5 & U1316); 
assign U1863 = ~(U1853 & SCAN_REG_0__SCAN_IN); 
assign U1869 = ~(U1369 & U1868); 
assign U1887 = ~(U1866 & TIMEBASE_REG_4__SCAN_IN); 
assign U1889 = ~(U1866 & TIMEBASE_REG_3__SCAN_IN); 
assign U1890 = ~(R745_U6 & U1317); 
assign U1891 = ~(U1866 & TIMEBASE_REG_2__SCAN_IN); 
assign U1892 = ~(R745_U9 & U1317); 
assign U1893 = ~(U1866 & TIMEBASE_REG_1__SCAN_IN); 
assign U1931 = ~(U1930 & U1649); 
assign U1950 = ~(U1949 & U1948); 
assign U1996 = ~(U1995 & S_REG_SCAN_IN); 
assign U2020 = ~(U2017 & U1524); 
assign U2032 = ~(U1626 & U1624 & U1629 & U2031 & U1369); 
assign U2128 = ~(U1866 & TIMEBASE_REG_5__SCAN_IN); 
assign U2130 = ~(U1866 & TIMEBASE_REG_0__SCAN_IN); 
assign U2162 = ~(U2012 & NLOSS_REG_SCAN_IN); 
assign U2172 = ~(U2034 & U1501); 
assign R745_U8 = ~(R745_U12 & R745_U24); 
assign R745_U22 = ~R745_U12; 
assign R745_U29 = ~(U1376 & R745_U12); 
assign U1322 = U1926 & U1541; 
assign U1323 = U1931 & U1541; 
assign U1374 = U2026 & U2027 & U2025 & U1373; 
assign U1386 = ~(U1373 & U1370 & U1582); 
assign U1394 = ~(U1658 & U1996); 
assign U1405 = ~(U1893 & U1892); 
assign U1406 = ~(U1891 & U1890); 
assign U1414 = ~(U1863 & U1862); 
assign U1415 = ~(U1861 & U1860); 
assign U1416 = ~(U1859 & U1858); 
assign U1417 = ~(U1857 & U1856); 
assign U1418 = ~(U1855 & U1854); 
assign U1567 = ~(U2131 & U2130); 
assign U1575 = ~(U2163 & U2162); 
assign U1647 = ~(U1621 & U1496 & U1541); 
assign U1838 = ~(U1309 & IND_REG_1__SCAN_IN & IND_REG_0__SCAN_IN); 
assign U1839 = ~(U1319 & U1837); 
assign U1840 = ~(U1836 & NL_REG_3__SCAN_IN); 
assign U1841 = ~(U1520 & U1319 & DATA_OUT_REG_1__SCAN_IN); 
assign U1842 = ~(U1517 & U1309 & IND_REG_1__SCAN_IN); 
assign U1843 = ~(U1836 & NL_REG_2__SCAN_IN); 
assign U1845 = ~(U1518 & U1309 & IND_REG_0__SCAN_IN); 
assign U1846 = ~(U1844 & U1319); 
assign U1847 = ~(U1836 & NL_REG_1__SCAN_IN); 
assign U1848 = ~(U1519 & U1520 & U1319); 
assign U1849 = ~(U1517 & U1518 & U1309); 
assign U1850 = ~(U1836 & NL_REG_0__SCAN_IN); 
assign U1870 = ~(U1622 & U1869); 
assign U1888 = ~(R745_U8 & U1317); 
assign U1906 = ~U1541; 
assign U1939 = ~(R745_U8 & U1926); 
assign U1954 = ~U1604; 
assign U2000 = ~U1607; 
assign U2112 = ~(U2020 & U1501); 
assign U2141 = ~(U1950 & U1541); 
assign U2143 = ~(U1956 & U1604); 
assign U2145 = ~(U1959 & U1604); 
assign U2147 = ~(U1962 & U1604); 
assign U2157 = ~(U2006 & U1607); 
assign U2171 = ~(U1622 & U2032); 
assign R745_U18 = ~(R745_U22 & R745_U19); 
assign R745_U30 = ~(R745_U22 & R745_U19); 
assign U1385 = ~(U2022 & U2021 & U1580 & U2112 & U2111); 
assign U1387 = ~(U2029 & U2030 & U2028 & U1583 & U1374); 
assign U1388 = ~(U1646 & U1643 & U1374 & U2172 & U2171); 
assign U1407 = ~(U1889 & U1888); 
assign U1419 = ~(U1850 & U1849 & U1848 & U1639); 
assign U1420 = ~(U1847 & U1846 & U1845 & U1639); 
assign U1421 = ~(U1843 & U1842 & U1841 & U1639); 
assign U1422 = ~(U1840 & U1839 & U1838 & U1639); 
assign U1533 = ~(U1866 & U1870); 
assign U1932 = ~(U1323 & TIMEBASE_REG_4__SCAN_IN); 
assign U1934 = ~(U1906 & COUNT_REG2_4__SCAN_IN); 
assign U1941 = ~(U1940 & U1938 & U1939); 
assign U1942 = ~(U1323 & TIMEBASE_REG_2__SCAN_IN); 
assign U1943 = ~(U1322 & R745_U6); 
assign U1944 = ~(U1906 & COUNT_REG2_2__SCAN_IN); 
assign U1945 = ~(U1323 & TIMEBASE_REG_1__SCAN_IN); 
assign U1946 = ~(U1322 & R745_U9); 
assign U1947 = ~(U1906 & COUNT_REG2_1__SCAN_IN); 
assign U2136 = ~(U1906 & COUNT_REG2_5__SCAN_IN); 
assign U2138 = ~(U1906 & COUNT_REG2_3__SCAN_IN); 
assign U2140 = ~(U1906 & COUNT_REG2_0__SCAN_IN); 
assign U2142 = ~(U1954 & SOUND_REG_2__SCAN_IN); 
assign U2144 = ~(U1954 & SOUND_REG_1__SCAN_IN); 
assign U2146 = ~(U1954 & SOUND_REG_0__SCAN_IN); 
assign U2156 = ~(U2000 & PLAY_REG_SCAN_IN); 
assign R745_U16 = ~(R745_U30 & R745_U29); 
assign R745_U23 = ~R745_U18; 
assign R745_U27 = ~(U1375 & R745_U18); 
assign U1313 = U1616 & U1533; 
assign U1400 = ~(U2141 & U2140 & U1647); 
assign U1401 = ~(U1946 & U1945 & U1947); 
assign U1402 = ~(U1943 & U1942 & U1944); 
assign U1569 = ~(U2143 & U2142); 
assign U1570 = ~(U2145 & U2144); 
assign U1571 = ~(U2147 & U2146); 
assign U1574 = ~(U2157 & U2156); 
assign U1871 = ~U1533; 
assign U1886 = ~(R745_U16 & U1317); 
assign U1933 = ~(U1322 & R745_U16); 
assign U2139 = ~(U1941 & U1541); 
assign R745_U28 = ~(R745_U23 & R745_U17); 
assign U1403 = ~(U1933 & U1932 & U1934); 
assign U1408 = ~(U1887 & U1886); 
assign U1568 = ~(U2139 & U2138); 
assign U1872 = ~(R730_U11 & U1313); 
assign U1873 = ~(U1871 & MAX_REG_4__SCAN_IN); 
assign U1874 = ~(R730_U12 & U1313); 
assign U1875 = ~(U1871 & MAX_REG_3__SCAN_IN); 
assign U1876 = ~(R730_U13 & U1313); 
assign U1877 = ~(U1871 & MAX_REG_2__SCAN_IN); 
assign U1878 = ~(R730_U14 & U1313); 
assign U1879 = ~(U1871 & MAX_REG_1__SCAN_IN); 
assign U1880 = ~(R730_U5 & U1313); 
assign U1881 = ~(U1871 & MAX_REG_0__SCAN_IN); 
assign R745_U15 = ~(R745_U28 & R745_U27); 
assign U1409 = ~(U1881 & U1880); 
assign U1410 = ~(U1879 & U1878); 
assign U1411 = ~(U1877 & U1876); 
assign U1412 = ~(U1875 & U1874); 
assign U1413 = ~(U1873 & U1872); 
assign U1540 = ~R745_U15; 
assign U1921 = ~(R745_U15 & U1920); 
assign U1885 = ~(U1611 & U1540); 
assign U1923 = ~(U1922 & U1921); 
assign U2129 = ~(U1885 & U1532); 
assign U2137 = ~(U1923 & U1541); 
assign U1404 = ~(U2137 & U2136 & U1647); 
assign U1566 = ~(U2129 & U2128); 
endmodule 
