module b06_C( EQL, CONT_EQL, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, U55, U56, U57, U58, U59, U60, U61, U62); 
input EQL, CONT_EQL, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN; 
output U55, U56, U57, U58, U59, U60, U61, U62; 
wire U54, U63, U64, U65, U66, U67, U68, U69, U70, U71, U72, U73, U74, U75, U76, U77, U78, U79, U80, U81, U82, U83, U84, U85, U86, U87, U88, U89, U90, U91, U92; 
assign U63 = STATE_REG_2__SCAN_IN & STATE_REG_1__SCAN_IN & STATE_REG_0__SCAN_IN; 
assign U64 = ~STATE_REG_1__SCAN_IN; 
assign U65 = ~EQL; 
assign U66 = ~(EQL & STATE_REG_1__SCAN_IN); 
assign U67 = ~STATE_REG_2__SCAN_IN; 
assign U68 = ~STATE_REG_0__SCAN_IN; 
assign U69 = STATE_REG_2__SCAN_IN | STATE_REG_0__SCAN_IN; 
assign U76 = ~(STATE_REG_2__SCAN_IN & STATE_REG_1__SCAN_IN); 
assign U77 = STATE_REG_1__SCAN_IN | STATE_REG_0__SCAN_IN; 
assign U88 = ~(STATE_REG_2__SCAN_IN & STATE_REG_0__SCAN_IN); 
assign U90 = ~(STATE_REG_1__SCAN_IN & STATE_REG_0__SCAN_IN); 
assign U70 = ~(U64 & U67 & STATE_REG_0__SCAN_IN); 
assign U71 = ~U66; 
assign U72 = ~(U68 & U64 & U65 & STATE_REG_2__SCAN_IN); 
assign U73 = ~U69; 
assign U78 = ~(U65 & U77); 
assign U81 = ~(EQL & U67 & STATE_REG_0__SCAN_IN); 
assign U84 = CONT_EQL | U63; 
assign U87 = ~(EQL & U68); 
assign U91 = ~(EQL & U64); 
assign U74 = ~U70; 
assign U75 = ~(U71 & STATE_REG_2__SCAN_IN); 
assign U80 = ~(U78 & STATE_REG_2__SCAN_IN); 
assign U82 = ~(U73 & STATE_REG_1__SCAN_IN); 
assign U83 = ~(U65 & U73 & STATE_REG_1__SCAN_IN); 
assign U85 = ~(U71 & U68); 
assign U86 = ~(U78 & STATE_REG_2__SCAN_IN); 
assign U89 = ~(U73 & U64); 
assign U92 = ~(U87 & STATE_REG_1__SCAN_IN); 
assign U54 = U90 & U89; 
assign U56 = ~(U82 & U81 & U72 & U66); 
assign U58 = ~(U88 & U69 & U92 & U91); 
assign U59 = ~(U86 & U70 & U85); 
assign U61 = ~(U72 & U75); 
assign U62 = ~(U84 & U83); 
assign U79 = ~(U74 & U65); 
assign U55 = ~(U54 & U78); 
assign U57 = ~(U80 & U79); 
assign U60 = ~(EQL & U76 & U54); 
endmodule 
