module b13_C( EOC, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_, DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_, DSR, TX_END_REG_SCAN_IN, S2_REG_0__SCAN_IN, S2_REG_1__SCAN_IN, CANALE_REG_3__SCAN_IN, CANALE_REG_2__SCAN_IN, CANALE_REG_1__SCAN_IN, CANALE_REG_0__SCAN_IN, CONTA_TMP_REG_3__SCAN_IN, CONTA_TMP_REG_2__SCAN_IN, CONTA_TMP_REG_1__SCAN_IN, CONTA_TMP_REG_0__SCAN_IN, ITFC_STATE_REG_1__SCAN_IN, ITFC_STATE_REG_0__SCAN_IN, OUT_REG_REG_7__SCAN_IN, OUT_REG_REG_6__SCAN_IN, OUT_REG_REG_5__SCAN_IN, OUT_REG_REG_4__SCAN_IN, OUT_REG_REG_3__SCAN_IN, OUT_REG_REG_2__SCAN_IN, OUT_REG_REG_1__SCAN_IN, OUT_REG_REG_0__SCAN_IN, NEXT_BIT_REG_3__SCAN_IN, NEXT_BIT_REG_2__SCAN_IN, NEXT_BIT_REG_1__SCAN_IN, NEXT_BIT_REG_0__SCAN_IN, TX_CONTA_REG_9__SCAN_IN, TX_CONTA_REG_8__SCAN_IN, TX_CONTA_REG_7__SCAN_IN, TX_CONTA_REG_6__SCAN_IN, TX_CONTA_REG_5__SCAN_IN, TX_CONTA_REG_4__SCAN_IN, TX_CONTA_REG_3__SCAN_IN, TX_CONTA_REG_2__SCAN_IN, TX_CONTA_REG_1__SCAN_IN, TX_CONTA_REG_0__SCAN_IN, LOAD_REG_SCAN_IN, SEND_DATA_REG_SCAN_IN, SEND_EN_REG_SCAN_IN, MUX_EN_REG_SCAN_IN, TRE_REG_SCAN_IN, LOAD_DATO_REG_SCAN_IN, SOC_REG_SCAN_IN, SEND_REG_SCAN_IN, MPX_REG_SCAN_IN, CONFIRM_REG_SCAN_IN, SHOT_REG_SCAN_IN, ADD_MPX2_REG_SCAN_IN, RDY_REG_SCAN_IN, ERROR_REG_SCAN_IN, S1_REG_2__SCAN_IN, S1_REG_1__SCAN_IN, S1_REG_0__SCAN_IN, U380, U381, U382, U383, U384, U385, U386, U387, U388, U389, U390, U391, U392, U393, U394, U395, U396, U397, U398, U399, U400, U401, U402, U403, U404, U405, U406, U407, U408, U409, U410, U411, U412, U413, U414, U415, U416, U417, U450, U451, U452, U453, U454, U455, U456, U457, U458, U459, U460, U461, U462, U463, U464); 
input EOC, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_, DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_, DSR, TX_END_REG_SCAN_IN, S2_REG_0__SCAN_IN, S2_REG_1__SCAN_IN, CANALE_REG_3__SCAN_IN, CANALE_REG_2__SCAN_IN, CANALE_REG_1__SCAN_IN, CANALE_REG_0__SCAN_IN, CONTA_TMP_REG_3__SCAN_IN, CONTA_TMP_REG_2__SCAN_IN, CONTA_TMP_REG_1__SCAN_IN, CONTA_TMP_REG_0__SCAN_IN, ITFC_STATE_REG_1__SCAN_IN, ITFC_STATE_REG_0__SCAN_IN, OUT_REG_REG_7__SCAN_IN, OUT_REG_REG_6__SCAN_IN, OUT_REG_REG_5__SCAN_IN, OUT_REG_REG_4__SCAN_IN, OUT_REG_REG_3__SCAN_IN, OUT_REG_REG_2__SCAN_IN, OUT_REG_REG_1__SCAN_IN, OUT_REG_REG_0__SCAN_IN, NEXT_BIT_REG_3__SCAN_IN, NEXT_BIT_REG_2__SCAN_IN, NEXT_BIT_REG_1__SCAN_IN, NEXT_BIT_REG_0__SCAN_IN, TX_CONTA_REG_9__SCAN_IN, TX_CONTA_REG_8__SCAN_IN, TX_CONTA_REG_7__SCAN_IN, TX_CONTA_REG_6__SCAN_IN, TX_CONTA_REG_5__SCAN_IN, TX_CONTA_REG_4__SCAN_IN, TX_CONTA_REG_3__SCAN_IN, TX_CONTA_REG_2__SCAN_IN, TX_CONTA_REG_1__SCAN_IN, TX_CONTA_REG_0__SCAN_IN, LOAD_REG_SCAN_IN, SEND_DATA_REG_SCAN_IN, SEND_EN_REG_SCAN_IN, MUX_EN_REG_SCAN_IN, TRE_REG_SCAN_IN, LOAD_DATO_REG_SCAN_IN, SOC_REG_SCAN_IN, SEND_REG_SCAN_IN, MPX_REG_SCAN_IN, CONFIRM_REG_SCAN_IN, SHOT_REG_SCAN_IN, ADD_MPX2_REG_SCAN_IN, RDY_REG_SCAN_IN, ERROR_REG_SCAN_IN, S1_REG_2__SCAN_IN, S1_REG_1__SCAN_IN, S1_REG_0__SCAN_IN; 
output U380, U381, U382, U383, U384, U385, U386, U387, U388, U389, U390, U391, U392, U393, U394, U395, U396, U397, U398, U399, U400, U401, U402, U403, U404, U405, U406, U407, U408, U409, U410, U411, U412, U413, U414, U415, U416, U417, U450, U451, U452, U453, U454, U455, U456, U457, U458, U459, U460, U461, U462, U463, U464; 
wire U375, U376, U377, U378, U379, U418, U419, U420, U421, U422, U423, U424, U425, U426, U427, U428, U429, U430, U431, U432, U433, U434, U435, U436, U437, U438, U439, U440, U441, U442, U443, U444, U445, U446, U447, U448, U449, U465, U466, U467, U468, U469, U470, U471, U472, U473, U474, U475, U476, U477, U478, U479, U480, U481, U482, U483, U484, U485, U486, U487, U488, U489, U490, U491, U492, U493, U494, U495, U496, U497, U498, U499, U500, U501, U502, U503, U504, U505, U506, U507, U508, U509, U510, U511, U512, U513, U514, U515, U516, U517, U518, U519, U520, U521, U522, U523, U524, U525, U526, U527, U528, U529, U530, U531, U532, U533, U534, U535, U536, U537, U538, U539, U540, U541, U542, U543, U544, U545, U546, U547, U548, U549, U550, U551, U552, U553, U554, U555, U556, U557, U558, U559, U560, U561, U562, U563, U564, U565, U566, U567, U568, U569, U570, U571, U572, U573, U574, U575, U576, U577, U578, U579, U580, U581, U582, U583, U584, U585, U586, U587, U588, U589, U590, U591, U592, U593, U594, U595, U596, U597, U598, U599, U600, U601, U602, U603, U604, U605, ADD_291_U5, ADD_291_U6, ADD_291_U7, ADD_291_U8, ADD_291_U9, ADD_291_U10, ADD_291_U11, ADD_291_U12, ADD_291_U13, ADD_291_U14, ADD_291_U15, ADD_291_U16, ADD_291_U17, ADD_291_U18, ADD_291_U19, ADD_291_U20, ADD_291_U21, ADD_291_U22, ADD_291_U23, ADD_291_U24, ADD_291_U25, ADD_291_U26, ADD_291_U27, ADD_291_U28, ADD_291_U29, ADD_291_U30, ADD_291_U31, ADD_291_U32, ADD_291_U33, ADD_291_U34, ADD_291_U35, ADD_291_U36, ADD_291_U37, ADD_291_U38, ADD_291_U39, ADD_291_U40, ADD_291_U41, ADD_291_U42, ADD_291_U43, ADD_291_U44, ADD_291_U45, ADD_291_U46, ADD_291_U47, ADD_291_U48, ADD_291_U49, ADD_291_U50, ADD_291_U51, ADD_291_U52, ADD_291_U53, ADD_291_U54, ADD_291_U55, ADD_291_U56, ADD_291_U57, GT_255_U6, GT_255_U7, GT_255_U8, GT_255_U9, GT_255_U10; 
assign U377 = NEXT_BIT_REG_2__SCAN_IN & NEXT_BIT_REG_1__SCAN_IN; 
assign U379 = CONTA_TMP_REG_1__SCAN_IN & CONTA_TMP_REG_0__SCAN_IN; 
assign U392 = LOAD_REG_SCAN_IN | TRE_REG_SCAN_IN | TX_END_REG_SCAN_IN; 
assign U418 = ~CONTA_TMP_REG_0__SCAN_IN; 
assign U419 = ~SEND_EN_REG_SCAN_IN; 
assign U422 = ~NEXT_BIT_REG_0__SCAN_IN; 
assign U424 = NEXT_BIT_REG_3__SCAN_IN | NEXT_BIT_REG_2__SCAN_IN; 
assign U425 = ~ITFC_STATE_REG_0__SCAN_IN; 
assign U426 = ~LOAD_REG_SCAN_IN; 
assign U427 = ~S1_REG_0__SCAN_IN; 
assign U428 = ~S1_REG_1__SCAN_IN; 
assign U429 = ~S1_REG_2__SCAN_IN; 
assign U430 = ~RDY_REG_SCAN_IN; 
assign U431 = ~(RDY_REG_SCAN_IN & S1_REG_1__SCAN_IN); 
assign U432 = ~SEND_REG_SCAN_IN; 
assign U433 = ~TRE_REG_SCAN_IN; 
assign U435 = ~ITFC_STATE_REG_1__SCAN_IN; 
assign U436 = ~S2_REG_1__SCAN_IN; 
assign U437 = ~CONFIRM_REG_SCAN_IN; 
assign U438 = ~MPX_REG_SCAN_IN; 
assign U440 = ~TX_END_REG_SCAN_IN; 
assign U441 = ~S2_REG_0__SCAN_IN; 
assign U442 = ~CONTA_TMP_REG_1__SCAN_IN; 
assign U445 = ~NEXT_BIT_REG_1__SCAN_IN; 
assign U446 = ~NEXT_BIT_REG_2__SCAN_IN; 
assign U447 = ~NEXT_BIT_REG_3__SCAN_IN; 
assign U449 = ~EOC; 
assign U485 = ~(S1_REG_2__SCAN_IN & S1_REG_1__SCAN_IN & S1_REG_0__SCAN_IN); 
assign U487 = ~(DSR & TRE_REG_SCAN_IN & SEND_REG_SCAN_IN); 
assign U490 = S1_REG_2__SCAN_IN | S1_REG_1__SCAN_IN | S1_REG_0__SCAN_IN; 
assign U500 = ITFC_STATE_REG_1__SCAN_IN | ITFC_STATE_REG_0__SCAN_IN; 
assign U501 = ~(ITFC_STATE_REG_1__SCAN_IN & ITFC_STATE_REG_0__SCAN_IN & TX_END_REG_SCAN_IN); 
assign U508 = ~(DSR & TRE_REG_SCAN_IN); 
assign U523 = ~(ITFC_STATE_REG_1__SCAN_IN & TX_END_REG_SCAN_IN); 
assign U524 = ~(ITFC_STATE_REG_0__SCAN_IN & TX_END_REG_SCAN_IN); 
assign U530 = NEXT_BIT_REG_2__SCAN_IN | NEXT_BIT_REG_1__SCAN_IN; 
assign U553 = ~(OUT_REG_REG_0__SCAN_IN & NEXT_BIT_REG_3__SCAN_IN); 
assign U558 = ~(OUT_REG_REG_1__SCAN_IN & NEXT_BIT_REG_3__SCAN_IN); 
assign U561 = ~(S1_REG_2__SCAN_IN & S1_REG_0__SCAN_IN); 
assign U563 = EOC | S1_REG_1__SCAN_IN; 
assign U568 = ~(LOAD_REG_SCAN_IN & TRE_REG_SCAN_IN); 
assign ADD_291_U5 = ~TX_CONTA_REG_0__SCAN_IN; 
assign ADD_291_U6 = ~TX_CONTA_REG_1__SCAN_IN; 
assign ADD_291_U7 = ~(TX_CONTA_REG_1__SCAN_IN & TX_CONTA_REG_0__SCAN_IN); 
assign ADD_291_U8 = ~TX_CONTA_REG_2__SCAN_IN; 
assign ADD_291_U10 = ~TX_CONTA_REG_3__SCAN_IN; 
assign ADD_291_U12 = ~TX_CONTA_REG_4__SCAN_IN; 
assign ADD_291_U14 = ~TX_CONTA_REG_5__SCAN_IN; 
assign ADD_291_U16 = ~TX_CONTA_REG_6__SCAN_IN; 
assign ADD_291_U18 = ~TX_CONTA_REG_7__SCAN_IN; 
assign ADD_291_U20 = ~TX_CONTA_REG_8__SCAN_IN; 
assign ADD_291_U30 = ~TX_CONTA_REG_9__SCAN_IN; 
assign GT_255_U9 = TX_CONTA_REG_2__SCAN_IN | TX_CONTA_REG_1__SCAN_IN | TX_CONTA_REG_0__SCAN_IN; 
assign U378 = U446 & NEXT_BIT_REG_1__SCAN_IN; 
assign U434 = ~(U427 & S1_REG_1__SCAN_IN); 
assign U439 = ~(U441 & CONFIRM_REG_SCAN_IN & S2_REG_1__SCAN_IN); 
assign U448 = ~(U445 & NEXT_BIT_REG_2__SCAN_IN); 
assign U465 = ~(U433 & LOAD_REG_SCAN_IN); 
assign U472 = ~(U441 & U436 & SEND_DATA_REG_SCAN_IN); 
assign U473 = ~U424; 
assign U477 = ~(U419 & TX_CONTA_REG_1__SCAN_IN); 
assign U479 = ~(U419 & TX_CONTA_REG_0__SCAN_IN); 
assign U480 = ~(U435 & ITFC_STATE_REG_0__SCAN_IN); 
assign U481 = ~(U425 & U435 & SHOT_REG_SCAN_IN); 
assign U483 = ~U431; 
assign U488 = ~(U440 & SEND_EN_REG_SCAN_IN); 
assign U489 = ~(U428 & U449 & S1_REG_2__SCAN_IN & S1_REG_0__SCAN_IN); 
assign U495 = ~(U425 & ITFC_STATE_REG_1__SCAN_IN); 
assign U497 = ~(U435 & ITFC_STATE_REG_0__SCAN_IN); 
assign U502 = ~(U500 & CONFIRM_REG_SCAN_IN); 
assign U503 = ~(U441 & U437 & S2_REG_1__SCAN_IN); 
assign U505 = ~(U436 & S2_REG_0__SCAN_IN); 
assign U509 = ~(U379 & CONTA_TMP_REG_2__SCAN_IN); 
assign U525 = ~(U524 & ITFC_STATE_REG_1__SCAN_IN); 
assign U526 = ~(U425 & SHOT_REG_SCAN_IN); 
assign U531 = ~(U530 & U422); 
assign U534 = ~(U419 & TX_CONTA_REG_9__SCAN_IN); 
assign U536 = ~(U419 & TX_CONTA_REG_8__SCAN_IN); 
assign U538 = ~(U419 & TX_CONTA_REG_7__SCAN_IN); 
assign U540 = ~(U419 & TX_CONTA_REG_6__SCAN_IN); 
assign U542 = ~(U419 & TX_CONTA_REG_5__SCAN_IN); 
assign U544 = ~(U419 & TX_CONTA_REG_4__SCAN_IN); 
assign U546 = ~(U419 & TX_CONTA_REG_3__SCAN_IN); 
assign U548 = ~(U419 & TX_CONTA_REG_2__SCAN_IN); 
assign U550 = ~(U377 & OUT_REG_REG_2__SCAN_IN); 
assign U556 = ~(U377 & OUT_REG_REG_3__SCAN_IN); 
assign U560 = ~(U438 & CONFIRM_REG_SCAN_IN); 
assign U562 = ~(U431 & U429); 
assign U567 = ~(U426 & ERROR_REG_SCAN_IN); 
assign U570 = ~(U508 & SEND_REG_SCAN_IN); 
assign U572 = ~(U425 & ITFC_STATE_REG_1__SCAN_IN); 
assign U573 = ~(U523 & ITFC_STATE_REG_0__SCAN_IN); 
assign U595 = ~(U424 & U422); 
assign U601 = ~(U436 & S2_REG_0__SCAN_IN); 
assign U602 = ~(U427 & S1_REG_2__SCAN_IN); 
assign U604 = ~(EOC & U428 & S1_REG_2__SCAN_IN); 
assign U605 = ~(U429 & U430 & S1_REG_1__SCAN_IN); 
assign ADD_291_U32 = ~ADD_291_U7; 
assign ADD_291_U54 = ~(ADD_291_U7 & TX_CONTA_REG_2__SCAN_IN); 
assign ADD_291_U56 = ~(ADD_291_U5 & TX_CONTA_REG_1__SCAN_IN); 
assign ADD_291_U57 = ~(ADD_291_U6 & TX_CONTA_REG_0__SCAN_IN); 
assign GT_255_U7 = GT_255_U9 & TX_CONTA_REG_3__SCAN_IN; 
assign U382 = ~(U439 & U472); 
assign U383 = ~(U434 & U561); 
assign U384 = ~(U605 & U604 & S1_REG_0__SCAN_IN); 
assign U388 = ~(U502 & U501); 
assign U394 = ~(U488 & U487); 
assign U409 = ~(U526 & U525); 
assign U452 = ~(U573 & U572); 
assign U471 = ~U448; 
assign U482 = ~(U480 & LOAD_REG_SCAN_IN); 
assign U484 = ~(U483 & S1_REG_0__SCAN_IN); 
assign U491 = ~(U489 & MUX_EN_REG_SCAN_IN); 
assign U492 = ~U434; 
assign U496 = ~(U495 & SEND_REG_SCAN_IN); 
assign U498 = ~U439; 
assign U499 = ~(U439 & MPX_REG_SCAN_IN); 
assign U504 = ~(U503 & SHOT_REG_SCAN_IN); 
assign U527 = ~U465; 
assign U532 = ~(U447 & U531); 
assign U549 = ~(U378 & OUT_REG_REG_6__SCAN_IN); 
assign U551 = ~(U473 & U445); 
assign U555 = ~(U378 & OUT_REG_REG_7__SCAN_IN); 
assign U564 = ~(U563 & U562); 
assign U566 = ~(U434 & SOC_REG_SCAN_IN); 
assign U569 = ~(U568 & U567); 
assign U574 = ~(U465 & OUT_REG_REG_7__SCAN_IN); 
assign U576 = ~(U465 & OUT_REG_REG_6__SCAN_IN); 
assign U578 = ~(U465 & OUT_REG_REG_5__SCAN_IN); 
assign U580 = ~(U465 & OUT_REG_REG_4__SCAN_IN); 
assign U582 = ~(U465 & OUT_REG_REG_3__SCAN_IN); 
assign U584 = ~(U465 & OUT_REG_REG_2__SCAN_IN); 
assign U586 = ~(U465 & OUT_REG_REG_1__SCAN_IN); 
assign U588 = ~(U465 & OUT_REG_REG_0__SCAN_IN); 
assign U594 = ~(U448 & NEXT_BIT_REG_0__SCAN_IN); 
assign U600 = ~(U560 & U441 & S2_REG_1__SCAN_IN); 
assign ADD_291_U9 = ~(ADD_291_U32 & TX_CONTA_REG_2__SCAN_IN); 
assign ADD_291_U29 = ~(ADD_291_U57 & ADD_291_U56); 
assign ADD_291_U55 = ~(ADD_291_U32 & ADD_291_U8); 
assign GT_255_U10 = GT_255_U7 | TX_CONTA_REG_4__SCAN_IN; 
assign U387 = ~(U505 & U504); 
assign U390 = ~(U497 & U496); 
assign U393 = ~(U491 & U490); 
assign U396 = ~(U482 & U481); 
assign U443 = ~(U492 & S1_REG_2__SCAN_IN); 
assign U463 = ~(U601 & U600); 
assign U466 = ~(U498 & U438); 
assign U486 = ~(U484 & SEND_DATA_REG_SCAN_IN); 
assign U506 = ~(U498 & MPX_REG_SCAN_IN); 
assign U552 = ~(U471 & OUT_REG_REG_4__SCAN_IN); 
assign U557 = ~(U471 & OUT_REG_REG_5__SCAN_IN); 
assign U565 = ~(U492 & U429); 
assign U571 = ~(U569 & U432); 
assign U575 = ~(DATA_IN_7_ & U527); 
assign U577 = ~(DATA_IN_6_ & U527); 
assign U579 = ~(DATA_IN_5_ & U527); 
assign U581 = ~(DATA_IN_4_ & U527); 
assign U583 = ~(DATA_IN_3_ & U527); 
assign U585 = ~(DATA_IN_2_ & U527); 
assign U587 = ~(DATA_IN_1_ & U527); 
assign U589 = ~(DATA_IN_0_ & U527); 
assign U603 = ~(U564 & S1_REG_0__SCAN_IN); 
assign ADD_291_U28 = ~(ADD_291_U55 & ADD_291_U54); 
assign ADD_291_U33 = ~ADD_291_U9; 
assign ADD_291_U52 = ~(ADD_291_U9 & TX_CONTA_REG_3__SCAN_IN); 
assign GT_255_U8 = GT_255_U10 & TX_CONTA_REG_6__SCAN_IN & TX_CONTA_REG_5__SCAN_IN; 
assign U389 = ~(U466 & U499); 
assign U395 = ~(U486 & U485); 
assign U450 = ~(U566 & U565); 
assign U451 = ~(U571 & U570); 
assign U453 = ~(U575 & U574); 
assign U454 = ~(U577 & U576); 
assign U455 = ~(U579 & U578); 
assign U456 = ~(U581 & U580); 
assign U457 = ~(U583 & U582); 
assign U458 = ~(U585 & U584); 
assign U459 = ~(U587 & U586); 
assign U460 = ~(U589 & U588); 
assign U464 = ~(U603 & U602); 
assign U467 = ~U466; 
assign U493 = ~U443; 
assign U494 = ~(U443 & LOAD_DATO_REG_SCAN_IN); 
assign U507 = ~(U506 & RDY_REG_SCAN_IN); 
assign U511 = ~(U443 & CANALE_REG_3__SCAN_IN); 
assign U513 = ~(U443 & CANALE_REG_2__SCAN_IN); 
assign U515 = ~(U443 & CANALE_REG_1__SCAN_IN); 
assign U516 = ~(U443 & CANALE_REG_0__SCAN_IN); 
assign U522 = ~(U443 & CONTA_TMP_REG_0__SCAN_IN); 
assign U554 = ~(U550 & U549 & U551 & U553 & U552); 
assign U559 = ~(U558 & U557 & U556 & U555); 
assign ADD_291_U11 = ~(ADD_291_U33 & TX_CONTA_REG_3__SCAN_IN); 
assign ADD_291_U53 = ~(ADD_291_U33 & ADD_291_U10); 
assign GT_255_U6 = GT_255_U8 | TX_CONTA_REG_9__SCAN_IN | TX_CONTA_REG_8__SCAN_IN | TX_CONTA_REG_7__SCAN_IN; 
assign U376 = U493 & U509; 
assign U385 = ~(U472 & U507); 
assign U386 = U467 | ADD_MPX2_REG_SCAN_IN; 
assign U391 = ~(U489 & U494); 
assign U420 = ~GT_255_U6; 
assign U421 = ~(GT_255_U6 & SEND_EN_REG_SCAN_IN); 
assign U517 = ~(U379 & U493 & CONTA_TMP_REG_2__SCAN_IN); 
assign U518 = ~(U493 & U379); 
assign U520 = ~(U493 & CONTA_TMP_REG_0__SCAN_IN); 
assign U598 = ~(U554 & NEXT_BIT_REG_0__SCAN_IN); 
assign U599 = ~(U559 & U422); 
assign ADD_291_U27 = ~(ADD_291_U53 & ADD_291_U52); 
assign ADD_291_U34 = ~ADD_291_U11; 
assign ADD_291_U50 = ~(ADD_291_U11 & TX_CONTA_REG_4__SCAN_IN); 
assign U375 = U420 & SEND_EN_REG_SCAN_IN; 
assign U417 = U517 & CONTA_TMP_REG_3__SCAN_IN; 
assign U444 = ~(U376 & U418); 
assign U468 = ~(U442 & U376 & CONTA_TMP_REG_0__SCAN_IN); 
assign U469 = ~(U376 & U379); 
assign U474 = ~U421; 
assign U510 = ~(U376 & CONTA_TMP_REG_3__SCAN_IN); 
assign U512 = ~(U376 & CONTA_TMP_REG_2__SCAN_IN); 
assign U519 = ~(U518 & CONTA_TMP_REG_2__SCAN_IN); 
assign U521 = ~(U520 & CONTA_TMP_REG_1__SCAN_IN); 
assign U596 = ~(U421 & NEXT_BIT_REG_0__SCAN_IN); 
assign ADD_291_U13 = ~(ADD_291_U34 & TX_CONTA_REG_4__SCAN_IN); 
assign ADD_291_U51 = ~(ADD_291_U34 & ADD_291_U12); 
assign U380 = ~(U599 & U598 & U474); 
assign U410 = ~(U444 & U522); 
assign U411 = ~(U468 & U521); 
assign U412 = ~(U469 & U519); 
assign U413 = ~(U444 & U516); 
assign U415 = ~(U512 & U469 & U513); 
assign U416 = ~(U511 & U510); 
assign U423 = ~(U474 & NEXT_BIT_REG_0__SCAN_IN); 
assign U470 = ~U444; 
assign U476 = ~(ADD_291_U29 & U375); 
assign U478 = ~(ADD_291_U5 & U375); 
assign U528 = ~(U595 & U594 & U474); 
assign U545 = ~(ADD_291_U27 & U375); 
assign U547 = ~(ADD_291_U28 & U375); 
assign U597 = ~(U474 & U532); 
assign ADD_291_U26 = ~(ADD_291_U51 & ADD_291_U50); 
assign ADD_291_U35 = ~ADD_291_U13; 
assign ADD_291_U48 = ~(ADD_291_U13 & TX_CONTA_REG_5__SCAN_IN); 
assign U397 = ~(U479 & U478); 
assign U398 = ~(U477 & U476); 
assign U399 = ~(U548 & U547); 
assign U400 = ~(U546 & U545); 
assign U462 = ~(U597 & U596); 
assign U475 = ~U423; 
assign U514 = ~(U470 & CONTA_TMP_REG_1__SCAN_IN); 
assign U529 = ~(U423 & NEXT_BIT_REG_1__SCAN_IN); 
assign U543 = ~(ADD_291_U26 & U375); 
assign U590 = ~(U423 & NEXT_BIT_REG_3__SCAN_IN); 
assign U592 = ~(U423 & NEXT_BIT_REG_2__SCAN_IN); 
assign ADD_291_U15 = ~(ADD_291_U35 & TX_CONTA_REG_5__SCAN_IN); 
assign ADD_291_U49 = ~(ADD_291_U35 & ADD_291_U14); 
assign U381 = U473 & U445 & U475; 
assign U401 = ~(U544 & U543); 
assign U407 = ~(U529 & U528); 
assign U414 = ~(U515 & U468 & U514); 
assign U591 = ~(U377 & U475); 
assign U593 = ~(U378 & U475); 
assign ADD_291_U25 = ~(ADD_291_U49 & ADD_291_U48); 
assign ADD_291_U36 = ~ADD_291_U15; 
assign ADD_291_U46 = ~(ADD_291_U15 & TX_CONTA_REG_6__SCAN_IN); 
assign U408 = ~(U593 & U592 & U448); 
assign U461 = ~(U591 & U590); 
assign U541 = ~(ADD_291_U25 & U375); 
assign ADD_291_U17 = ~(ADD_291_U36 & TX_CONTA_REG_6__SCAN_IN); 
assign ADD_291_U47 = ~(ADD_291_U36 & ADD_291_U16); 
assign U402 = ~(U542 & U541); 
assign ADD_291_U24 = ~(ADD_291_U47 & ADD_291_U46); 
assign ADD_291_U37 = ~ADD_291_U17; 
assign ADD_291_U44 = ~(ADD_291_U17 & TX_CONTA_REG_7__SCAN_IN); 
assign U539 = ~(ADD_291_U24 & U375); 
assign ADD_291_U19 = ~(ADD_291_U37 & TX_CONTA_REG_7__SCAN_IN); 
assign ADD_291_U45 = ~(ADD_291_U37 & ADD_291_U18); 
assign U403 = ~(U540 & U539); 
assign ADD_291_U23 = ~(ADD_291_U45 & ADD_291_U44); 
assign ADD_291_U38 = ~ADD_291_U19; 
assign ADD_291_U42 = ~(ADD_291_U19 & TX_CONTA_REG_8__SCAN_IN); 
assign U537 = ~(ADD_291_U23 & U375); 
assign ADD_291_U31 = ~(ADD_291_U38 & TX_CONTA_REG_8__SCAN_IN); 
assign ADD_291_U43 = ~(ADD_291_U38 & ADD_291_U20); 
assign U404 = ~(U538 & U537); 
assign ADD_291_U22 = ~(ADD_291_U43 & ADD_291_U42); 
assign ADD_291_U39 = ~ADD_291_U31; 
assign ADD_291_U40 = ~(ADD_291_U31 & TX_CONTA_REG_9__SCAN_IN); 
assign U535 = ~(ADD_291_U22 & U375); 
assign ADD_291_U41 = ~(ADD_291_U39 & ADD_291_U30); 
assign U405 = ~(U536 & U535); 
assign ADD_291_U21 = ~(ADD_291_U41 & ADD_291_U40); 
assign U533 = ~(ADD_291_U21 & U375); 
assign U406 = ~(U534 & U533); 
endmodule 
