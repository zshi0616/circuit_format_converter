module b17_C( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U212, U213, U216, U217, U218, U219, U220, U221, U222, U223, U224, U225, U226, U227, U228, U229, U230, U231, U232, U233, U234, U235, U236, U237, U238, U239, U240, U241, U242, U243, U244, U245, U246, U247, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, U280, U281, U282, U347, U348, U349, U350, U351, U352, U353, U354, U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U365, U366, U367, U368, U369, U370, U371, U372, U373, U374, U375, U376, P3_U2633, P3_U2634, P3_U2635, P3_U2636, P3_U2637, P3_U2638, P3_U2639, P3_U2640, P3_U2641, P3_U2642, P3_U2643, P3_U2644, P3_U2645, P3_U2646, P3_U2647, P3_U2648, P3_U2649, P3_U2650, P3_U2651, P3_U2652, P3_U2653, P3_U2654, P3_U2655, P3_U2656, P3_U2657, P3_U2658, P3_U2659, P3_U2660, P3_U2661, P3_U2662, P3_U2663, P3_U2664, P3_U2665, P3_U2666, P3_U2667, P3_U2668, P3_U2669, P3_U2670, P3_U2671, P3_U2672, P3_U2673, P3_U2674, P3_U2675, P3_U2676, P3_U2677, P3_U2678, P3_U2679, P3_U2680, P3_U2681, P3_U2682, P3_U2683, P3_U2684, P3_U2685, P3_U2686, P3_U2687, P3_U2688, P3_U2689, P3_U2690, P3_U2691, P3_U2692, P3_U2693, P3_U2694, P3_U2695, P3_U2696, P3_U2697, P3_U2698, P3_U2699, P3_U2700, P3_U2701, P3_U2702, P3_U2703, P3_U2704, P3_U2705, P3_U2706, P3_U2707, P3_U2708, P3_U2709, P3_U2710, P3_U2711, P3_U2712, P3_U2713, P3_U2714, P3_U2715, P3_U2716, P3_U2717, P3_U2718, P3_U2719, P3_U2720, P3_U2721, P3_U2722, P3_U2723, P3_U2724, P3_U2725, P3_U2726, P3_U2727, P3_U2728, P3_U2729, P3_U2730, P3_U2731, P3_U2732, P3_U2733, P3_U2734, P3_U2735, P3_U2736, P3_U2737, P3_U2738, P3_U2739, P3_U2740, P3_U2741, P3_U2742, P3_U2743, P3_U2744, P3_U2745, P3_U2746, P3_U2747, P3_U2748, P3_U2749, P3_U2750, P3_U2751, P3_U2752, P3_U2753, P3_U2754, P3_U2755, P3_U2756, P3_U2757, P3_U2758, P3_U2759, P3_U2760, P3_U2761, P3_U2762, P3_U2763, P3_U2764, P3_U2765, P3_U2766, P3_U2767, P3_U2768, P3_U2769, P3_U2770, P3_U2771, P3_U2772, P3_U2773, P3_U2774, P3_U2775, P3_U2776, P3_U2777, P3_U2778, P3_U2779, P3_U2780, P3_U2781, P3_U2782, P3_U2783, P3_U2784, P3_U2785, P3_U2786, P3_U2787, P3_U2788, P3_U2789, P3_U2790, P3_U2791, P3_U2792, P3_U2793, P3_U2794, P3_U2795, P3_U2796, P3_U2797, P3_U2798, P3_U2799, P3_U2800, P3_U2801, P3_U2802, P3_U2803, P3_U2804, P3_U2805, P3_U2806, P3_U2807, P3_U2808, P3_U2809, P3_U2810, P3_U2811, P3_U2812, P3_U2813, P3_U2814, P3_U2815, P3_U2816, P3_U2817, P3_U2818, P3_U2819, P3_U2820, P3_U2821, P3_U2822, P3_U2823, P3_U2824, P3_U2825, P3_U2826, P3_U2827, P3_U2828, P3_U2829, P3_U2830, P3_U2831, P3_U2832, P3_U2833, P3_U2834, P3_U2835, P3_U2836, P3_U2837, P3_U2838, P3_U2839, P3_U2840, P3_U2841, P3_U2842, P3_U2843, P3_U2844, P3_U2845, P3_U2846, P3_U2847, P3_U2848, P3_U2849, P3_U2850, P3_U2851, P3_U2852, P3_U2853, P3_U2854, P3_U2855, P3_U2856, P3_U2857, P3_U2858, P3_U2859, P3_U2860, P3_U2861, P3_U2862, P3_U2863, P3_U2864, P3_U2865, P3_U2866, P3_U2867, P3_U2868, P3_U2869, P3_U2870, P3_U2871, P3_U2872, P3_U2873, P3_U2874, P3_U2875, P3_U2876, P3_U2877, P3_U2878, P3_U2879, P3_U2880, P3_U2881, P3_U2882, P3_U2883, P3_U2884, P3_U2885, P3_U2886, P3_U2887, P3_U2888, P3_U2889, P3_U2890, P3_U2891, P3_U2892, P3_U2893, P3_U2894, P3_U2895, P3_U2896, P3_U2897, P3_U2898, P3_U2899, P3_U2900, P3_U2901, P3_U2902, P3_U2903, P3_U2904, P3_U2905, P3_U2906, P3_U2907, P3_U2908, P3_U2909, P3_U2910, P3_U2911, P3_U2912, P3_U2913, P3_U2914, P3_U2915, P3_U2916, P3_U2917, P3_U2918, P3_U2919, P3_U2920, P3_U2921, P3_U2922, P3_U2923, P3_U2924, P3_U2925, P3_U2926, P3_U2927, P3_U2928, P3_U2929, P3_U2930, P3_U2931, P3_U2932, P3_U2933, P3_U2934, P3_U2935, P3_U2936, P3_U2937, P3_U2938, P3_U2939, P3_U2940, P3_U2941, P3_U2942, P3_U2943, P3_U2944, P3_U2945, P3_U2946, P3_U2947, P3_U2948, P3_U2949, P3_U2950, P3_U2951, P3_U2952, P3_U2953, P3_U2954, P3_U2955, P3_U2956, P3_U2957, P3_U2958, P3_U2959, P3_U2960, P3_U2961, P3_U2962, P3_U2963, P3_U2964, P3_U2965, P3_U2966, P3_U2967, P3_U2968, P3_U2969, P3_U2970, P3_U2971, P3_U2972, P3_U2973, P3_U2974, P3_U2975, P3_U2976, P3_U2977, P3_U2978, P3_U2979, P3_U2980, P3_U2981, P3_U2982, P3_U2983, P3_U2984, P3_U2985, P3_U2986, P3_U2987, P3_U2988, P3_U2989, P3_U2990, P3_U2991, P3_U2992, P3_U2993, P3_U2994, P3_U2995, P3_U2996, P3_U2997, P3_U2998, P3_U2999, P3_U3000, P3_U3001, P3_U3002, P3_U3003, P3_U3004, P3_U3005, P3_U3006, P3_U3007, P3_U3008, P3_U3009, P3_U3010, P3_U3011, P3_U3012, P3_U3013, P3_U3014, P3_U3015, P3_U3016, P3_U3017, P3_U3018, P3_U3019, P3_U3020, P3_U3021, P3_U3022, P3_U3023, P3_U3024, P3_U3025, P3_U3026, P3_U3027, P3_U3028, P3_U3029, P3_U3030, P3_U3031, P3_U3032, P3_U3033, P3_U3034, P3_U3035, P3_U3036, P3_U3037, P3_U3038, P3_U3039, P3_U3040, P3_U3041, P3_U3042, P3_U3043, P3_U3044, P3_U3045, P3_U3046, P3_U3047, P3_U3048, P3_U3049, P3_U3050, P3_U3051, P3_U3052, P3_U3053, P3_U3054, P3_U3055, P3_U3056, P3_U3057, P3_U3058, P3_U3059, P3_U3060, P3_U3061, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3280, P3_U3281, P3_U3282, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U3292, P3_U3293, P3_U3294, P3_U3295, P3_U3296, P3_U3297, P3_U3298, P3_U3299, P2_U2814, P2_U2815, P2_U2816, P2_U2817, P2_U2818, P2_U2819, P2_U2820, P2_U2821, P2_U2822, P2_U2823, P2_U2824, P2_U2825, P2_U2826, P2_U2827, P2_U2828, P2_U2829, P2_U2830, P2_U2831, P2_U2832, P2_U2833, P2_U2834, P2_U2835, P2_U2836, P2_U2837, P2_U2838, P2_U2839, P2_U2840, P2_U2841, P2_U2842, P2_U2843, P2_U2844, P2_U2845, P2_U2846, P2_U2847, P2_U2848, P2_U2849, P2_U2850, P2_U2851, P2_U2852, P2_U2853, P2_U2854, P2_U2855, P2_U2856, P2_U2857, P2_U2858, P2_U2859, P2_U2860, P2_U2861, P2_U2862, P2_U2863, P2_U2864, P2_U2865, P2_U2866, P2_U2867, P2_U2868, P2_U2869, P2_U2870, P2_U2871, P2_U2872, P2_U2873, P2_U2874, P2_U2875, P2_U2876, P2_U2877, P2_U2878, P2_U2879, P2_U2880, P2_U2881, P2_U2882, P2_U2883, P2_U2884, P2_U2885, P2_U2886, P2_U2887, P2_U2888, P2_U2889, P2_U2890, P2_U2891, P2_U2892, P2_U2893, P2_U2894, P2_U2895, P2_U2896, P2_U2897, P2_U2898, P2_U2899, P2_U2900, P2_U2901, P2_U2902, P2_U2903, P2_U2904, P2_U2905, P2_U2906, P2_U2907, P2_U2908, P2_U2909, P2_U2910, P2_U2911, P2_U2912, P2_U2913, P2_U2914, P2_U2915, P2_U2916, P2_U2917, P2_U2918, P2_U2919, P2_U2920, P2_U2921, P2_U2922, P2_U2923, P2_U2924, P2_U2925, P2_U2926, P2_U2927, P2_U2928, P2_U2929, P2_U2930, P2_U2931, P2_U2932, P2_U2933, P2_U2934, P2_U2935, P2_U2936, P2_U2937, P2_U2938, P2_U2939, P2_U2940, P2_U2941, P2_U2942, P2_U2943, P2_U2944, P2_U2945, P2_U2946, P2_U2947, P2_U2948, P2_U2949, P2_U2950, P2_U2951, P2_U2952, P2_U2953, P2_U2954, P2_U2955, P2_U2956, P2_U2957, P2_U2958, P2_U2959, P2_U2960, P2_U2961, P2_U2962, P2_U2963, P2_U2964, P2_U2965, P2_U2966, P2_U2967, P2_U2968, P2_U2969, P2_U2970, P2_U2971, P2_U2972, P2_U2973, P2_U2974, P2_U2975, P2_U2976, P2_U2977, P2_U2978, P2_U2979, P2_U2980, P2_U2981, P2_U2982, P2_U2983, P2_U2984, P2_U2985, P2_U2986, P2_U2987, P2_U2988, P2_U2989, P2_U2990, P2_U2991, P2_U2992, P2_U2993, P2_U2994, P2_U2995, P2_U2996, P2_U2997, P2_U2998, P2_U2999, P2_U3000, P2_U3001, P2_U3002, P2_U3003, P2_U3004, P2_U3005, P2_U3006, P2_U3007, P2_U3008, P2_U3009, P2_U3010, P2_U3011, P2_U3012, P2_U3013, P2_U3014, P2_U3015, P2_U3016, P2_U3017, P2_U3018, P2_U3019, P2_U3020, P2_U3021, P2_U3022, P2_U3023, P2_U3024, P2_U3025, P2_U3026, P2_U3027, P2_U3028, P2_U3029, P2_U3030, P2_U3031, P2_U3032, P2_U3033, P2_U3034, P2_U3035, P2_U3036, P2_U3037, P2_U3038, P2_U3039, P2_U3040, P2_U3041, P2_U3042, P2_U3043, P2_U3044, P2_U3045, P2_U3046, P2_U3047, P2_U3048, P2_U3049, P2_U3050, P2_U3051, P2_U3052, P2_U3053, P2_U3054, P2_U3055, P2_U3056, P2_U3057, P2_U3058, P2_U3059, P2_U3060, P2_U3061, P2_U3062, P2_U3063, P2_U3064, P2_U3065, P2_U3066, P2_U3067, P2_U3068, P2_U3069, P2_U3070, P2_U3071, P2_U3072, P2_U3073, P2_U3074, P2_U3075, P2_U3076, P2_U3077, P2_U3078, P2_U3079, P2_U3080, P2_U3081, P2_U3082, P2_U3083, P2_U3084, P2_U3085, P2_U3086, P2_U3087, P2_U3088, P2_U3089, P2_U3090, P2_U3091, P2_U3092, P2_U3093, P2_U3094, P2_U3095, P2_U3096, P2_U3097, P2_U3098, P2_U3099, P2_U3100, P2_U3101, P2_U3102, P2_U3103, P2_U3104, P2_U3105, P2_U3106, P2_U3107, P2_U3108, P2_U3109, P2_U3110, P2_U3111, P2_U3112, P2_U3113, P2_U3114, P2_U3115, P2_U3116, P2_U3117, P2_U3118, P2_U3119, P2_U3120, P2_U3121, P2_U3122, P2_U3123, P2_U3124, P2_U3125, P2_U3126, P2_U3127, P2_U3128, P2_U3129, P2_U3130, P2_U3131, P2_U3132, P2_U3133, P2_U3134, P2_U3135, P2_U3136, P2_U3137, P2_U3138, P2_U3139, P2_U3140, P2_U3141, P2_U3142, P2_U3143, P2_U3144, P2_U3145, P2_U3146, P2_U3147, P2_U3148, P2_U3149, P2_U3150, P2_U3151, P2_U3152, P2_U3153, P2_U3154, P2_U3155, P2_U3156, P2_U3157, P2_U3158, P2_U3159, P2_U3160, P2_U3161, P2_U3162, P2_U3163, P2_U3164, P2_U3165, P2_U3166, P2_U3167, P2_U3168, P2_U3169, P2_U3170, P2_U3171, P2_U3172, P2_U3173, P2_U3174, P2_U3175, P2_U3176, P2_U3177, P2_U3178, P2_U3179, P2_U3180, P2_U3181, P2_U3182, P2_U3183, P2_U3184, P2_U3185, P2_U3186, P2_U3187, P2_U3188, P2_U3189, P2_U3190, P2_U3191, P2_U3192, P2_U3193, P2_U3194, P2_U3195, P2_U3196, P2_U3197, P2_U3198, P2_U3199, P2_U3200, P2_U3201, P2_U3202, P2_U3203, P2_U3204, P2_U3205, P2_U3206, P2_U3207, P2_U3208, P2_U3209, P2_U3210, P2_U3211, P2_U3212, P2_U3213, P2_U3214, P2_U3215, P2_U3216, P2_U3217, P2_U3218, P2_U3219, P2_U3220, P2_U3221, P2_U3222, P2_U3223, P2_U3224, P2_U3225, P2_U3226, P2_U3227, P2_U3228, P2_U3229, P2_U3230, P2_U3231, P2_U3232, P2_U3233, P2_U3234, P2_U3235, P2_U3236, P2_U3237, P2_U3238, P2_U3239, P2_U3240, P2_U3241, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3591, P2_U3592, P2_U3593, P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3608, P2_U3609, P2_U3610, P2_U3611, P2_U3612, P1_U2801, P1_U2802, P1_U2803, P1_U2804, P1_U2805, P1_U2806, P1_U2807, P1_U2808, P1_U2809, P1_U2810, P1_U2811, P1_U2812, P1_U2813, P1_U2814, P1_U2815, P1_U2816, P1_U2817, P1_U2818, P1_U2819, P1_U2820, P1_U2821, P1_U2822, P1_U2823, P1_U2824, P1_U2825, P1_U2826, P1_U2827, P1_U2828, P1_U2829, P1_U2830, P1_U2831, P1_U2832, P1_U2833, P1_U2834, P1_U2835, P1_U2836, P1_U2837, P1_U2838, P1_U2839, P1_U2840, P1_U2841, P1_U2842, P1_U2843, P1_U2844, P1_U2845, P1_U2846, P1_U2847, P1_U2848, P1_U2849, P1_U2850, P1_U2851, P1_U2852, P1_U2853, P1_U2854, P1_U2855, P1_U2856, P1_U2857, P1_U2858, P1_U2859, P1_U2860, P1_U2861, P1_U2862, P1_U2863, P1_U2864, P1_U2865, P1_U2866, P1_U2867, P1_U2868, P1_U2869, P1_U2870, P1_U2871, P1_U2872, P1_U2873, P1_U2874, P1_U2875, P1_U2876, P1_U2877, P1_U2878, P1_U2879, P1_U2880, P1_U2881, P1_U2882, P1_U2883, P1_U2884, P1_U2885, P1_U2886, P1_U2887, P1_U2888, P1_U2889, P1_U2890, P1_U2891, P1_U2892, P1_U2893, P1_U2894, P1_U2895, P1_U2896, P1_U2897, P1_U2898, P1_U2899, P1_U2900, P1_U2901, P1_U2902, P1_U2903, P1_U2904, P1_U2905, P1_U2906, P1_U2907, P1_U2908, P1_U2909, P1_U2910, P1_U2911, P1_U2912, P1_U2913, P1_U2914, P1_U2915, P1_U2916, P1_U2917, P1_U2918, P1_U2919, P1_U2920, P1_U2921, P1_U2922, P1_U2923, P1_U2924, P1_U2925, P1_U2926, P1_U2927, P1_U2928, P1_U2929, P1_U2930, P1_U2931, P1_U2932, P1_U2933, P1_U2934, P1_U2935, P1_U2936, P1_U2937, P1_U2938, P1_U2939, P1_U2940, P1_U2941, P1_U2942, P1_U2943, P1_U2944, P1_U2945, P1_U2946, P1_U2947, P1_U2948, P1_U2949, P1_U2950, P1_U2951, P1_U2952, P1_U2953, P1_U2954, P1_U2955, P1_U2956, P1_U2957, P1_U2958, P1_U2959, P1_U2960, P1_U2961, P1_U2962, P1_U2963, P1_U2964, P1_U2965, P1_U2966, P1_U2967, P1_U2968, P1_U2969, P1_U2970, P1_U2971, P1_U2972, P1_U2973, P1_U2974, P1_U2975, P1_U2976, P1_U2977, P1_U2978, P1_U2979, P1_U2980, P1_U2981, P1_U2982, P1_U2983, P1_U2984, P1_U2985, P1_U2986, P1_U2987, P1_U2988, P1_U2989, P1_U2990, P1_U2991, P1_U2992, P1_U2993, P1_U2994, P1_U2995, P1_U2996, P1_U2997, P1_U2998, P1_U2999, P1_U3000, P1_U3001, P1_U3002, P1_U3003, P1_U3004, P1_U3005, P1_U3006, P1_U3007, P1_U3008, P1_U3009, P1_U3010, P1_U3011, P1_U3012, P1_U3013, P1_U3014, P1_U3015, P1_U3016, P1_U3017, P1_U3018, P1_U3019, P1_U3020, P1_U3021, P1_U3022, P1_U3023, P1_U3024, P1_U3025, P1_U3026, P1_U3027, P1_U3028, P1_U3029, P1_U3030, P1_U3031, P1_U3032, P1_U3033, P1_U3034, P1_U3035, P1_U3036, P1_U3037, P1_U3038, P1_U3039, P1_U3040, P1_U3041, P1_U3042, P1_U3043, P1_U3044, P1_U3045, P1_U3046, P1_U3047, P1_U3048, P1_U3049, P1_U3050, P1_U3051, P1_U3052, P1_U3053, P1_U3054, P1_U3055, P1_U3056, P1_U3057, P1_U3058, P1_U3059, P1_U3060, P1_U3061, P1_U3062, P1_U3063, P1_U3064, P1_U3065, P1_U3066, P1_U3067, P1_U3068, P1_U3069, P1_U3070, P1_U3071, P1_U3072, P1_U3073, P1_U3074, P1_U3075, P1_U3076, P1_U3077, P1_U3078, P1_U3079, P1_U3080, P1_U3081, P1_U3082, P1_U3083, P1_U3084, P1_U3085, P1_U3086, P1_U3087, P1_U3088, P1_U3089, P1_U3090, P1_U3091, P1_U3092, P1_U3093, P1_U3094, P1_U3095, P1_U3096, P1_U3097, P1_U3098, P1_U3099, P1_U3100, P1_U3101, P1_U3102, P1_U3103, P1_U3104, P1_U3105, P1_U3106, P1_U3107, P1_U3108, P1_U3109, P1_U3110, P1_U3111, P1_U3112, P1_U3113, P1_U3114, P1_U3115, P1_U3116, P1_U3117, P1_U3118, P1_U3119, P1_U3120, P1_U3121, P1_U3122, P1_U3123, P1_U3124, P1_U3125, P1_U3126, P1_U3127, P1_U3128, P1_U3129, P1_U3130, P1_U3131, P1_U3132, P1_U3133, P1_U3134, P1_U3135, P1_U3136, P1_U3137, P1_U3138, P1_U3139, P1_U3140, P1_U3141, P1_U3142, P1_U3143, P1_U3144, P1_U3145, P1_U3146, P1_U3147, P1_U3148, P1_U3149, P1_U3150, P1_U3151, P1_U3152, P1_U3153, P1_U3154, P1_U3155, P1_U3156, P1_U3157, P1_U3158, P1_U3159, P1_U3160, P1_U3161, P1_U3162, P1_U3163, P1_U3164, P1_U3165, P1_U3166, P1_U3167, P1_U3168, P1_U3169, P1_U3170, P1_U3171, P1_U3172, P1_U3173, P1_U3174, P1_U3175, P1_U3176, P1_U3177, P1_U3178, P1_U3179, P1_U3180, P1_U3181, P1_U3182, P1_U3183, P1_U3184, P1_U3185, P1_U3186, P1_U3187, P1_U3188, P1_U3189, P1_U3190, P1_U3191, P1_U3192, P1_U3193, P1_U3194, P1_U3195, P1_U3196, P1_U3197, P1_U3198, P1_U3199, P1_U3200, P1_U3201, P1_U3202, P1_U3203, P1_U3204, P1_U3205, P1_U3206, P1_U3207, P1_U3208, P1_U3209, P1_U3210, P1_U3211, P1_U3212, P1_U3213, P1_U3214, P1_U3215, P1_U3216, P1_U3217, P1_U3218, P1_U3219, P1_U3220, P1_U3221, P1_U3222, P1_U3223, P1_U3224, P1_U3225, P1_U3226, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3464, P1_U3465, P1_U3466, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3481, P1_U3482, P1_U3483, P1_U3484, P1_U3485, P1_U3486, P1_U3487); 
input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN; 
output U212, U213, U216, U217, U218, U219, U220, U221, U222, U223, U224, U225, U226, U227, U228, U229, U230, U231, U232, U233, U234, U235, U236, U237, U238, U239, U240, U241, U242, U243, U244, U245, U246, U247, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, U280, U281, U282, U347, U348, U349, U350, U351, U352, U353, U354, U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U365, U366, U367, U368, U369, U370, U371, U372, U373, U374, U375, U376, P3_U2633, P3_U2634, P3_U2635, P3_U2636, P3_U2637, P3_U2638, P3_U2639, P3_U2640, P3_U2641, P3_U2642, P3_U2643, P3_U2644, P3_U2645, P3_U2646, P3_U2647, P3_U2648, P3_U2649, P3_U2650, P3_U2651, P3_U2652, P3_U2653, P3_U2654, P3_U2655, P3_U2656, P3_U2657, P3_U2658, P3_U2659, P3_U2660, P3_U2661, P3_U2662, P3_U2663, P3_U2664, P3_U2665, P3_U2666, P3_U2667, P3_U2668, P3_U2669, P3_U2670, P3_U2671, P3_U2672, P3_U2673, P3_U2674, P3_U2675, P3_U2676, P3_U2677, P3_U2678, P3_U2679, P3_U2680, P3_U2681, P3_U2682, P3_U2683, P3_U2684, P3_U2685, P3_U2686, P3_U2687, P3_U2688, P3_U2689, P3_U2690, P3_U2691, P3_U2692, P3_U2693, P3_U2694, P3_U2695, P3_U2696, P3_U2697, P3_U2698, P3_U2699, P3_U2700, P3_U2701, P3_U2702, P3_U2703, P3_U2704, P3_U2705, P3_U2706, P3_U2707, P3_U2708, P3_U2709, P3_U2710, P3_U2711, P3_U2712, P3_U2713, P3_U2714, P3_U2715, P3_U2716, P3_U2717, P3_U2718, P3_U2719, P3_U2720, P3_U2721, P3_U2722, P3_U2723, P3_U2724, P3_U2725, P3_U2726, P3_U2727, P3_U2728, P3_U2729, P3_U2730, P3_U2731, P3_U2732, P3_U2733, P3_U2734, P3_U2735, P3_U2736, P3_U2737, P3_U2738, P3_U2739, P3_U2740, P3_U2741, P3_U2742, P3_U2743, P3_U2744, P3_U2745, P3_U2746, P3_U2747, P3_U2748, P3_U2749, P3_U2750, P3_U2751, P3_U2752, P3_U2753, P3_U2754, P3_U2755, P3_U2756, P3_U2757, P3_U2758, P3_U2759, P3_U2760, P3_U2761, P3_U2762, P3_U2763, P3_U2764, P3_U2765, P3_U2766, P3_U2767, P3_U2768, P3_U2769, P3_U2770, P3_U2771, P3_U2772, P3_U2773, P3_U2774, P3_U2775, P3_U2776, P3_U2777, P3_U2778, P3_U2779, P3_U2780, P3_U2781, P3_U2782, P3_U2783, P3_U2784, P3_U2785, P3_U2786, P3_U2787, P3_U2788, P3_U2789, P3_U2790, P3_U2791, P3_U2792, P3_U2793, P3_U2794, P3_U2795, P3_U2796, P3_U2797, P3_U2798, P3_U2799, P3_U2800, P3_U2801, P3_U2802, P3_U2803, P3_U2804, P3_U2805, P3_U2806, P3_U2807, P3_U2808, P3_U2809, P3_U2810, P3_U2811, P3_U2812, P3_U2813, P3_U2814, P3_U2815, P3_U2816, P3_U2817, P3_U2818, P3_U2819, P3_U2820, P3_U2821, P3_U2822, P3_U2823, P3_U2824, P3_U2825, P3_U2826, P3_U2827, P3_U2828, P3_U2829, P3_U2830, P3_U2831, P3_U2832, P3_U2833, P3_U2834, P3_U2835, P3_U2836, P3_U2837, P3_U2838, P3_U2839, P3_U2840, P3_U2841, P3_U2842, P3_U2843, P3_U2844, P3_U2845, P3_U2846, P3_U2847, P3_U2848, P3_U2849, P3_U2850, P3_U2851, P3_U2852, P3_U2853, P3_U2854, P3_U2855, P3_U2856, P3_U2857, P3_U2858, P3_U2859, P3_U2860, P3_U2861, P3_U2862, P3_U2863, P3_U2864, P3_U2865, P3_U2866, P3_U2867, P3_U2868, P3_U2869, P3_U2870, P3_U2871, P3_U2872, P3_U2873, P3_U2874, P3_U2875, P3_U2876, P3_U2877, P3_U2878, P3_U2879, P3_U2880, P3_U2881, P3_U2882, P3_U2883, P3_U2884, P3_U2885, P3_U2886, P3_U2887, P3_U2888, P3_U2889, P3_U2890, P3_U2891, P3_U2892, P3_U2893, P3_U2894, P3_U2895, P3_U2896, P3_U2897, P3_U2898, P3_U2899, P3_U2900, P3_U2901, P3_U2902, P3_U2903, P3_U2904, P3_U2905, P3_U2906, P3_U2907, P3_U2908, P3_U2909, P3_U2910, P3_U2911, P3_U2912, P3_U2913, P3_U2914, P3_U2915, P3_U2916, P3_U2917, P3_U2918, P3_U2919, P3_U2920, P3_U2921, P3_U2922, P3_U2923, P3_U2924, P3_U2925, P3_U2926, P3_U2927, P3_U2928, P3_U2929, P3_U2930, P3_U2931, P3_U2932, P3_U2933, P3_U2934, P3_U2935, P3_U2936, P3_U2937, P3_U2938, P3_U2939, P3_U2940, P3_U2941, P3_U2942, P3_U2943, P3_U2944, P3_U2945, P3_U2946, P3_U2947, P3_U2948, P3_U2949, P3_U2950, P3_U2951, P3_U2952, P3_U2953, P3_U2954, P3_U2955, P3_U2956, P3_U2957, P3_U2958, P3_U2959, P3_U2960, P3_U2961, P3_U2962, P3_U2963, P3_U2964, P3_U2965, P3_U2966, P3_U2967, P3_U2968, P3_U2969, P3_U2970, P3_U2971, P3_U2972, P3_U2973, P3_U2974, P3_U2975, P3_U2976, P3_U2977, P3_U2978, P3_U2979, P3_U2980, P3_U2981, P3_U2982, P3_U2983, P3_U2984, P3_U2985, P3_U2986, P3_U2987, P3_U2988, P3_U2989, P3_U2990, P3_U2991, P3_U2992, P3_U2993, P3_U2994, P3_U2995, P3_U2996, P3_U2997, P3_U2998, P3_U2999, P3_U3000, P3_U3001, P3_U3002, P3_U3003, P3_U3004, P3_U3005, P3_U3006, P3_U3007, P3_U3008, P3_U3009, P3_U3010, P3_U3011, P3_U3012, P3_U3013, P3_U3014, P3_U3015, P3_U3016, P3_U3017, P3_U3018, P3_U3019, P3_U3020, P3_U3021, P3_U3022, P3_U3023, P3_U3024, P3_U3025, P3_U3026, P3_U3027, P3_U3028, P3_U3029, P3_U3030, P3_U3031, P3_U3032, P3_U3033, P3_U3034, P3_U3035, P3_U3036, P3_U3037, P3_U3038, P3_U3039, P3_U3040, P3_U3041, P3_U3042, P3_U3043, P3_U3044, P3_U3045, P3_U3046, P3_U3047, P3_U3048, P3_U3049, P3_U3050, P3_U3051, P3_U3052, P3_U3053, P3_U3054, P3_U3055, P3_U3056, P3_U3057, P3_U3058, P3_U3059, P3_U3060, P3_U3061, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3280, P3_U3281, P3_U3282, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U3292, P3_U3293, P3_U3294, P3_U3295, P3_U3296, P3_U3297, P3_U3298, P3_U3299, P2_U2814, P2_U2815, P2_U2816, P2_U2817, P2_U2818, P2_U2819, P2_U2820, P2_U2821, P2_U2822, P2_U2823, P2_U2824, P2_U2825, P2_U2826, P2_U2827, P2_U2828, P2_U2829, P2_U2830, P2_U2831, P2_U2832, P2_U2833, P2_U2834, P2_U2835, P2_U2836, P2_U2837, P2_U2838, P2_U2839, P2_U2840, P2_U2841, P2_U2842, P2_U2843, P2_U2844, P2_U2845, P2_U2846, P2_U2847, P2_U2848, P2_U2849, P2_U2850, P2_U2851, P2_U2852, P2_U2853, P2_U2854, P2_U2855, P2_U2856, P2_U2857, P2_U2858, P2_U2859, P2_U2860, P2_U2861, P2_U2862, P2_U2863, P2_U2864, P2_U2865, P2_U2866, P2_U2867, P2_U2868, P2_U2869, P2_U2870, P2_U2871, P2_U2872, P2_U2873, P2_U2874, P2_U2875, P2_U2876, P2_U2877, P2_U2878, P2_U2879, P2_U2880, P2_U2881, P2_U2882, P2_U2883, P2_U2884, P2_U2885, P2_U2886, P2_U2887, P2_U2888, P2_U2889, P2_U2890, P2_U2891, P2_U2892, P2_U2893, P2_U2894, P2_U2895, P2_U2896, P2_U2897, P2_U2898, P2_U2899, P2_U2900, P2_U2901, P2_U2902, P2_U2903, P2_U2904, P2_U2905, P2_U2906, P2_U2907, P2_U2908, P2_U2909, P2_U2910, P2_U2911, P2_U2912, P2_U2913, P2_U2914, P2_U2915, P2_U2916, P2_U2917, P2_U2918, P2_U2919, P2_U2920, P2_U2921, P2_U2922, P2_U2923, P2_U2924, P2_U2925, P2_U2926, P2_U2927, P2_U2928, P2_U2929, P2_U2930, P2_U2931, P2_U2932, P2_U2933, P2_U2934, P2_U2935, P2_U2936, P2_U2937, P2_U2938, P2_U2939, P2_U2940, P2_U2941, P2_U2942, P2_U2943, P2_U2944, P2_U2945, P2_U2946, P2_U2947, P2_U2948, P2_U2949, P2_U2950, P2_U2951, P2_U2952, P2_U2953, P2_U2954, P2_U2955, P2_U2956, P2_U2957, P2_U2958, P2_U2959, P2_U2960, P2_U2961, P2_U2962, P2_U2963, P2_U2964, P2_U2965, P2_U2966, P2_U2967, P2_U2968, P2_U2969, P2_U2970, P2_U2971, P2_U2972, P2_U2973, P2_U2974, P2_U2975, P2_U2976, P2_U2977, P2_U2978, P2_U2979, P2_U2980, P2_U2981, P2_U2982, P2_U2983, P2_U2984, P2_U2985, P2_U2986, P2_U2987, P2_U2988, P2_U2989, P2_U2990, P2_U2991, P2_U2992, P2_U2993, P2_U2994, P2_U2995, P2_U2996, P2_U2997, P2_U2998, P2_U2999, P2_U3000, P2_U3001, P2_U3002, P2_U3003, P2_U3004, P2_U3005, P2_U3006, P2_U3007, P2_U3008, P2_U3009, P2_U3010, P2_U3011, P2_U3012, P2_U3013, P2_U3014, P2_U3015, P2_U3016, P2_U3017, P2_U3018, P2_U3019, P2_U3020, P2_U3021, P2_U3022, P2_U3023, P2_U3024, P2_U3025, P2_U3026, P2_U3027, P2_U3028, P2_U3029, P2_U3030, P2_U3031, P2_U3032, P2_U3033, P2_U3034, P2_U3035, P2_U3036, P2_U3037, P2_U3038, P2_U3039, P2_U3040, P2_U3041, P2_U3042, P2_U3043, P2_U3044, P2_U3045, P2_U3046, P2_U3047, P2_U3048, P2_U3049, P2_U3050, P2_U3051, P2_U3052, P2_U3053, P2_U3054, P2_U3055, P2_U3056, P2_U3057, P2_U3058, P2_U3059, P2_U3060, P2_U3061, P2_U3062, P2_U3063, P2_U3064, P2_U3065, P2_U3066, P2_U3067, P2_U3068, P2_U3069, P2_U3070, P2_U3071, P2_U3072, P2_U3073, P2_U3074, P2_U3075, P2_U3076, P2_U3077, P2_U3078, P2_U3079, P2_U3080, P2_U3081, P2_U3082, P2_U3083, P2_U3084, P2_U3085, P2_U3086, P2_U3087, P2_U3088, P2_U3089, P2_U3090, P2_U3091, P2_U3092, P2_U3093, P2_U3094, P2_U3095, P2_U3096, P2_U3097, P2_U3098, P2_U3099, P2_U3100, P2_U3101, P2_U3102, P2_U3103, P2_U3104, P2_U3105, P2_U3106, P2_U3107, P2_U3108, P2_U3109, P2_U3110, P2_U3111, P2_U3112, P2_U3113, P2_U3114, P2_U3115, P2_U3116, P2_U3117, P2_U3118, P2_U3119, P2_U3120, P2_U3121, P2_U3122, P2_U3123, P2_U3124, P2_U3125, P2_U3126, P2_U3127, P2_U3128, P2_U3129, P2_U3130, P2_U3131, P2_U3132, P2_U3133, P2_U3134, P2_U3135, P2_U3136, P2_U3137, P2_U3138, P2_U3139, P2_U3140, P2_U3141, P2_U3142, P2_U3143, P2_U3144, P2_U3145, P2_U3146, P2_U3147, P2_U3148, P2_U3149, P2_U3150, P2_U3151, P2_U3152, P2_U3153, P2_U3154, P2_U3155, P2_U3156, P2_U3157, P2_U3158, P2_U3159, P2_U3160, P2_U3161, P2_U3162, P2_U3163, P2_U3164, P2_U3165, P2_U3166, P2_U3167, P2_U3168, P2_U3169, P2_U3170, P2_U3171, P2_U3172, P2_U3173, P2_U3174, P2_U3175, P2_U3176, P2_U3177, P2_U3178, P2_U3179, P2_U3180, P2_U3181, P2_U3182, P2_U3183, P2_U3184, P2_U3185, P2_U3186, P2_U3187, P2_U3188, P2_U3189, P2_U3190, P2_U3191, P2_U3192, P2_U3193, P2_U3194, P2_U3195, P2_U3196, P2_U3197, P2_U3198, P2_U3199, P2_U3200, P2_U3201, P2_U3202, P2_U3203, P2_U3204, P2_U3205, P2_U3206, P2_U3207, P2_U3208, P2_U3209, P2_U3210, P2_U3211, P2_U3212, P2_U3213, P2_U3214, P2_U3215, P2_U3216, P2_U3217, P2_U3218, P2_U3219, P2_U3220, P2_U3221, P2_U3222, P2_U3223, P2_U3224, P2_U3225, P2_U3226, P2_U3227, P2_U3228, P2_U3229, P2_U3230, P2_U3231, P2_U3232, P2_U3233, P2_U3234, P2_U3235, P2_U3236, P2_U3237, P2_U3238, P2_U3239, P2_U3240, P2_U3241, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3591, P2_U3592, P2_U3593, P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3608, P2_U3609, P2_U3610, P2_U3611, P2_U3612, P1_U2801, P1_U2802, P1_U2803, P1_U2804, P1_U2805, P1_U2806, P1_U2807, P1_U2808, P1_U2809, P1_U2810, P1_U2811, P1_U2812, P1_U2813, P1_U2814, P1_U2815, P1_U2816, P1_U2817, P1_U2818, P1_U2819, P1_U2820, P1_U2821, P1_U2822, P1_U2823, P1_U2824, P1_U2825, P1_U2826, P1_U2827, P1_U2828, P1_U2829, P1_U2830, P1_U2831, P1_U2832, P1_U2833, P1_U2834, P1_U2835, P1_U2836, P1_U2837, P1_U2838, P1_U2839, P1_U2840, P1_U2841, P1_U2842, P1_U2843, P1_U2844, P1_U2845, P1_U2846, P1_U2847, P1_U2848, P1_U2849, P1_U2850, P1_U2851, P1_U2852, P1_U2853, P1_U2854, P1_U2855, P1_U2856, P1_U2857, P1_U2858, P1_U2859, P1_U2860, P1_U2861, P1_U2862, P1_U2863, P1_U2864, P1_U2865, P1_U2866, P1_U2867, P1_U2868, P1_U2869, P1_U2870, P1_U2871, P1_U2872, P1_U2873, P1_U2874, P1_U2875, P1_U2876, P1_U2877, P1_U2878, P1_U2879, P1_U2880, P1_U2881, P1_U2882, P1_U2883, P1_U2884, P1_U2885, P1_U2886, P1_U2887, P1_U2888, P1_U2889, P1_U2890, P1_U2891, P1_U2892, P1_U2893, P1_U2894, P1_U2895, P1_U2896, P1_U2897, P1_U2898, P1_U2899, P1_U2900, P1_U2901, P1_U2902, P1_U2903, P1_U2904, P1_U2905, P1_U2906, P1_U2907, P1_U2908, P1_U2909, P1_U2910, P1_U2911, P1_U2912, P1_U2913, P1_U2914, P1_U2915, P1_U2916, P1_U2917, P1_U2918, P1_U2919, P1_U2920, P1_U2921, P1_U2922, P1_U2923, P1_U2924, P1_U2925, P1_U2926, P1_U2927, P1_U2928, P1_U2929, P1_U2930, P1_U2931, P1_U2932, P1_U2933, P1_U2934, P1_U2935, P1_U2936, P1_U2937, P1_U2938, P1_U2939, P1_U2940, P1_U2941, P1_U2942, P1_U2943, P1_U2944, P1_U2945, P1_U2946, P1_U2947, P1_U2948, P1_U2949, P1_U2950, P1_U2951, P1_U2952, P1_U2953, P1_U2954, P1_U2955, P1_U2956, P1_U2957, P1_U2958, P1_U2959, P1_U2960, P1_U2961, P1_U2962, P1_U2963, P1_U2964, P1_U2965, P1_U2966, P1_U2967, P1_U2968, P1_U2969, P1_U2970, P1_U2971, P1_U2972, P1_U2973, P1_U2974, P1_U2975, P1_U2976, P1_U2977, P1_U2978, P1_U2979, P1_U2980, P1_U2981, P1_U2982, P1_U2983, P1_U2984, P1_U2985, P1_U2986, P1_U2987, P1_U2988, P1_U2989, P1_U2990, P1_U2991, P1_U2992, P1_U2993, P1_U2994, P1_U2995, P1_U2996, P1_U2997, P1_U2998, P1_U2999, P1_U3000, P1_U3001, P1_U3002, P1_U3003, P1_U3004, P1_U3005, P1_U3006, P1_U3007, P1_U3008, P1_U3009, P1_U3010, P1_U3011, P1_U3012, P1_U3013, P1_U3014, P1_U3015, P1_U3016, P1_U3017, P1_U3018, P1_U3019, P1_U3020, P1_U3021, P1_U3022, P1_U3023, P1_U3024, P1_U3025, P1_U3026, P1_U3027, P1_U3028, P1_U3029, P1_U3030, P1_U3031, P1_U3032, P1_U3033, P1_U3034, P1_U3035, P1_U3036, P1_U3037, P1_U3038, P1_U3039, P1_U3040, P1_U3041, P1_U3042, P1_U3043, P1_U3044, P1_U3045, P1_U3046, P1_U3047, P1_U3048, P1_U3049, P1_U3050, P1_U3051, P1_U3052, P1_U3053, P1_U3054, P1_U3055, P1_U3056, P1_U3057, P1_U3058, P1_U3059, P1_U3060, P1_U3061, P1_U3062, P1_U3063, P1_U3064, P1_U3065, P1_U3066, P1_U3067, P1_U3068, P1_U3069, P1_U3070, P1_U3071, P1_U3072, P1_U3073, P1_U3074, P1_U3075, P1_U3076, P1_U3077, P1_U3078, P1_U3079, P1_U3080, P1_U3081, P1_U3082, P1_U3083, P1_U3084, P1_U3085, P1_U3086, P1_U3087, P1_U3088, P1_U3089, P1_U3090, P1_U3091, P1_U3092, P1_U3093, P1_U3094, P1_U3095, P1_U3096, P1_U3097, P1_U3098, P1_U3099, P1_U3100, P1_U3101, P1_U3102, P1_U3103, P1_U3104, P1_U3105, P1_U3106, P1_U3107, P1_U3108, P1_U3109, P1_U3110, P1_U3111, P1_U3112, P1_U3113, P1_U3114, P1_U3115, P1_U3116, P1_U3117, P1_U3118, P1_U3119, P1_U3120, P1_U3121, P1_U3122, P1_U3123, P1_U3124, P1_U3125, P1_U3126, P1_U3127, P1_U3128, P1_U3129, P1_U3130, P1_U3131, P1_U3132, P1_U3133, P1_U3134, P1_U3135, P1_U3136, P1_U3137, P1_U3138, P1_U3139, P1_U3140, P1_U3141, P1_U3142, P1_U3143, P1_U3144, P1_U3145, P1_U3146, P1_U3147, P1_U3148, P1_U3149, P1_U3150, P1_U3151, P1_U3152, P1_U3153, P1_U3154, P1_U3155, P1_U3156, P1_U3157, P1_U3158, P1_U3159, P1_U3160, P1_U3161, P1_U3162, P1_U3163, P1_U3164, P1_U3165, P1_U3166, P1_U3167, P1_U3168, P1_U3169, P1_U3170, P1_U3171, P1_U3172, P1_U3173, P1_U3174, P1_U3175, P1_U3176, P1_U3177, P1_U3178, P1_U3179, P1_U3180, P1_U3181, P1_U3182, P1_U3183, P1_U3184, P1_U3185, P1_U3186, P1_U3187, P1_U3188, P1_U3189, P1_U3190, P1_U3191, P1_U3192, P1_U3193, P1_U3194, P1_U3195, P1_U3196, P1_U3197, P1_U3198, P1_U3199, P1_U3200, P1_U3201, P1_U3202, P1_U3203, P1_U3204, P1_U3205, P1_U3206, P1_U3207, P1_U3208, P1_U3209, P1_U3210, P1_U3211, P1_U3212, P1_U3213, P1_U3214, P1_U3215, P1_U3216, P1_U3217, P1_U3218, P1_U3219, P1_U3220, P1_U3221, P1_U3222, P1_U3223, P1_U3224, P1_U3225, P1_U3226, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3464, P1_U3465, P1_U3466, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3481, P1_U3482, P1_U3483, P1_U3484, P1_U3485, P1_U3486, P1_U3487; 
wire U207, U208, U209, U210, U211, U214, U215, U248, U249, U250, U283, U284, U285, U286, U287, U288, U289, U290, U291, U292, U293, U294, U295, U296, U297, U298, U299, U300, U301, U302, U303, U304, U305, U306, U307, U308, U309, U310, U311, U312, U313, U314, U315, U316, U317, U318, U319, U320, U321, U322, U323, U324, U325, U326, U327, U328, U329, U330, U331, U332, U333, U334, U335, U336, U337, U338, U339, U340, U341, U342, U343, U344, U345, U346, U377, U378, U379, U380, U381, U382, U383, U384, U385, U386, U387, U388, U389, U390, U391, U392, U393, U394, U395, U396, U397, U398, U399, U400, U401, U402, U403, U404, U405, U406, U407, U408, U409, U410, U411, U412, U413, U414, U415, U416, U417, U418, U419, U420, U421, U422, U423, U424, U425, U426, U427, U428, U429, U430, U431, U432, U433, U434, U435, U436, U437, U438, U439, U440, U441, U442, U443, U444, U445, U446, U447, U448, U449, U450, U451, U452, U453, U454, U455, U456, U457, U458, U459, U460, U461, U462, U463, U464, U465, U466, U467, U468, U469, U470, U471, U472, U473, U474, U475, U476, U477, U478, U479, U480, U481, U482, U483, U484, U485, U486, U487, U488, U489, U490, U491, U492, U493, U494, U495, U496, U497, U498, U499, U500, U501, U502, U503, U504, U505, U506, U507, U508, U509, U510, U511, U512, U513, U514, U515, U516, U517, U518, U519, U520, U521, U522, U523, U524, U525, U526, U527, U528, U529, U530, U531, U532, U533, U534, U535, U536, U537, U538, U539, U540, U541, U542, U543, U544, U545, U546, U547, U548, U549, U550, U551, U552, U553, U554, U555, U556, U557, U558, U559, U560, U561, U562, U563, U564, U565, U566, U567, U568, U569, U570, U571, U572, U573, U574, U575, U576, U577, U578, U579, U580, U581, U582, U583, U584, U585, U586, U587, U588, U589, U590, U591, U592, U593, U594, U595, U596, U597, U598, U599, U600, U601, U602, U603, U604, U605, U606, U607, U608, U609, U610, U611, U612, U613, U614, U615, U616, U617, U618, U619, U620, U621, U622, U623, U624, U625, U626, U627, U628, U629, U630, U631, U632, U633, U634, U635, U636, U637, U638, U639, U640, U641, U642, U643, U644, U645, U646, U647, U648, U649, U650, U651, U652, U653, U654, U655, U656, U657, U658, U659, U660, U661, U662, U663, U664, U665, U666, U667, U668, U669, U670, U671, U672, U673, U674, U675, U676, U677, U678, U679, U680, U681, U682, U683, U684, U685, U686, U687, U688, U689, U690, U691, U692, U693, U694, U695, U696, U697, U698, U699, U700, U701, U702, U703, U704, U705, U706, U707, U708, U709, U710, U711, U712, U713, U714, U715, U716, U717, U718, U719, U720, U721, U722, U723, U724, U725, U726, U727, U728, U729, U730, U731, U732, U733, U734, U735, U736, P3_U2352, P3_U2353, P3_U2354, P3_U2355, P3_U2356, P3_U2357, P3_U2358, P3_U2359, P3_U2360, P3_U2361, P3_U2362, P3_U2363, P3_U2364, P3_U2365, P3_U2366, P3_U2367, P3_U2368, P3_U2369, P3_U2370, P3_U2371, P3_U2372, P3_U2373, P3_U2374, P3_U2375, P3_U2376, P3_U2377, P3_U2378, P3_U2379, P3_U2380, P3_U2381, P3_U2382, P3_U2383, P3_U2384, P3_U2385, P3_U2386, P3_U2387, P3_U2388, P3_U2389, P3_U2390, P3_U2391, P3_U2392, P3_U2393, P3_U2394, P3_U2395, P3_U2396, P3_U2397, P3_U2398, P3_U2399, P3_U2400, P3_U2401, P3_U2402, P3_U2403, P3_U2404, P3_U2405, P3_U2406, P3_U2407, P3_U2408, P3_U2409, P3_U2410, P3_U2411, P3_U2412, P3_U2413, P3_U2414, P3_U2415, P3_U2416, P3_U2417, P3_U2418, P3_U2419, P3_U2420, P3_U2421, P3_U2422, P3_U2423, P3_U2424, P3_U2425, P3_U2426, P3_U2427, P3_U2428, P3_U2429, P3_U2430, P3_U2431, P3_U2432, P3_U2433, P3_U2434, P3_U2435, P3_U2436, P3_U2437, P3_U2438, P3_U2439, P3_U2440, P3_U2441, P3_U2442, P3_U2443, P3_U2444, P3_U2445, P3_U2446, P3_U2447, P3_U2448, P3_U2449, P3_U2450, P3_U2451, P3_U2452, P3_U2453, P3_U2454, P3_U2455, P3_U2456, P3_U2457, P3_U2458, P3_U2459, P3_U2460, P3_U2461, P3_U2462, P3_U2463, P3_U2464, P3_U2465, P3_U2466, P3_U2467, P3_U2468, P3_U2469, P3_U2470, P3_U2471, P3_U2472, P3_U2473, P3_U2474, P3_U2475, P3_U2476, P3_U2477, P3_U2478, P3_U2479, P3_U2480, P3_U2481, P3_U2482, P3_U2483, P3_U2484, P3_U2485, P3_U2486, P3_U2487, P3_U2488, P3_U2489, P3_U2490, P3_U2491, P3_U2492, P3_U2493, P3_U2494, P3_U2495, P3_U2496, P3_U2497, P3_U2498, P3_U2499, P3_U2500, P3_U2501, P3_U2502, P3_U2503, P3_U2504, P3_U2505, P3_U2506, P3_U2507, P3_U2508, P3_U2509, P3_U2510, P3_U2511, P3_U2512, P3_U2513, P3_U2514, P3_U2515, P3_U2516, P3_U2517, P3_U2518, P3_U2519, P3_U2520, P3_U2521, P3_U2522, P3_U2523, P3_U2524, P3_U2525, P3_U2526, P3_U2527, P3_U2528, P3_U2529, P3_U2530, P3_U2531, P3_U2532, P3_U2533, P3_U2534, P3_U2535, P3_U2536, P3_U2537, P3_U2538, P3_U2539, P3_U2540, P3_U2541, P3_U2542, P3_U2543, P3_U2544, P3_U2545, P3_U2546, P3_U2547, P3_U2548, P3_U2549, P3_U2550, P3_U2551, P3_U2552, P3_U2553, P3_U2554, P3_U2555, P3_U2556, P3_U2557, P3_U2558, P3_U2559, P3_U2560, P3_U2561, P3_U2562, P3_U2563, P3_U2564, P3_U2565, P3_U2566, P3_U2567, P3_U2568, P3_U2569, P3_U2570, P3_U2571, P3_U2572, P3_U2573, P3_U2574, P3_U2575, P3_U2576, P3_U2577, P3_U2578, P3_U2579, P3_U2580, P3_U2581, P3_U2582, P3_U2583, P3_U2584, P3_U2585, P3_U2586, P3_U2587, P3_U2588, P3_U2589, P3_U2590, P3_U2591, P3_U2592, P3_U2593, P3_U2594, P3_U2595, P3_U2596, P3_U2597, P3_U2598, P3_U2599, P3_U2600, P3_U2601, P3_U2602, P3_U2603, P3_U2604, P3_U2605, P3_U2606, P3_U2607, P3_U2608, P3_U2609, P3_U2610, P3_U2611, P3_U2612, P3_U2613, P3_U2614, P3_U2615, P3_U2616, P3_U2617, P3_U2618, P3_U2619, P3_U2620, P3_U2621, P3_U2622, P3_U2623, P3_U2624, P3_U2625, P3_U2626, P3_U2627, P3_U2628, P3_U2629, P3_U2630, P3_U2631, P3_U2632, P3_U3062, P3_U3063, P3_U3064, P3_U3065, P3_U3066, P3_U3067, P3_U3068, P3_U3069, P3_U3070, P3_U3071, P3_U3072, P3_U3073, P3_U3074, P3_U3075, P3_U3076, P3_U3077, P3_U3078, P3_U3079, P3_U3080, P3_U3081, P3_U3082, P3_U3083, P3_U3084, P3_U3085, P3_U3086, P3_U3087, P3_U3088, P3_U3089, P3_U3090, P3_U3091, P3_U3092, P3_U3093, P3_U3094, P3_U3095, P3_U3096, P3_U3097, P3_U3098, P3_U3099, P3_U3100, P3_U3101, P3_U3102, P3_U3103, P3_U3104, P3_U3105, P3_U3106, P3_U3107, P3_U3108, P3_U3109, P3_U3110, P3_U3111, P3_U3112, P3_U3113, P3_U3114, P3_U3115, P3_U3116, P3_U3117, P3_U3118, P3_U3119, P3_U3120, P3_U3121, P3_U3122, P3_U3123, P3_U3124, P3_U3125, P3_U3126, P3_U3127, P3_U3128, P3_U3129, P3_U3130, P3_U3131, P3_U3132, P3_U3133, P3_U3134, P3_U3135, P3_U3136, P3_U3137, P3_U3138, P3_U3139, P3_U3140, P3_U3141, P3_U3142, P3_U3143, P3_U3144, P3_U3145, P3_U3146, P3_U3147, P3_U3148, P3_U3149, P3_U3150, P3_U3151, P3_U3152, P3_U3153, P3_U3154, P3_U3155, P3_U3156, P3_U3157, P3_U3158, P3_U3159, P3_U3160, P3_U3161, P3_U3162, P3_U3163, P3_U3164, P3_U3165, P3_U3166, P3_U3167, P3_U3168, P3_U3169, P3_U3170, P3_U3171, P3_U3172, P3_U3173, P3_U3174, P3_U3175, P3_U3176, P3_U3177, P3_U3178, P3_U3179, P3_U3180, P3_U3181, P3_U3182, P3_U3183, P3_U3184, P3_U3185, P3_U3186, P3_U3187, P3_U3188, P3_U3189, P3_U3190, P3_U3191, P3_U3192, P3_U3193, P3_U3194, P3_U3195, P3_U3196, P3_U3197, P3_U3198, P3_U3199, P3_U3200, P3_U3201, P3_U3202, P3_U3203, P3_U3204, P3_U3205, P3_U3206, P3_U3207, P3_U3208, P3_U3209, P3_U3210, P3_U3211, P3_U3212, P3_U3213, P3_U3214, P3_U3215, P3_U3216, P3_U3217, P3_U3218, P3_U3219, P3_U3220, P3_U3221, P3_U3222, P3_U3223, P3_U3224, P3_U3225, P3_U3226, P3_U3227, P3_U3228, P3_U3229, P3_U3230, P3_U3231, P3_U3232, P3_U3233, P3_U3234, P3_U3235, P3_U3236, P3_U3237, P3_U3238, P3_U3239, P3_U3240, P3_U3241, P3_U3242, P3_U3243, P3_U3244, P3_U3245, P3_U3246, P3_U3247, P3_U3248, P3_U3249, P3_U3250, P3_U3251, P3_U3252, P3_U3253, P3_U3254, P3_U3255, P3_U3256, P3_U3257, P3_U3258, P3_U3259, P3_U3260, P3_U3261, P3_U3262, P3_U3263, P3_U3264, P3_U3265, P3_U3266, P3_U3267, P3_U3268, P3_U3269, P3_U3270, P3_U3271, P3_U3272, P3_U3273, P3_U3278, P3_U3279, P3_U3283, P3_U3286, P3_U3287, P3_U3291, P3_U3300, P3_U3301, P3_U3302, P3_U3303, P3_U3304, P3_U3305, P3_U3306, P3_U3307, P3_U3308, P3_U3309, P3_U3310, P3_U3311, P3_U3312, P3_U3313, P3_U3314, P3_U3315, P3_U3316, P3_U3317, P3_U3318, P3_U3319, P3_U3320, P3_U3321, P3_U3322, P3_U3323, P3_U3324, P3_U3325, P3_U3326, P3_U3327, P3_U3328, P3_U3329, P3_U3330, P3_U3331, P3_U3332, P3_U3333, P3_U3334, P3_U3335, P3_U3336, P3_U3337, P3_U3338, P3_U3339, P3_U3340, P3_U3341, P3_U3342, P3_U3343, P3_U3344, P3_U3345, P3_U3346, P3_U3347, P3_U3348, P3_U3349, P3_U3350, P3_U3351, P3_U3352, P3_U3353, P3_U3354, P3_U3355, P3_U3356, P3_U3357, P3_U3358, P3_U3359, P3_U3360, P3_U3361, P3_U3362, P3_U3363, P3_U3364, P3_U3365, P3_U3366, P3_U3367, P3_U3368, P3_U3369, P3_U3370, P3_U3371, P3_U3372, P3_U3373, P3_U3374, P3_U3375, P3_U3376, P3_U3377, P3_U3378, P3_U3379, P3_U3380, P3_U3381, P3_U3382, P3_U3383, P3_U3384, P3_U3385, P3_U3386, P3_U3387, P3_U3388, P3_U3389, P3_U3390, P3_U3391, P3_U3392, P3_U3393, P3_U3394, P3_U3395, P3_U3396, P3_U3397, P3_U3398, P3_U3399, P3_U3400, P3_U3401, P3_U3402, P3_U3403, P3_U3404, P3_U3405, P3_U3406, P3_U3407, P3_U3408, P3_U3409, P3_U3410, P3_U3411, P3_U3412, P3_U3413, P3_U3414, P3_U3415, P3_U3416, P3_U3417, P3_U3418, P3_U3419, P3_U3420, P3_U3421, P3_U3422, P3_U3423, P3_U3424, P3_U3425, P3_U3426, P3_U3427, P3_U3428, P3_U3429, P3_U3430, P3_U3431, P3_U3432, P3_U3433, P3_U3434, P3_U3435, P3_U3436, P3_U3437, P3_U3438, P3_U3439, P3_U3440, P3_U3441, P3_U3442, P3_U3443, P3_U3444, P3_U3445, P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3523, P3_U3524, P3_U3525, P3_U3526, P3_U3527, P3_U3528, P3_U3529, P3_U3530, P3_U3531, P3_U3532, P3_U3533, P3_U3534, P3_U3535, P3_U3536, P3_U3537, P3_U3538, P3_U3539, P3_U3540, P3_U3541, P3_U3542, P3_U3543, P3_U3544, P3_U3545, P3_U3546, P3_U3547, P3_U3548, P3_U3549, P3_U3550, P3_U3551, P3_U3552, P3_U3553, P3_U3554, P3_U3555, P3_U3556, P3_U3557, P3_U3558, P3_U3559, P3_U3560, P3_U3561, P3_U3562, P3_U3563, P3_U3564, P3_U3565, P3_U3566, P3_U3567, P3_U3568, P3_U3569, P3_U3570, P3_U3571, P3_U3572, P3_U3573, P3_U3574, P3_U3575, P3_U3576, P3_U3577, P3_U3578, P3_U3579, P3_U3580, P3_U3581, P3_U3582, P3_U3583, P3_U3584, P3_U3585, P3_U3586, P3_U3587, P3_U3588, P3_U3589, P3_U3590, P3_U3591, P3_U3592, P3_U3593, P3_U3594, P3_U3595, P3_U3596, P3_U3597, P3_U3598, P3_U3599, P3_U3600, P3_U3601, P3_U3602, P3_U3603, P3_U3604, P3_U3605, P3_U3606, P3_U3607, P3_U3608, P3_U3609, P3_U3610, P3_U3611, P3_U3612, P3_U3613, P3_U3614, P3_U3615, P3_U3616, P3_U3617, P3_U3618, P3_U3619, P3_U3620, P3_U3621, P3_U3622, P3_U3623, P3_U3624, P3_U3625, P3_U3626, P3_U3627, P3_U3628, P3_U3629, P3_U3630, P3_U3631, P3_U3632, P3_U3633, P3_U3634, P3_U3635, P3_U3636, P3_U3637, P3_U3638, P3_U3639, P3_U3640, P3_U3641, P3_U3642, P3_U3643, P3_U3644, P3_U3645, P3_U3646, P3_U3647, P3_U3648, P3_U3649, P3_U3650, P3_U3651, P3_U3652, P3_U3653, P3_U3654, P3_U3655, P3_U3656, P3_U3657, P3_U3658, P3_U3659, P3_U3660, P3_U3661, P3_U3662, P3_U3663, P3_U3664, P3_U3665, P3_U3666, P3_U3667, P3_U3668, P3_U3669, P3_U3670, P3_U3671, P3_U3672, P3_U3673, P3_U3674, P3_U3675, P3_U3676, P3_U3677, P3_U3678, P3_U3679, P3_U3680, P3_U3681, P3_U3682, P3_U3683, P3_U3684, P3_U3685, P3_U3686, P3_U3687, P3_U3688, P3_U3689, P3_U3690, P3_U3691, P3_U3692, P3_U3693, P3_U3694, P3_U3695, P3_U3696, P3_U3697, P3_U3698, P3_U3699, P3_U3700, P3_U3701, P3_U3702, P3_U3703, P3_U3704, P3_U3705, P3_U3706, P3_U3707, P3_U3708, P3_U3709, P3_U3710, P3_U3711, P3_U3712, P3_U3713, P3_U3714, P3_U3715, P3_U3716, P3_U3717, P3_U3718, P3_U3719, P3_U3720, P3_U3721, P3_U3722, P3_U3723, P3_U3724, P3_U3725, P3_U3726, P3_U3727, P3_U3728, P3_U3729, P3_U3730, P3_U3731, P3_U3732, P3_U3733, P3_U3734, P3_U3735, P3_U3736, P3_U3737, P3_U3738, P3_U3739, P3_U3740, P3_U3741, P3_U3742, P3_U3743, P3_U3744, P3_U3745, P3_U3746, P3_U3747, P3_U3748, P3_U3749, P3_U3750, P3_U3751, P3_U3752, P3_U3753, P3_U3754, P3_U3755, P3_U3756, P3_U3757, P3_U3758, P3_U3759, P3_U3760, P3_U3761, P3_U3762, P3_U3763, P3_U3764, P3_U3765, P3_U3766, P3_U3767, P3_U3768, P3_U3769, P3_U3770, P3_U3771, P3_U3772, P3_U3773, P3_U3774, P3_U3775, P3_U3776, P3_U3777, P3_U3778, P3_U3779, P3_U3780, P3_U3781, P3_U3782, P3_U3783, P3_U3784, P3_U3785, P3_U3786, P3_U3787, P3_U3788, P3_U3789, P3_U3790, P3_U3791, P3_U3792, P3_U3793, P3_U3794, P3_U3795, P3_U3796, P3_U3797, P3_U3798, P3_U3799, P3_U3800, P3_U3801, P3_U3802, P3_U3803, P3_U3804, P3_U3805, P3_U3806, P3_U3807, P3_U3808, P3_U3809, P3_U3810, P3_U3811, P3_U3812, P3_U3813, P3_U3814, P3_U3815, P3_U3816, P3_U3817, P3_U3818, P3_U3819, P3_U3820, P3_U3821, P3_U3822, P3_U3823, P3_U3824, P3_U3825, P3_U3826, P3_U3827, P3_U3828, P3_U3829, P3_U3830, P3_U3831, P3_U3832, P3_U3833, P3_U3834, P3_U3835, P3_U3836, P3_U3837, P3_U3838, P3_U3839, P3_U3840, P3_U3841, P3_U3842, P3_U3843, P3_U3844, P3_U3845, P3_U3846, P3_U3847, P3_U3848, P3_U3849, P3_U3850, P3_U3851, P3_U3852, P3_U3853, P3_U3854, P3_U3855, P3_U3856, P3_U3857, P3_U3858, P3_U3859, P3_U3860, P3_U3861, P3_U3862, P3_U3863, P3_U3864, P3_U3865, P3_U3866, P3_U3867, P3_U3868, P3_U3869, P3_U3870, P3_U3871, P3_U3872, P3_U3873, P3_U3874, P3_U3875, P3_U3876, P3_U3877, P3_U3878, P3_U3879, P3_U3880, P3_U3881, P3_U3882, P3_U3883, P3_U3884, P3_U3885, P3_U3886, P3_U3887, P3_U3888, P3_U3889, P3_U3890, P3_U3891, P3_U3892, P3_U3893, P3_U3894, P3_U3895, P3_U3896, P3_U3897, P3_U3898, P3_U3899, P3_U3900, P3_U3901, P3_U3902, P3_U3903, P3_U3904, P3_U3905, P3_U3906, P3_U3907, P3_U3908, P3_U3909, P3_U3910, P3_U3911, P3_U3912, P3_U3913, P3_U3914, P3_U3915, P3_U3916, P3_U3917, P3_U3918, P3_U3919, P3_U3920, P3_U3921, P3_U3922, P3_U3923, P3_U3924, P3_U3925, P3_U3926, P3_U3927, P3_U3928, P3_U3929, P3_U3930, P3_U3931, P3_U3932, P3_U3933, P3_U3934, P3_U3935, P3_U3936, P3_U3937, P3_U3938, P3_U3939, P3_U3940, P3_U3941, P3_U3942, P3_U3943, P3_U3944, P3_U3945, P3_U3946, P3_U3947, P3_U3948, P3_U3949, P3_U3950, P3_U3951, P3_U3952, P3_U3953, P3_U3954, P3_U3955, P3_U3956, P3_U3957, P3_U3958, P3_U3959, P3_U3960, P3_U3961, P3_U3962, P3_U3963, P3_U3964, P3_U3965, P3_U3966, P3_U3967, P3_U3968, P3_U3969, P3_U3970, P3_U3971, P3_U3972, P3_U3973, P3_U3974, P3_U3975, P3_U3976, P3_U3977, P3_U3978, P3_U3979, P3_U3980, P3_U3981, P3_U3982, P3_U3983, P3_U3984, P3_U3985, P3_U3986, P3_U3987, P3_U3988, P3_U3989, P3_U3990, P3_U3991, P3_U3992, P3_U3993, P3_U3994, P3_U3995, P3_U3996, P3_U3997, P3_U3998, P3_U3999, P3_U4000, P3_U4001, P3_U4002, P3_U4003, P3_U4004, P3_U4005, P3_U4006, P3_U4007, P3_U4008, P3_U4009, P3_U4010, P3_U4011, P3_U4012, P3_U4013, P3_U4014, P3_U4015, P3_U4016, P3_U4017, P3_U4018, P3_U4019, P3_U4020, P3_U4021, P3_U4022, P3_U4023, P3_U4024, P3_U4025, P3_U4026, P3_U4027, P3_U4028, P3_U4029, P3_U4030, P3_U4031, P3_U4032, P3_U4033, P3_U4034, P3_U4035, P3_U4036, P3_U4037, P3_U4038, P3_U4039, P3_U4040, P3_U4041, P3_U4042, P3_U4043, P3_U4044, P3_U4045, P3_U4046, P3_U4047, P3_U4048, P3_U4049, P3_U4050, P3_U4051, P3_U4052, P3_U4053, P3_U4054, P3_U4055, P3_U4056, P3_U4057, P3_U4058, P3_U4059, P3_U4060, P3_U4061, P3_U4062, P3_U4063, P3_U4064, P3_U4065, P3_U4066, P3_U4067, P3_U4068, P3_U4069, P3_U4070, P3_U4071, P3_U4072, P3_U4073, P3_U4074, P3_U4075, P3_U4076, P3_U4077, P3_U4078, P3_U4079, P3_U4080, P3_U4081, P3_U4082, P3_U4083, P3_U4084, P3_U4085, P3_U4086, P3_U4087, P3_U4088, P3_U4089, P3_U4090, P3_U4091, P3_U4092, P3_U4093, P3_U4094, P3_U4095, P3_U4096, P3_U4097, P3_U4098, P3_U4099, P3_U4100, P3_U4101, P3_U4102, P3_U4103, P3_U4104, P3_U4105, P3_U4106, P3_U4107, P3_U4108, P3_U4109, P3_U4110, P3_U4111, P3_U4112, P3_U4113, P3_U4114, P3_U4115, P3_U4116, P3_U4117, P3_U4118, P3_U4119, P3_U4120, P3_U4121, P3_U4122, P3_U4123, P3_U4124, P3_U4125, P3_U4126, P3_U4127, P3_U4128, P3_U4129, P3_U4130, P3_U4131, P3_U4132, P3_U4133, P3_U4134, P3_U4135, P3_U4136, P3_U4137, P3_U4138, P3_U4139, P3_U4140, P3_U4141, P3_U4142, P3_U4143, P3_U4144, P3_U4145, P3_U4146, P3_U4147, P3_U4148, P3_U4149, P3_U4150, P3_U4151, P3_U4152, P3_U4153, P3_U4154, P3_U4155, P3_U4156, P3_U4157, P3_U4158, P3_U4159, P3_U4160, P3_U4161, P3_U4162, P3_U4163, P3_U4164, P3_U4165, P3_U4166, P3_U4167, P3_U4168, P3_U4169, P3_U4170, P3_U4171, P3_U4172, P3_U4173, P3_U4174, P3_U4175, P3_U4176, P3_U4177, P3_U4178, P3_U4179, P3_U4180, P3_U4181, P3_U4182, P3_U4183, P3_U4184, P3_U4185, P3_U4186, P3_U4187, P3_U4188, P3_U4189, P3_U4190, P3_U4191, P3_U4192, P3_U4193, P3_U4194, P3_U4195, P3_U4196, P3_U4197, P3_U4198, P3_U4199, P3_U4200, P3_U4201, P3_U4202, P3_U4203, P3_U4204, P3_U4205, P3_U4206, P3_U4207, P3_U4208, P3_U4209, P3_U4210, P3_U4211, P3_U4212, P3_U4213, P3_U4214, P3_U4215, P3_U4216, P3_U4217, P3_U4218, P3_U4219, P3_U4220, P3_U4221, P3_U4222, P3_U4223, P3_U4224, P3_U4225, P3_U4226, P3_U4227, P3_U4228, P3_U4229, P3_U4230, P3_U4231, P3_U4232, P3_U4233, P3_U4234, P3_U4235, P3_U4236, P3_U4237, P3_U4238, P3_U4239, P3_U4240, P3_U4241, P3_U4242, P3_U4243, P3_U4244, P3_U4245, P3_U4246, P3_U4247, P3_U4248, P3_U4249, P3_U4250, P3_U4251, P3_U4252, P3_U4253, P3_U4254, P3_U4255, P3_U4256, P3_U4257, P3_U4258, P3_U4259, P3_U4260, P3_U4261, P3_U4262, P3_U4263, P3_U4264, P3_U4265, P3_U4266, P3_U4267, P3_U4268, P3_U4269, P3_U4270, P3_U4271, P3_U4272, P3_U4273, P3_U4274, P3_U4275, P3_U4276, P3_U4277, P3_U4278, P3_U4279, P3_U4280, P3_U4281, P3_U4282, P3_U4283, P3_U4284, P3_U4285, P3_U4286, P3_U4287, P3_U4288, P3_U4289, P3_U4290, P3_U4291, P3_U4292, P3_U4293, P3_U4294, P3_U4295, P3_U4296, P3_U4297, P3_U4298, P3_U4299, P3_U4300, P3_U4301, P3_U4302, P3_U4303, P3_U4304, P3_U4305, P3_U4306, P3_U4307, P3_U4308, P3_U4309, P3_U4310, P3_U4311, P3_U4312, P3_U4313, P3_U4314, P3_U4315, P3_U4316, P3_U4317, P3_U4318, P3_U4319, P3_U4320, P3_U4321, P3_U4322, P3_U4323, P3_U4324, P3_U4325, P3_U4326, P3_U4327, P3_U4328, P3_U4329, P3_U4330, P3_U4331, P3_U4332, P3_U4333, P3_U4334, P3_U4335, P3_U4336, P3_U4337, P3_U4338, P3_U4339, P3_U4340, P3_U4341, P3_U4342, P3_U4343, P3_U4344, P3_U4345, P3_U4346, P3_U4347, P3_U4348, P3_U4349, P3_U4350, P3_U4351, P3_U4352, P3_U4353, P3_U4354, P3_U4355, P3_U4356, P3_U4357, P3_U4358, P3_U4359, P3_U4360, P3_U4361, P3_U4362, P3_U4363, P3_U4364, P3_U4365, P3_U4366, P3_U4367, P3_U4368, P3_U4369, P3_U4370, P3_U4371, P3_U4372, P3_U4373, P3_U4374, P3_U4375, P3_U4376, P3_U4377, P3_U4378, P3_U4379, P3_U4380, P3_U4381, P3_U4382, P3_U4383, P3_U4384, P3_U4385, P3_U4386, P3_U4387, P3_U4388, P3_U4389, P3_U4390, P3_U4391, P3_U4392, P3_U4393, P3_U4394, P3_U4395, P3_U4396, P3_U4397, P3_U4398, P3_U4399, P3_U4400, P3_U4401, P3_U4402, P3_U4403, P3_U4404, P3_U4405, P3_U4406, P3_U4407, P3_U4408, P3_U4409, P3_U4410, P3_U4411, P3_U4412, P3_U4413, P3_U4414, P3_U4415, P3_U4416, P3_U4417, P3_U4418, P3_U4419, P3_U4420, P3_U4421, P3_U4422, P3_U4423, P3_U4424, P3_U4425, P3_U4426, P3_U4427, P3_U4428, P3_U4429, P3_U4430, P3_U4431, P3_U4432, P3_U4433, P3_U4434, P3_U4435, P3_U4436, P3_U4437, P3_U4438, P3_U4439, P3_U4440, P3_U4441, P3_U4442, P3_U4443, P3_U4444, P3_U4445, P3_U4446, P3_U4447, P3_U4448, P3_U4449, P3_U4450, P3_U4451, P3_U4452, P3_U4453, P3_U4454, P3_U4455, P3_U4456, P3_U4457, P3_U4458, P3_U4459, P3_U4460, P3_U4461, P3_U4462, P3_U4463, P3_U4464, P3_U4465, P3_U4466, P3_U4467, P3_U4468, P3_U4469, P3_U4470, P3_U4471, P3_U4472, P3_U4473, P3_U4474, P3_U4475, P3_U4476, P3_U4477, P3_U4478, P3_U4479, P3_U4480, P3_U4481, P3_U4482, P3_U4483, P3_U4484, P3_U4485, P3_U4486, P3_U4487, P3_U4488, P3_U4489, P3_U4490, P3_U4491, P3_U4492, P3_U4493, P3_U4494, P3_U4495, P3_U4496, P3_U4497, P3_U4498, P3_U4499, P3_U4500, P3_U4501, P3_U4502, P3_U4503, P3_U4504, P3_U4505, P3_U4506, P3_U4507, P3_U4508, P3_U4509, P3_U4510, P3_U4511, P3_U4512, P3_U4513, P3_U4514, P3_U4515, P3_U4516, P3_U4517, P3_U4518, P3_U4519, P3_U4520, P3_U4521, P3_U4522, P3_U4523, P3_U4524, P3_U4525, P3_U4526, P3_U4527, P3_U4528, P3_U4529, P3_U4530, P3_U4531, P3_U4532, P3_U4533, P3_U4534, P3_U4535, P3_U4536, P3_U4537, P3_U4538, P3_U4539, P3_U4540, P3_U4541, P3_U4542, P3_U4543, P3_U4544, P3_U4545, P3_U4546, P3_U4547, P3_U4548, P3_U4549, P3_U4550, P3_U4551, P3_U4552, P3_U4553, P3_U4554, P3_U4555, P3_U4556, P3_U4557, P3_U4558, P3_U4559, P3_U4560, P3_U4561, P3_U4562, P3_U4563, P3_U4564, P3_U4565, P3_U4566, P3_U4567, P3_U4568, P3_U4569, P3_U4570, P3_U4571, P3_U4572, P3_U4573, P3_U4574, P3_U4575, P3_U4576, P3_U4577, P3_U4578, P3_U4579, P3_U4580, P3_U4581, P3_U4582, P3_U4583, P3_U4584, P3_U4585, P3_U4586, P3_U4587, P3_U4588, P3_U4589, P3_U4590, P3_U4591, P3_U4592, P3_U4593, P3_U4594, P3_U4595, P3_U4596, P3_U4597, P3_U4598, P3_U4599, P3_U4600, P3_U4601, P3_U4602, P3_U4603, P3_U4604, P3_U4605, P3_U4606, P3_U4607, P3_U4608, P3_U4609, P3_U4610, P3_U4611, P3_U4612, P3_U4613, P3_U4614, P3_U4615, P3_U4616, P3_U4617, P3_U4618, P3_U4619, P3_U4620, P3_U4621, P3_U4622, P3_U4623, P3_U4624, P3_U4625, P3_U4626, P3_U4627, P3_U4628, P3_U4629, P3_U4630, P3_U4631, P3_U4632, P3_U4633, P3_U4634, P3_U4635, P3_U4636, P3_U4637, P3_U4638, P3_U4639, P3_U4640, P3_U4641, P3_U4642, P3_U4643, P3_U4644, P3_U4645, P3_U4646, P3_U4647, P3_U4648, P3_U4649, P3_U4650, P3_U4651, P3_U4652, P3_U4653, P3_U4654, P3_U4655, P3_U4656, P3_U4657, P3_U4658, P3_U4659, P3_U4660, P3_U4661, P3_U4662, P3_U4663, P3_U4664, P3_U4665, P3_U4666, P3_U4667, P3_U4668, P3_U4669, P3_U4670, P3_U4671, P3_U4672, P3_U4673, P3_U4674, P3_U4675, P3_U4676, P3_U4677, P3_U4678, P3_U4679, P3_U4680, P3_U4681, P3_U4682, P3_U4683, P3_U4684, P3_U4685, P3_U4686, P3_U4687, P3_U4688, P3_U4689, P3_U4690, P3_U4691, P3_U4692, P3_U4693, P3_U4694, P3_U4695, P3_U4696, P3_U4697, P3_U4698, P3_U4699, P3_U4700, P3_U4701, P3_U4702, P3_U4703, P3_U4704, P3_U4705, P3_U4706, P3_U4707, P3_U4708, P3_U4709, P3_U4710, P3_U4711, P3_U4712, P3_U4713, P3_U4714, P3_U4715, P3_U4716, P3_U4717, P3_U4718, P3_U4719, P3_U4720, P3_U4721, P3_U4722, P3_U4723, P3_U4724, P3_U4725, P3_U4726, P3_U4727, P3_U4728, P3_U4729, P3_U4730, P3_U4731, P3_U4732, P3_U4733, P3_U4734, P3_U4735, P3_U4736, P3_U4737, P3_U4738, P3_U4739, P3_U4740, P3_U4741, P3_U4742, P3_U4743, P3_U4744, P3_U4745, P3_U4746, P3_U4747, P3_U4748, P3_U4749, P3_U4750, P3_U4751, P3_U4752, P3_U4753, P3_U4754, P3_U4755, P3_U4756, P3_U4757, P3_U4758, P3_U4759, P3_U4760, P3_U4761, P3_U4762, P3_U4763, P3_U4764, P3_U4765, P3_U4766, P3_U4767, P3_U4768, P3_U4769, P3_U4770, P3_U4771, P3_U4772, P3_U4773, P3_U4774, P3_U4775, P3_U4776, P3_U4777, P3_U4778, P3_U4779, P3_U4780, P3_U4781, P3_U4782, P3_U4783, P3_U4784, P3_U4785, P3_U4786, P3_U4787, P3_U4788, P3_U4789, P3_U4790, P3_U4791, P3_U4792, P3_U4793, P3_U4794, P3_U4795, P3_U4796, P3_U4797, P3_U4798, P3_U4799, P3_U4800, P3_U4801, P3_U4802, P3_U4803, P3_U4804, P3_U4805, P3_U4806, P3_U4807, P3_U4808, P3_U4809, P3_U4810, P3_U4811, P3_U4812, P3_U4813, P3_U4814, P3_U4815, P3_U4816, P3_U4817, P3_U4818, P3_U4819, P3_U4820, P3_U4821, P3_U4822, P3_U4823, P3_U4824, P3_U4825, P3_U4826, P3_U4827, P3_U4828, P3_U4829, P3_U4830, P3_U4831, P3_U4832, P3_U4833, P3_U4834, P3_U4835, P3_U4836, P3_U4837, P3_U4838, P3_U4839, P3_U4840, P3_U4841, P3_U4842, P3_U4843, P3_U4844, P3_U4845, P3_U4846, P3_U4847, P3_U4848, P3_U4849, P3_U4850, P3_U4851, P3_U4852, P3_U4853, P3_U4854, P3_U4855, P3_U4856, P3_U4857, P3_U4858, P3_U4859, P3_U4860, P3_U4861, P3_U4862, P3_U4863, P3_U4864, P3_U4865, P3_U4866, P3_U4867, P3_U4868, P3_U4869, P3_U4870, P3_U4871, P3_U4872, P3_U4873, P3_U4874, P3_U4875, P3_U4876, P3_U4877, P3_U4878, P3_U4879, P3_U4880, P3_U4881, P3_U4882, P3_U4883, P3_U4884, P3_U4885, P3_U4886, P3_U4887, P3_U4888, P3_U4889, P3_U4890, P3_U4891, P3_U4892, P3_U4893, P3_U4894, P3_U4895, P3_U4896, P3_U4897, P3_U4898, P3_U4899, P3_U4900, P3_U4901, P3_U4902, P3_U4903, P3_U4904, P3_U4905, P3_U4906, P3_U4907, P3_U4908, P3_U4909, P3_U4910, P3_U4911, P3_U4912, P3_U4913, P3_U4914, P3_U4915, P3_U4916, P3_U4917, P3_U4918, P3_U4919, P3_U4920, P3_U4921, P3_U4922, P3_U4923, P3_U4924, P3_U4925, P3_U4926, P3_U4927, P3_U4928, P3_U4929, P3_U4930, P3_U4931, P3_U4932, P3_U4933, P3_U4934, P3_U4935, P3_U4936, P3_U4937, P3_U4938, P3_U4939, P3_U4940, P3_U4941, P3_U4942, P3_U4943, P3_U4944, P3_U4945, P3_U4946, P3_U4947, P3_U4948, P3_U4949, P3_U4950, P3_U4951, P3_U4952, P3_U4953, P3_U4954, P3_U4955, P3_U4956, P3_U4957, P3_U4958, P3_U4959, P3_U4960, P3_U4961, P3_U4962, P3_U4963, P3_U4964, P3_U4965, P3_U4966, P3_U4967, P3_U4968, P3_U4969, P3_U4970, P3_U4971, P3_U4972, P3_U4973, P3_U4974, P3_U4975, P3_U4976, P3_U4977, P3_U4978, P3_U4979, P3_U4980, P3_U4981, P3_U4982, P3_U4983, P3_U4984, P3_U4985, P3_U4986, P3_U4987, P3_U4988, P3_U4989, P3_U4990, P3_U4991, P3_U4992, P3_U4993, P3_U4994, P3_U4995, P3_U4996, P3_U4997, P3_U4998, P3_U4999, P3_U5000, P3_U5001, P3_U5002, P3_U5003, P3_U5004, P3_U5005, P3_U5006, P3_U5007, P3_U5008, P3_U5009, P3_U5010, P3_U5011, P3_U5012, P3_U5013, P3_U5014, P3_U5015, P3_U5016, P3_U5017, P3_U5018, P3_U5019, P3_U5020, P3_U5021, P3_U5022, P3_U5023, P3_U5024, P3_U5025, P3_U5026, P3_U5027, P3_U5028, P3_U5029, P3_U5030, P3_U5031, P3_U5032, P3_U5033, P3_U5034, P3_U5035, P3_U5036, P3_U5037, P3_U5038, P3_U5039, P3_U5040, P3_U5041, P3_U5042, P3_U5043, P3_U5044, P3_U5045, P3_U5046, P3_U5047, P3_U5048, P3_U5049, P3_U5050, P3_U5051, P3_U5052, P3_U5053, P3_U5054, P3_U5055, P3_U5056, P3_U5057, P3_U5058, P3_U5059, P3_U5060, P3_U5061, P3_U5062, P3_U5063, P3_U5064, P3_U5065, P3_U5066, P3_U5067, P3_U5068, P3_U5069, P3_U5070, P3_U5071, P3_U5072, P3_U5073, P3_U5074, P3_U5075, P3_U5076, P3_U5077, P3_U5078, P3_U5079, P3_U5080, P3_U5081, P3_U5082, P3_U5083, P3_U5084, P3_U5085, P3_U5086, P3_U5087, P3_U5088, P3_U5089, P3_U5090, P3_U5091, P3_U5092, P3_U5093, P3_U5094, P3_U5095, P3_U5096, P3_U5097, P3_U5098, P3_U5099, P3_U5100, P3_U5101, P3_U5102, P3_U5103, P3_U5104, P3_U5105, P3_U5106, P3_U5107, P3_U5108, P3_U5109, P3_U5110, P3_U5111, P3_U5112, P3_U5113, P3_U5114, P3_U5115, P3_U5116, P3_U5117, P3_U5118, P3_U5119, P3_U5120, P3_U5121, P3_U5122, P3_U5123, P3_U5124, P3_U5125, P3_U5126, P3_U5127, P3_U5128, P3_U5129, P3_U5130, P3_U5131, P3_U5132, P3_U5133, P3_U5134, P3_U5135, P3_U5136, P3_U5137, P3_U5138, P3_U5139, P3_U5140, P3_U5141, P3_U5142, P3_U5143, P3_U5144, P3_U5145, P3_U5146, P3_U5147, P3_U5148, P3_U5149, P3_U5150, P3_U5151, P3_U5152, P3_U5153, P3_U5154, P3_U5155, P3_U5156, P3_U5157, P3_U5158, P3_U5159, P3_U5160, P3_U5161, P3_U5162, P3_U5163, P3_U5164, P3_U5165, P3_U5166, P3_U5167, P3_U5168, P3_U5169, P3_U5170, P3_U5171, P3_U5172, P3_U5173, P3_U5174, P3_U5175, P3_U5176, P3_U5177, P3_U5178, P3_U5179, P3_U5180, P3_U5181, P3_U5182, P3_U5183, P3_U5184, P3_U5185, P3_U5186, P3_U5187, P3_U5188, P3_U5189, P3_U5190, P3_U5191, P3_U5192, P3_U5193, P3_U5194, P3_U5195, P3_U5196, P3_U5197, P3_U5198, P3_U5199, P3_U5200, P3_U5201, P3_U5202, P3_U5203, P3_U5204, P3_U5205, P3_U5206, P3_U5207, P3_U5208, P3_U5209, P3_U5210, P3_U5211, P3_U5212, P3_U5213, P3_U5214, P3_U5215, P3_U5216, P3_U5217, P3_U5218, P3_U5219, P3_U5220, P3_U5221, P3_U5222, P3_U5223, P3_U5224, P3_U5225, P3_U5226, P3_U5227, P3_U5228, P3_U5229, P3_U5230, P3_U5231, P3_U5232, P3_U5233, P3_U5234, P3_U5235, P3_U5236, P3_U5237, P3_U5238, P3_U5239, P3_U5240, P3_U5241, P3_U5242, P3_U5243, P3_U5244, P3_U5245, P3_U5246, P3_U5247, P3_U5248, P3_U5249, P3_U5250, P3_U5251, P3_U5252, P3_U5253, P3_U5254, P3_U5255, P3_U5256, P3_U5257, P3_U5258, P3_U5259, P3_U5260, P3_U5261, P3_U5262, P3_U5263, P3_U5264, P3_U5265, P3_U5266, P3_U5267, P3_U5268, P3_U5269, P3_U5270, P3_U5271, P3_U5272, P3_U5273, P3_U5274, P3_U5275, P3_U5276, P3_U5277, P3_U5278, P3_U5279, P3_U5280, P3_U5281, P3_U5282, P3_U5283, P3_U5284, P3_U5285, P3_U5286, P3_U5287, P3_U5288, P3_U5289, P3_U5290, P3_U5291, P3_U5292, P3_U5293, P3_U5294, P3_U5295, P3_U5296, P3_U5297, P3_U5298, P3_U5299, P3_U5300, P3_U5301, P3_U5302, P3_U5303, P3_U5304, P3_U5305, P3_U5306, P3_U5307, P3_U5308, P3_U5309, P3_U5310, P3_U5311, P3_U5312, P3_U5313, P3_U5314, P3_U5315, P3_U5316, P3_U5317, P3_U5318, P3_U5319, P3_U5320, P3_U5321, P3_U5322, P3_U5323, P3_U5324, P3_U5325, P3_U5326, P3_U5327, P3_U5328, P3_U5329, P3_U5330, P3_U5331, P3_U5332, P3_U5333, P3_U5334, P3_U5335, P3_U5336, P3_U5337, P3_U5338, P3_U5339, P3_U5340, P3_U5341, P3_U5342, P3_U5343, P3_U5344, P3_U5345, P3_U5346, P3_U5347, P3_U5348, P3_U5349, P3_U5350, P3_U5351, P3_U5352, P3_U5353, P3_U5354, P3_U5355, P3_U5356, P3_U5357, P3_U5358, P3_U5359, P3_U5360, P3_U5361, P3_U5362, P3_U5363, P3_U5364, P3_U5365, P3_U5366, P3_U5367, P3_U5368, P3_U5369, P3_U5370, P3_U5371, P3_U5372, P3_U5373, P3_U5374, P3_U5375, P3_U5376, P3_U5377, P3_U5378, P3_U5379, P3_U5380, P3_U5381, P3_U5382, P3_U5383, P3_U5384, P3_U5385, P3_U5386, P3_U5387, P3_U5388, P3_U5389, P3_U5390, P3_U5391, P3_U5392, P3_U5393, P3_U5394, P3_U5395, P3_U5396, P3_U5397, P3_U5398, P3_U5399, P3_U5400, P3_U5401, P3_U5402, P3_U5403, P3_U5404, P3_U5405, P3_U5406, P3_U5407, P3_U5408, P3_U5409, P3_U5410, P3_U5411, P3_U5412, P3_U5413, P3_U5414, P3_U5415, P3_U5416, P3_U5417, P3_U5418, P3_U5419, P3_U5420, P3_U5421, P3_U5422, P3_U5423, P3_U5424, P3_U5425, P3_U5426, P3_U5427, P3_U5428, P3_U5429, P3_U5430, P3_U5431, P3_U5432, P3_U5433, P3_U5434, P3_U5435, P3_U5436, P3_U5437, P3_U5438, P3_U5439, P3_U5440, P3_U5441, P3_U5442, P3_U5443, P3_U5444, P3_U5445, P3_U5446, P3_U5447, P3_U5448, P3_U5449, P3_U5450, P3_U5451, P3_U5452, P3_U5453, P3_U5454, P3_U5455, P3_U5456, P3_U5457, P3_U5458, P3_U5459, P3_U5460, P3_U5461, P3_U5462, P3_U5463, P3_U5464, P3_U5465, P3_U5466, P3_U5467, P3_U5468, P3_U5469, P3_U5470, P3_U5471, P3_U5472, P3_U5473, P3_U5474, P3_U5475, P3_U5476, P3_U5477, P3_U5478, P3_U5479, P3_U5480, P3_U5481, P3_U5482, P3_U5483, P3_U5484, P3_U5485, P3_U5486, P3_U5487, P3_U5488, P3_U5489, P3_U5490, P3_U5491, P3_U5492, P3_U5493, P3_U5494, P3_U5495, P3_U5496, P3_U5497, P3_U5498, P3_U5499, P3_U5500, P3_U5501, P3_U5502, P3_U5503, P3_U5504, P3_U5505, P3_U5506, P3_U5507, P3_U5508, P3_U5509, P3_U5510, P3_U5511, P3_U5512, P3_U5513, P3_U5514, P3_U5515, P3_U5516, P3_U5517, P3_U5518, P3_U5519, P3_U5520, P3_U5521, P3_U5522, P3_U5523, P3_U5524, P3_U5525, P3_U5526, P3_U5527, P3_U5528, P3_U5529, P3_U5530, P3_U5531, P3_U5532, P3_U5533, P3_U5534, P3_U5535, P3_U5536, P3_U5537, P3_U5538, P3_U5539, P3_U5540, P3_U5541, P3_U5542, P3_U5543, P3_U5544, P3_U5545, P3_U5546, P3_U5547, P3_U5548, P3_U5549, P3_U5550, P3_U5551, P3_U5552, P3_U5553, P3_U5554, P3_U5555, P3_U5556, P3_U5557, P3_U5558, P3_U5559, P3_U5560, P3_U5561, P3_U5562, P3_U5563, P3_U5564, P3_U5565, P3_U5566, P3_U5567, P3_U5568, P3_U5569, P3_U5570, P3_U5571, P3_U5572, P3_U5573, P3_U5574, P3_U5575, P3_U5576, P3_U5577, P3_U5578, P3_U5579, P3_U5580, P3_U5581, P3_U5582, P3_U5583, P3_U5584, P3_U5585, P3_U5586, P3_U5587, P3_U5588, P3_U5589, P3_U5590, P3_U5591, P3_U5592, P3_U5593, P3_U5594, P3_U5595, P3_U5596, P3_U5597, P3_U5598, P3_U5599, P3_U5600, P3_U5601, P3_U5602, P3_U5603, P3_U5604, P3_U5605, P3_U5606, P3_U5607, P3_U5608, P3_U5609, P3_U5610, P3_U5611, P3_U5612, P3_U5613, P3_U5614, P3_U5615, P3_U5616, P3_U5617, P3_U5618, P3_U5619, P3_U5620, P3_U5621, P3_U5622, P3_U5623, P3_U5624, P3_U5625, P3_U5626, P3_U5627, P3_U5628, P3_U5629, P3_U5630, P3_U5631, P3_U5632, P3_U5633, P3_U5634, P3_U5635, P3_U5636, P3_U5637, P3_U5638, P3_U5639, P3_U5640, P3_U5641, P3_U5642, P3_U5643, P3_U5644, P3_U5645, P3_U5646, P3_U5647, P3_U5648, P3_U5649, P3_U5650, P3_U5651, P3_U5652, P3_U5653, P3_U5654, P3_U5655, P3_U5656, P3_U5657, P3_U5658, P3_U5659, P3_U5660, P3_U5661, P3_U5662, P3_U5663, P3_U5664, P3_U5665, P3_U5666, P3_U5667, P3_U5668, P3_U5669, P3_U5670, P3_U5671, P3_U5672, P3_U5673, P3_U5674, P3_U5675, P3_U5676, P3_U5677, P3_U5678, P3_U5679, P3_U5680, P3_U5681, P3_U5682, P3_U5683, P3_U5684, P3_U5685, P3_U5686, P3_U5687, P3_U5688, P3_U5689, P3_U5690, P3_U5691, P3_U5692, P3_U5693, P3_U5694, P3_U5695, P3_U5696, P3_U5697, P3_U5698, P3_U5699, P3_U5700, P3_U5701, P3_U5702, P3_U5703, P3_U5704, P3_U5705, P3_U5706, P3_U5707, P3_U5708, P3_U5709, P3_U5710, P3_U5711, P3_U5712, P3_U5713, P3_U5714, P3_U5715, P3_U5716, P3_U5717, P3_U5718, P3_U5719, P3_U5720, P3_U5721, P3_U5722, P3_U5723, P3_U5724, P3_U5725, P3_U5726, P3_U5727, P3_U5728, P3_U5729, P3_U5730, P3_U5731, P3_U5732, P3_U5733, P3_U5734, P3_U5735, P3_U5736, P3_U5737, P3_U5738, P3_U5739, P3_U5740, P3_U5741, P3_U5742, P3_U5743, P3_U5744, P3_U5745, P3_U5746, P3_U5747, P3_U5748, P3_U5749, P3_U5750, P3_U5751, P3_U5752, P3_U5753, P3_U5754, P3_U5755, P3_U5756, P3_U5757, P3_U5758, P3_U5759, P3_U5760, P3_U5761, P3_U5762, P3_U5763, P3_U5764, P3_U5765, P3_U5766, P3_U5767, P3_U5768, P3_U5769, P3_U5770, P3_U5771, P3_U5772, P3_U5773, P3_U5774, P3_U5775, P3_U5776, P3_U5777, P3_U5778, P3_U5779, P3_U5780, P3_U5781, P3_U5782, P3_U5783, P3_U5784, P3_U5785, P3_U5786, P3_U5787, P3_U5788, P3_U5789, P3_U5790, P3_U5791, P3_U5792, P3_U5793, P3_U5794, P3_U5795, P3_U5796, P3_U5797, P3_U5798, P3_U5799, P3_U5800, P3_U5801, P3_U5802, P3_U5803, P3_U5804, P3_U5805, P3_U5806, P3_U5807, P3_U5808, P3_U5809, P3_U5810, P3_U5811, P3_U5812, P3_U5813, P3_U5814, P3_U5815, P3_U5816, P3_U5817, P3_U5818, P3_U5819, P3_U5820, P3_U5821, P3_U5822, P3_U5823, P3_U5824, P3_U5825, P3_U5826, P3_U5827, P3_U5828, P3_U5829, P3_U5830, P3_U5831, P3_U5832, P3_U5833, P3_U5834, P3_U5835, P3_U5836, P3_U5837, P3_U5838, P3_U5839, P3_U5840, P3_U5841, P3_U5842, P3_U5843, P3_U5844, P3_U5845, P3_U5846, P3_U5847, P3_U5848, P3_U5849, P3_U5850, P3_U5851, P3_U5852, P3_U5853, P3_U5854, P3_U5855, P3_U5856, P3_U5857, P3_U5858, P3_U5859, P3_U5860, P3_U5861, P3_U5862, P3_U5863, P3_U5864, P3_U5865, P3_U5866, P3_U5867, P3_U5868, P3_U5869, P3_U5870, P3_U5871, P3_U5872, P3_U5873, P3_U5874, P3_U5875, P3_U5876, P3_U5877, P3_U5878, P3_U5879, P3_U5880, P3_U5881, P3_U5882, P3_U5883, P3_U5884, P3_U5885, P3_U5886, P3_U5887, P3_U5888, P3_U5889, P3_U5890, P3_U5891, P3_U5892, P3_U5893, P3_U5894, P3_U5895, P3_U5896, P3_U5897, P3_U5898, P3_U5899, P3_U5900, P3_U5901, P3_U5902, P3_U5903, P3_U5904, P3_U5905, P3_U5906, P3_U5907, P3_U5908, P3_U5909, P3_U5910, P3_U5911, P3_U5912, P3_U5913, P3_U5914, P3_U5915, P3_U5916, P3_U5917, P3_U5918, P3_U5919, P3_U5920, P3_U5921, P3_U5922, P3_U5923, P3_U5924, P3_U5925, P3_U5926, P3_U5927, P3_U5928, P3_U5929, P3_U5930, P3_U5931, P3_U5932, P3_U5933, P3_U5934, P3_U5935, P3_U5936, P3_U5937, P3_U5938, P3_U5939, P3_U5940, P3_U5941, P3_U5942, P3_U5943, P3_U5944, P3_U5945, P3_U5946, P3_U5947, P3_U5948, P3_U5949, P3_U5950, P3_U5951, P3_U5952, P3_U5953, P3_U5954, P3_U5955, P3_U5956, P3_U5957, P3_U5958, P3_U5959, P3_U5960, P3_U5961, P3_U5962, P3_U5963, P3_U5964, P3_U5965, P3_U5966, P3_U5967, P3_U5968, P3_U5969, P3_U5970, P3_U5971, P3_U5972, P3_U5973, P3_U5974, P3_U5975, P3_U5976, P3_U5977, P3_U5978, P3_U5979, P3_U5980, P3_U5981, P3_U5982, P3_U5983, P3_U5984, P3_U5985, P3_U5986, P3_U5987, P3_U5988, P3_U5989, P3_U5990, P3_U5991, P3_U5992, P3_U5993, P3_U5994, P3_U5995, P3_U5996, P3_U5997, P3_U5998, P3_U5999, P3_U6000, P3_U6001, P3_U6002, P3_U6003, P3_U6004, P3_U6005, P3_U6006, P3_U6007, P3_U6008, P3_U6009, P3_U6010, P3_U6011, P3_U6012, P3_U6013, P3_U6014, P3_U6015, P3_U6016, P3_U6017, P3_U6018, P3_U6019, P3_U6020, P3_U6021, P3_U6022, P3_U6023, P3_U6024, P3_U6025, P3_U6026, P3_U6027, P3_U6028, P3_U6029, P3_U6030, P3_U6031, P3_U6032, P3_U6033, P3_U6034, P3_U6035, P3_U6036, P3_U6037, P3_U6038, P3_U6039, P3_U6040, P3_U6041, P3_U6042, P3_U6043, P3_U6044, P3_U6045, P3_U6046, P3_U6047, P3_U6048, P3_U6049, P3_U6050, P3_U6051, P3_U6052, P3_U6053, P3_U6054, P3_U6055, P3_U6056, P3_U6057, P3_U6058, P3_U6059, P3_U6060, P3_U6061, P3_U6062, P3_U6063, P3_U6064, P3_U6065, P3_U6066, P3_U6067, P3_U6068, P3_U6069, P3_U6070, P3_U6071, P3_U6072, P3_U6073, P3_U6074, P3_U6075, P3_U6076, P3_U6077, P3_U6078, P3_U6079, P3_U6080, P3_U6081, P3_U6082, P3_U6083, P3_U6084, P3_U6085, P3_U6086, P3_U6087, P3_U6088, P3_U6089, P3_U6090, P3_U6091, P3_U6092, P3_U6093, P3_U6094, P3_U6095, P3_U6096, P3_U6097, P3_U6098, P3_U6099, P3_U6100, P3_U6101, P3_U6102, P3_U6103, P3_U6104, P3_U6105, P3_U6106, P3_U6107, P3_U6108, P3_U6109, P3_U6110, P3_U6111, P3_U6112, P3_U6113, P3_U6114, P3_U6115, P3_U6116, P3_U6117, P3_U6118, P3_U6119, P3_U6120, P3_U6121, P3_U6122, P3_U6123, P3_U6124, P3_U6125, P3_U6126, P3_U6127, P3_U6128, P3_U6129, P3_U6130, P3_U6131, P3_U6132, P3_U6133, P3_U6134, P3_U6135, P3_U6136, P3_U6137, P3_U6138, P3_U6139, P3_U6140, P3_U6141, P3_U6142, P3_U6143, P3_U6144, P3_U6145, P3_U6146, P3_U6147, P3_U6148, P3_U6149, P3_U6150, P3_U6151, P3_U6152, P3_U6153, P3_U6154, P3_U6155, P3_U6156, P3_U6157, P3_U6158, P3_U6159, P3_U6160, P3_U6161, P3_U6162, P3_U6163, P3_U6164, P3_U6165, P3_U6166, P3_U6167, P3_U6168, P3_U6169, P3_U6170, P3_U6171, P3_U6172, P3_U6173, P3_U6174, P3_U6175, P3_U6176, P3_U6177, P3_U6178, P3_U6179, P3_U6180, P3_U6181, P3_U6182, P3_U6183, P3_U6184, P3_U6185, P3_U6186, P3_U6187, P3_U6188, P3_U6189, P3_U6190, P3_U6191, P3_U6192, P3_U6193, P3_U6194, P3_U6195, P3_U6196, P3_U6197, P3_U6198, P3_U6199, P3_U6200, P3_U6201, P3_U6202, P3_U6203, P3_U6204, P3_U6205, P3_U6206, P3_U6207, P3_U6208, P3_U6209, P3_U6210, P3_U6211, P3_U6212, P3_U6213, P3_U6214, P3_U6215, P3_U6216, P3_U6217, P3_U6218, P3_U6219, P3_U6220, P3_U6221, P3_U6222, P3_U6223, P3_U6224, P3_U6225, P3_U6226, P3_U6227, P3_U6228, P3_U6229, P3_U6230, P3_U6231, P3_U6232, P3_U6233, P3_U6234, P3_U6235, P3_U6236, P3_U6237, P3_U6238, P3_U6239, P3_U6240, P3_U6241, P3_U6242, P3_U6243, P3_U6244, P3_U6245, P3_U6246, P3_U6247, P3_U6248, P3_U6249, P3_U6250, P3_U6251, P3_U6252, P3_U6253, P3_U6254, P3_U6255, P3_U6256, P3_U6257, P3_U6258, P3_U6259, P3_U6260, P3_U6261, P3_U6262, P3_U6263, P3_U6264, P3_U6265, P3_U6266, P3_U6267, P3_U6268, P3_U6269, P3_U6270, P3_U6271, P3_U6272, P3_U6273, P3_U6274, P3_U6275, P3_U6276, P3_U6277, P3_U6278, P3_U6279, P3_U6280, P3_U6281, P3_U6282, P3_U6283, P3_U6284, P3_U6285, P3_U6286, P3_U6287, P3_U6288, P3_U6289, P3_U6290, P3_U6291, P3_U6292, P3_U6293, P3_U6294, P3_U6295, P3_U6296, P3_U6297, P3_U6298, P3_U6299, P3_U6300, P3_U6301, P3_U6302, P3_U6303, P3_U6304, P3_U6305, P3_U6306, P3_U6307, P3_U6308, P3_U6309, P3_U6310, P3_U6311, P3_U6312, P3_U6313, P3_U6314, P3_U6315, P3_U6316, P3_U6317, P3_U6318, P3_U6319, P3_U6320, P3_U6321, P3_U6322, P3_U6323, P3_U6324, P3_U6325, P3_U6326, P3_U6327, P3_U6328, P3_U6329, P3_U6330, P3_U6331, P3_U6332, P3_U6333, P3_U6334, P3_U6335, P3_U6336, P3_U6337, P3_U6338, P3_U6339, P3_U6340, P3_U6341, P3_U6342, P3_U6343, P3_U6344, P3_U6345, P3_U6346, P3_U6347, P3_U6348, P3_U6349, P3_U6350, P3_U6351, P3_U6352, P3_U6353, P3_U6354, P3_U6355, P3_U6356, P3_U6357, P3_U6358, P3_U6359, P3_U6360, P3_U6361, P3_U6362, P3_U6363, P3_U6364, P3_U6365, P3_U6366, P3_U6367, P3_U6368, P3_U6369, P3_U6370, P3_U6371, P3_U6372, P3_U6373, P3_U6374, P3_U6375, P3_U6376, P3_U6377, P3_U6378, P3_U6379, P3_U6380, P3_U6381, P3_U6382, P3_U6383, P3_U6384, P3_U6385, P3_U6386, P3_U6387, P3_U6388, P3_U6389, P3_U6390, P3_U6391, P3_U6392, P3_U6393, P3_U6394, P3_U6395, P3_U6396, P3_U6397, P3_U6398, P3_U6399, P3_U6400, P3_U6401, P3_U6402, P3_U6403, P3_U6404, P3_U6405, P3_U6406, P3_U6407, P3_U6408, P3_U6409, P3_U6410, P3_U6411, P3_U6412, P3_U6413, P3_U6414, P3_U6415, P3_U6416, P3_U6417, P3_U6418, P3_U6419, P3_U6420, P3_U6421, P3_U6422, P3_U6423, P3_U6424, P3_U6425, P3_U6426, P3_U6427, P3_U6428, P3_U6429, P3_U6430, P3_U6431, P3_U6432, P3_U6433, P3_U6434, P3_U6435, P3_U6436, P3_U6437, P3_U6438, P3_U6439, P3_U6440, P3_U6441, P3_U6442, P3_U6443, P3_U6444, P3_U6445, P3_U6446, P3_U6447, P3_U6448, P3_U6449, P3_U6450, P3_U6451, P3_U6452, P3_U6453, P3_U6454, P3_U6455, P3_U6456, P3_U6457, P3_U6458, P3_U6459, P3_U6460, P3_U6461, P3_U6462, P3_U6463, P3_U6464, P3_U6465, P3_U6466, P3_U6467, P3_U6468, P3_U6469, P3_U6470, P3_U6471, P3_U6472, P3_U6473, P3_U6474, P3_U6475, P3_U6476, P3_U6477, P3_U6478, P3_U6479, P3_U6480, P3_U6481, P3_U6482, P3_U6483, P3_U6484, P3_U6485, P3_U6486, P3_U6487, P3_U6488, P3_U6489, P3_U6490, P3_U6491, P3_U6492, P3_U6493, P3_U6494, P3_U6495, P3_U6496, P3_U6497, P3_U6498, P3_U6499, P3_U6500, P3_U6501, P3_U6502, P3_U6503, P3_U6504, P3_U6505, P3_U6506, P3_U6507, P3_U6508, P3_U6509, P3_U6510, P3_U6511, P3_U6512, P3_U6513, P3_U6514, P3_U6515, P3_U6516, P3_U6517, P3_U6518, P3_U6519, P3_U6520, P3_U6521, P3_U6522, P3_U6523, P3_U6524, P3_U6525, P3_U6526, P3_U6527, P3_U6528, P3_U6529, P3_U6530, P3_U6531, P3_U6532, P3_U6533, P3_U6534, P3_U6535, P3_U6536, P3_U6537, P3_U6538, P3_U6539, P3_U6540, P3_U6541, P3_U6542, P3_U6543, P3_U6544, P3_U6545, P3_U6546, P3_U6547, P3_U6548, P3_U6549, P3_U6550, P3_U6551, P3_U6552, P3_U6553, P3_U6554, P3_U6555, P3_U6556, P3_U6557, P3_U6558, P3_U6559, P3_U6560, P3_U6561, P3_U6562, P3_U6563, P3_U6564, P3_U6565, P3_U6566, P3_U6567, P3_U6568, P3_U6569, P3_U6570, P3_U6571, P3_U6572, P3_U6573, P3_U6574, P3_U6575, P3_U6576, P3_U6577, P3_U6578, P3_U6579, P3_U6580, P3_U6581, P3_U6582, P3_U6583, P3_U6584, P3_U6585, P3_U6586, P3_U6587, P3_U6588, P3_U6589, P3_U6590, P3_U6591, P3_U6592, P3_U6593, P3_U6594, P3_U6595, P3_U6596, P3_U6597, P3_U6598, P3_U6599, P3_U6600, P3_U6601, P3_U6602, P3_U6603, P3_U6604, P3_U6605, P3_U6606, P3_U6607, P3_U6608, P3_U6609, P3_U6610, P3_U6611, P3_U6612, P3_U6613, P3_U6614, P3_U6615, P3_U6616, P3_U6617, P3_U6618, P3_U6619, P3_U6620, P3_U6621, P3_U6622, P3_U6623, P3_U6624, P3_U6625, P3_U6626, P3_U6627, P3_U6628, P3_U6629, P3_U6630, P3_U6631, P3_U6632, P3_U6633, P3_U6634, P3_U6635, P3_U6636, P3_U6637, P3_U6638, P3_U6639, P3_U6640, P3_U6641, P3_U6642, P3_U6643, P3_U6644, P3_U6645, P3_U6646, P3_U6647, P3_U6648, P3_U6649, P3_U6650, P3_U6651, P3_U6652, P3_U6653, P3_U6654, P3_U6655, P3_U6656, P3_U6657, P3_U6658, P3_U6659, P3_U6660, P3_U6661, P3_U6662, P3_U6663, P3_U6664, P3_U6665, P3_U6666, P3_U6667, P3_U6668, P3_U6669, P3_U6670, P3_U6671, P3_U6672, P3_U6673, P3_U6674, P3_U6675, P3_U6676, P3_U6677, P3_U6678, P3_U6679, P3_U6680, P3_U6681, P3_U6682, P3_U6683, P3_U6684, P3_U6685, P3_U6686, P3_U6687, P3_U6688, P3_U6689, P3_U6690, P3_U6691, P3_U6692, P3_U6693, P3_U6694, P3_U6695, P3_U6696, P3_U6697, P3_U6698, P3_U6699, P3_U6700, P3_U6701, P3_U6702, P3_U6703, P3_U6704, P3_U6705, P3_U6706, P3_U6707, P3_U6708, P3_U6709, P3_U6710, P3_U6711, P3_U6712, P3_U6713, P3_U6714, P3_U6715, P3_U6716, P3_U6717, P3_U6718, P3_U6719, P3_U6720, P3_U6721, P3_U6722, P3_U6723, P3_U6724, P3_U6725, P3_U6726, P3_U6727, P3_U6728, P3_U6729, P3_U6730, P3_U6731, P3_U6732, P3_U6733, P3_U6734, P3_U6735, P3_U6736, P3_U6737, P3_U6738, P3_U6739, P3_U6740, P3_U6741, P3_U6742, P3_U6743, P3_U6744, P3_U6745, P3_U6746, P3_U6747, P3_U6748, P3_U6749, P3_U6750, P3_U6751, P3_U6752, P3_U6753, P3_U6754, P3_U6755, P3_U6756, P3_U6757, P3_U6758, P3_U6759, P3_U6760, P3_U6761, P3_U6762, P3_U6763, P3_U6764, P3_U6765, P3_U6766, P3_U6767, P3_U6768, P3_U6769, P3_U6770, P3_U6771, P3_U6772, P3_U6773, P3_U6774, P3_U6775, P3_U6776, P3_U6777, P3_U6778, P3_U6779, P3_U6780, P3_U6781, P3_U6782, P3_U6783, P3_U6784, P3_U6785, P3_U6786, P3_U6787, P3_U6788, P3_U6789, P3_U6790, P3_U6791, P3_U6792, P3_U6793, P3_U6794, P3_U6795, P3_U6796, P3_U6797, P3_U6798, P3_U6799, P3_U6800, P3_U6801, P3_U6802, P3_U6803, P3_U6804, P3_U6805, P3_U6806, P3_U6807, P3_U6808, P3_U6809, P3_U6810, P3_U6811, P3_U6812, P3_U6813, P3_U6814, P3_U6815, P3_U6816, P3_U6817, P3_U6818, P3_U6819, P3_U6820, P3_U6821, P3_U6822, P3_U6823, P3_U6824, P3_U6825, P3_U6826, P3_U6827, P3_U6828, P3_U6829, P3_U6830, P3_U6831, P3_U6832, P3_U6833, P3_U6834, P3_U6835, P3_U6836, P3_U6837, P3_U6838, P3_U6839, P3_U6840, P3_U6841, P3_U6842, P3_U6843, P3_U6844, P3_U6845, P3_U6846, P3_U6847, P3_U6848, P3_U6849, P3_U6850, P3_U6851, P3_U6852, P3_U6853, P3_U6854, P3_U6855, P3_U6856, P3_U6857, P3_U6858, P3_U6859, P3_U6860, P3_U6861, P3_U6862, P3_U6863, P3_U6864, P3_U6865, P3_U6866, P3_U6867, P3_U6868, P3_U6869, P3_U6870, P3_U6871, P3_U6872, P3_U6873, P3_U6874, P3_U6875, P3_U6876, P3_U6877, P3_U6878, P3_U6879, P3_U6880, P3_U6881, P3_U6882, P3_U6883, P3_U6884, P3_U6885, P3_U6886, P3_U6887, P3_U6888, P3_U6889, P3_U6890, P3_U6891, P3_U6892, P3_U6893, P3_U6894, P3_U6895, P3_U6896, P3_U6897, P3_U6898, P3_U6899, P3_U6900, P3_U6901, P3_U6902, P3_U6903, P3_U6904, P3_U6905, P3_U6906, P3_U6907, P3_U6908, P3_U6909, P3_U6910, P3_U6911, P3_U6912, P3_U6913, P3_U6914, P3_U6915, P3_U6916, P3_U6917, P3_U6918, P3_U6919, P3_U6920, P3_U6921, P3_U6922, P3_U6923, P3_U6924, P3_U6925, P3_U6926, P3_U6927, P3_U6928, P3_U6929, P3_U6930, P3_U6931, P3_U6932, P3_U6933, P3_U6934, P3_U6935, P3_U6936, P3_U6937, P3_U6938, P3_U6939, P3_U6940, P3_U6941, P3_U6942, P3_U6943, P3_U6944, P3_U6945, P3_U6946, P3_U6947, P3_U6948, P3_U6949, P3_U6950, P3_U6951, P3_U6952, P3_U6953, P3_U6954, P3_U6955, P3_U6956, P3_U6957, P3_U6958, P3_U6959, P3_U6960, P3_U6961, P3_U6962, P3_U6963, P3_U6964, P3_U6965, P3_U6966, P3_U6967, P3_U6968, P3_U6969, P3_U6970, P3_U6971, P3_U6972, P3_U6973, P3_U6974, P3_U6975, P3_U6976, P3_U6977, P3_U6978, P3_U6979, P3_U6980, P3_U6981, P3_U6982, P3_U6983, P3_U6984, P3_U6985, P3_U6986, P3_U6987, P3_U6988, P3_U6989, P3_U6990, P3_U6991, P3_U6992, P3_U6993, P3_U6994, P3_U6995, P3_U6996, P3_U6997, P3_U6998, P3_U6999, P3_U7000, P3_U7001, P3_U7002, P3_U7003, P3_U7004, P3_U7005, P3_U7006, P3_U7007, P3_U7008, P3_U7009, P3_U7010, P3_U7011, P3_U7012, P3_U7013, P3_U7014, P3_U7015, P3_U7016, P3_U7017, P3_U7018, P3_U7019, P3_U7020, P3_U7021, P3_U7022, P3_U7023, P3_U7024, P3_U7025, P3_U7026, P3_U7027, P3_U7028, P3_U7029, P3_U7030, P3_U7031, P3_U7032, P3_U7033, P3_U7034, P3_U7035, P3_U7036, P3_U7037, P3_U7038, P3_U7039, P3_U7040, P3_U7041, P3_U7042, P3_U7043, P3_U7044, P3_U7045, P3_U7046, P3_U7047, P3_U7048, P3_U7049, P3_U7050, P3_U7051, P3_U7052, P3_U7053, P3_U7054, P3_U7055, P3_U7056, P3_U7057, P3_U7058, P3_U7059, P3_U7060, P3_U7061, P3_U7062, P3_U7063, P3_U7064, P3_U7065, P3_U7066, P3_U7067, P3_U7068, P3_U7069, P3_U7070, P3_U7071, P3_U7072, P3_U7073, P3_U7074, P3_U7075, P3_U7076, P3_U7077, P3_U7078, P3_U7079, P3_U7080, P3_U7081, P3_U7082, P3_U7083, P3_U7084, P3_U7085, P3_U7086, P3_U7087, P3_U7088, P3_U7089, P3_U7090, P3_U7091, P3_U7092, P3_U7093, P3_U7094, P3_U7095, P3_U7096, P3_U7097, P3_U7098, P3_U7099, P3_U7100, P3_U7101, P3_U7102, P3_U7103, P3_U7104, P3_U7105, P3_U7106, P3_U7107, P3_U7108, P3_U7109, P3_U7110, P3_U7111, P3_U7112, P3_U7113, P3_U7114, P3_U7115, P3_U7116, P3_U7117, P3_U7118, P3_U7119, P3_U7120, P3_U7121, P3_U7122, P3_U7123, P3_U7124, P3_U7125, P3_U7126, P3_U7127, P3_U7128, P3_U7129, P3_U7130, P3_U7131, P3_U7132, P3_U7133, P3_U7134, P3_U7135, P3_U7136, P3_U7137, P3_U7138, P3_U7139, P3_U7140, P3_U7141, P3_U7142, P3_U7143, P3_U7144, P3_U7145, P3_U7146, P3_U7147, P3_U7148, P3_U7149, P3_U7150, P3_U7151, P3_U7152, P3_U7153, P3_U7154, P3_U7155, P3_U7156, P3_U7157, P3_U7158, P3_U7159, P3_U7160, P3_U7161, P3_U7162, P3_U7163, P3_U7164, P3_U7165, P3_U7166, P3_U7167, P3_U7168, P3_U7169, P3_U7170, P3_U7171, P3_U7172, P3_U7173, P3_U7174, P3_U7175, P3_U7176, P3_U7177, P3_U7178, P3_U7179, P3_U7180, P3_U7181, P3_U7182, P3_U7183, P3_U7184, P3_U7185, P3_U7186, P3_U7187, P3_U7188, P3_U7189, P3_U7190, P3_U7191, P3_U7192, P3_U7193, P3_U7194, P3_U7195, P3_U7196, P3_U7197, P3_U7198, P3_U7199, P3_U7200, P3_U7201, P3_U7202, P3_U7203, P3_U7204, P3_U7205, P3_U7206, P3_U7207, P3_U7208, P3_U7209, P3_U7210, P3_U7211, P3_U7212, P3_U7213, P3_U7214, P3_U7215, P3_U7216, P3_U7217, P3_U7218, P3_U7219, P3_U7220, P3_U7221, P3_U7222, P3_U7223, P3_U7224, P3_U7225, P3_U7226, P3_U7227, P3_U7228, P3_U7229, P3_U7230, P3_U7231, P3_U7232, P3_U7233, P3_U7234, P3_U7235, P3_U7236, P3_U7237, P3_U7238, P3_U7239, P3_U7240, P3_U7241, P3_U7242, P3_U7243, P3_U7244, P3_U7245, P3_U7246, P3_U7247, P3_U7248, P3_U7249, P3_U7250, P3_U7251, P3_U7252, P3_U7253, P3_U7254, P3_U7255, P3_U7256, P3_U7257, P3_U7258, P3_U7259, P3_U7260, P3_U7261, P3_U7262, P3_U7263, P3_U7264, P3_U7265, P3_U7266, P3_U7267, P3_U7268, P3_U7269, P3_U7270, P3_U7271, P3_U7272, P3_U7273, P3_U7274, P3_U7275, P3_U7276, P3_U7277, P3_U7278, P3_U7279, P3_U7280, P3_U7281, P3_U7282, P3_U7283, P3_U7284, P3_U7285, P3_U7286, P3_U7287, P3_U7288, P3_U7289, P3_U7290, P3_U7291, P3_U7292, P3_U7293, P3_U7294, P3_U7295, P3_U7296, P3_U7297, P3_U7298, P3_U7299, P3_U7300, P3_U7301, P3_U7302, P3_U7303, P3_U7304, P3_U7305, P3_U7306, P3_U7307, P3_U7308, P3_U7309, P3_U7310, P3_U7311, P3_U7312, P3_U7313, P3_U7314, P3_U7315, P3_U7316, P3_U7317, P3_U7318, P3_U7319, P3_U7320, P3_U7321, P3_U7322, P3_U7323, P3_U7324, P3_U7325, P3_U7326, P3_U7327, P3_U7328, P3_U7329, P3_U7330, P3_U7331, P3_U7332, P3_U7333, P3_U7334, P3_U7335, P3_U7336, P3_U7337, P3_U7338, P3_U7339, P3_U7340, P3_U7341, P3_U7342, P3_U7343, P3_U7344, P3_U7345, P3_U7346, P3_U7347, P3_U7348, P3_U7349, P3_U7350, P3_U7351, P3_U7352, P3_U7353, P3_U7354, P3_U7355, P3_U7356, P3_U7357, P3_U7358, P3_U7359, P3_U7360, P3_U7361, P3_U7362, P3_U7363, P3_U7364, P3_U7365, P3_U7366, P3_U7367, P3_U7368, P3_U7369, P3_U7370, P3_U7371, P3_U7372, P3_U7373, P3_U7374, P3_U7375, P3_U7376, P3_U7377, P3_U7378, P3_U7379, P3_U7380, P3_U7381, P3_U7382, P3_U7383, P3_U7384, P3_U7385, P3_U7386, P3_U7387, P3_U7388, P3_U7389, P3_U7390, P3_U7391, P3_U7392, P3_U7393, P3_U7394, P3_U7395, P3_U7396, P3_U7397, P3_U7398, P3_U7399, P3_U7400, P3_U7401, P3_U7402, P3_U7403, P3_U7404, P3_U7405, P3_U7406, P3_U7407, P3_U7408, P3_U7409, P3_U7410, P3_U7411, P3_U7412, P3_U7413, P3_U7414, P3_U7415, P3_U7416, P3_U7417, P3_U7418, P3_U7419, P3_U7420, P3_U7421, P3_U7422, P3_U7423, P3_U7424, P3_U7425, P3_U7426, P3_U7427, P3_U7428, P3_U7429, P3_U7430, P3_U7431, P3_U7432, P3_U7433, P3_U7434, P3_U7435, P3_U7436, P3_U7437, P3_U7438, P3_U7439, P3_U7440, P3_U7441, P3_U7442, P3_U7443, P3_U7444, P3_U7445, P3_U7446, P3_U7447, P3_U7448, P3_U7449, P3_U7450, P3_U7451, P3_U7452, P3_U7453, P3_U7454, P3_U7455, P3_U7456, P3_U7457, P3_U7458, P3_U7459, P3_U7460, P3_U7461, P3_U7462, P3_U7463, P3_U7464, P3_U7465, P3_U7466, P3_U7467, P3_U7468, P3_U7469, P3_U7470, P3_U7471, P3_U7472, P3_U7473, P3_U7474, P3_U7475, P3_U7476, P3_U7477, P3_U7478, P3_U7479, P3_U7480, P3_U7481, P3_U7482, P3_U7483, P3_U7484, P3_U7485, P3_U7486, P3_U7487, P3_U7488, P3_U7489, P3_U7490, P3_U7491, P3_U7492, P3_U7493, P3_U7494, P3_U7495, P3_U7496, P3_U7497, P3_U7498, P3_U7499, P3_U7500, P3_U7501, P3_U7502, P3_U7503, P3_U7504, P3_U7505, P3_U7506, P3_U7507, P3_U7508, P3_U7509, P3_U7510, P3_U7511, P3_U7512, P3_U7513, P3_U7514, P3_U7515, P3_U7516, P3_U7517, P3_U7518, P3_U7519, P3_U7520, P3_U7521, P3_U7522, P3_U7523, P3_U7524, P3_U7525, P3_U7526, P3_U7527, P3_U7528, P3_U7529, P3_U7530, P3_U7531, P3_U7532, P3_U7533, P3_U7534, P3_U7535, P3_U7536, P3_U7537, P3_U7538, P3_U7539, P3_U7540, P3_U7541, P3_U7542, P3_U7543, P3_U7544, P3_U7545, P3_U7546, P3_U7547, P3_U7548, P3_U7549, P3_U7550, P3_U7551, P3_U7552, P3_U7553, P3_U7554, P3_U7555, P3_U7556, P3_U7557, P3_U7558, P3_U7559, P3_U7560, P3_U7561, P3_U7562, P3_U7563, P3_U7564, P3_U7565, P3_U7566, P3_U7567, P3_U7568, P3_U7569, P3_U7570, P3_U7571, P3_U7572, P3_U7573, P3_U7574, P3_U7575, P3_U7576, P3_U7577, P3_U7578, P3_U7579, P3_U7580, P3_U7581, P3_U7582, P3_U7583, P3_U7584, P3_U7585, P3_U7586, P3_U7587, P3_U7588, P3_U7589, P3_U7590, P3_U7591, P3_U7592, P3_U7593, P3_U7594, P3_U7595, P3_U7596, P3_U7597, P3_U7598, P3_U7599, P3_U7600, P3_U7601, P3_U7602, P3_U7603, P3_U7604, P3_U7605, P3_U7606, P3_U7607, P3_U7608, P3_U7609, P3_U7610, P3_U7611, P3_U7612, P3_U7613, P3_U7614, P3_U7615, P3_U7616, P3_U7617, P3_U7618, P3_U7619, P3_U7620, P3_U7621, P3_U7622, P3_U7623, P3_U7624, P3_U7625, P3_U7626, P3_U7627, P3_U7628, P3_U7629, P3_U7630, P3_U7631, P3_U7632, P3_U7633, P3_U7634, P3_U7635, P3_U7636, P3_U7637, P3_U7638, P3_U7639, P3_U7640, P3_U7641, P3_U7642, P3_U7643, P3_U7644, P3_U7645, P3_U7646, P3_U7647, P3_U7648, P3_U7649, P3_U7650, P3_U7651, P3_U7652, P3_U7653, P3_U7654, P3_U7655, P3_U7656, P3_U7657, P3_U7658, P3_U7659, P3_U7660, P3_U7661, P3_U7662, P3_U7663, P3_U7664, P3_U7665, P3_U7666, P3_U7667, P3_U7668, P3_U7669, P3_U7670, P3_U7671, P3_U7672, P3_U7673, P3_U7674, P3_U7675, P3_U7676, P3_U7677, P3_U7678, P3_U7679, P3_U7680, P3_U7681, P3_U7682, P3_U7683, P3_U7684, P3_U7685, P3_U7686, P3_U7687, P3_U7688, P3_U7689, P3_U7690, P3_U7691, P3_U7692, P3_U7693, P3_U7694, P3_U7695, P3_U7696, P3_U7697, P3_U7698, P3_U7699, P3_U7700, P3_U7701, P3_U7702, P3_U7703, P3_U7704, P3_U7705, P3_U7706, P3_U7707, P3_U7708, P3_U7709, P3_U7710, P3_U7711, P3_U7712, P3_U7713, P3_U7714, P3_U7715, P3_U7716, P3_U7717, P3_U7718, P3_U7719, P3_U7720, P3_U7721, P3_U7722, P3_U7723, P3_U7724, P3_U7725, P3_U7726, P3_U7727, P3_U7728, P3_U7729, P3_U7730, P3_U7731, P3_U7732, P3_U7733, P3_U7734, P3_U7735, P3_U7736, P3_U7737, P3_U7738, P3_U7739, P3_U7740, P3_U7741, P3_U7742, P3_U7743, P3_U7744, P3_U7745, P3_U7746, P3_U7747, P3_U7748, P3_U7749, P3_U7750, P3_U7751, P3_U7752, P3_U7753, P3_U7754, P3_U7755, P3_U7756, P3_U7757, P3_U7758, P3_U7759, P3_U7760, P3_U7761, P3_U7762, P3_U7763, P3_U7764, P3_U7765, P3_U7766, P3_U7767, P3_U7768, P3_U7769, P3_U7770, P3_U7771, P3_U7772, P3_U7773, P3_U7774, P3_U7775, P3_U7776, P3_U7777, P3_U7778, P3_U7779, P3_U7780, P3_U7781, P3_U7782, P3_U7783, P3_U7784, P3_U7785, P3_U7786, P3_U7787, P3_U7788, P3_U7789, P3_U7790, P3_U7791, P3_U7792, P3_U7793, P3_U7794, P3_U7795, P3_U7796, P3_U7797, P3_U7798, P3_U7799, P3_U7800, P3_U7801, P3_U7802, P3_U7803, P3_U7804, P3_U7805, P3_U7806, P3_U7807, P3_U7808, P3_U7809, P3_U7810, P3_U7811, P3_U7812, P3_U7813, P3_U7814, P3_U7815, P3_U7816, P3_U7817, P3_U7818, P3_U7819, P3_U7820, P3_U7821, P3_U7822, P3_U7823, P3_U7824, P3_U7825, P3_U7826, P3_U7827, P3_U7828, P3_U7829, P3_U7830, P3_U7831, P3_U7832, P3_U7833, P3_U7834, P3_U7835, P3_U7836, P3_U7837, P3_U7838, P3_U7839, P3_U7840, P3_U7841, P3_U7842, P3_U7843, P3_U7844, P3_U7845, P3_U7846, P3_U7847, P3_U7848, P3_U7849, P3_U7850, P3_U7851, P3_U7852, P3_U7853, P3_U7854, P3_U7855, P3_U7856, P3_U7857, P3_U7858, P3_U7859, P3_U7860, P3_U7861, P3_U7862, P3_U7863, P3_U7864, P3_U7865, P3_U7866, P3_U7867, P3_U7868, P3_U7869, P3_U7870, P3_U7871, P3_U7872, P3_U7873, P3_U7874, P3_U7875, P3_U7876, P3_U7877, P3_U7878, P3_U7879, P3_U7880, P3_U7881, P3_U7882, P3_U7883, P3_U7884, P3_U7885, P3_U7886, P3_U7887, P3_U7888, P3_U7889, P3_U7890, P3_U7891, P3_U7892, P3_U7893, P3_U7894, P3_U7895, P3_U7896, P3_U7897, P3_U7898, P3_U7899, P3_U7900, P3_U7901, P3_U7902, P3_U7903, P3_U7904, P3_U7905, P3_U7906, P3_U7907, P3_U7908, P3_U7909, P3_U7910, P3_U7911, P3_U7912, P3_U7913, P3_U7914, P3_U7915, P3_U7916, P3_U7917, P3_U7918, P3_U7919, P3_U7920, P3_U7921, P3_U7922, P3_U7923, P3_U7924, P3_U7925, P3_U7926, P3_U7927, P3_U7928, P3_U7929, P3_U7930, P3_U7931, P3_U7932, P3_U7933, P3_U7934, P3_U7935, P3_U7936, P3_U7937, P3_U7938, P3_U7939, P3_U7940, P3_U7941, P3_U7942, P3_U7943, P3_U7944, P3_U7945, P3_U7946, P3_U7947, P3_U7948, P3_U7949, P3_U7950, P3_U7951, P3_U7952, P3_U7953, P3_U7954, P3_U7955, P3_U7956, P3_U7957, P3_U7958, P3_U7959, P3_U7960, P3_U7961, P3_U7962, P3_U7963, P3_U7964, P3_U7965, P3_U7966, P3_U7967, P3_U7968, P3_U7969, P3_U7970, P3_U7971, P3_U7972, P3_U7973, P3_U7974, P3_U7975, P3_U7976, P3_U7977, P3_U7978, P3_U7979, P3_U7980, P3_U7981, P3_U7982, P3_U7983, P3_U7984, P3_U7985, P3_U7986, P3_U7987, P3_U7988, P3_U7989, P3_U7990, P3_U7991, P3_U7992, P3_U7993, P3_U7994, P3_U7995, P3_U7996, P3_U7997, P3_U7998, P3_U7999, P3_U8000, P3_U8001, P3_U8002, P3_U8003, P3_U8004, P3_U8005, P3_U8006, P3_U8007, P3_U8008, P3_U8009, P3_U8010, P3_U8011, P3_U8012, P3_U8013, P3_U8014, P3_U8015, P3_U8016, P3_U8017, P3_U8018, P3_U8019, P3_U8020, P3_U8021, P3_U8022, P3_U8023, P3_U8024, P3_U8025, P3_U8026, P3_U8027, P3_U8028, P3_U8029, P3_U8030, P3_U8031, P3_U8032, P3_U8033, P3_U8034, P3_U8035, P3_U8036, P3_U8037, P3_U8038, P3_U8039, P3_U8040, P3_U8041, P3_U8042, P3_U8043, P3_U8044, P3_U8045, P3_U8046, P3_U8047, P3_U8048, P3_U8049, P3_U8050, P3_U8051, P3_U8052, P3_U8053, P2_U2352, P2_U2353, P2_U2354, P2_U2355, P2_U2356, P2_U2357, P2_U2358, P2_U2359, P2_U2360, P2_U2361, P2_U2362, P2_U2363, P2_U2364, P2_U2365, P2_U2366, P2_U2367, P2_U2368, P2_U2369, P2_U2370, P2_U2371, P2_U2372, P2_U2373, P2_U2374, P2_U2375, P2_U2376, P2_U2377, P2_U2378, P2_U2379, P2_U2380, P2_U2381, P2_U2382, P2_U2383, P2_U2384, P2_U2385, P2_U2386, P2_U2387, P2_U2388, P2_U2389, P2_U2390, P2_U2391, P2_U2392, P2_U2393, P2_U2394, P2_U2395, P2_U2396, P2_U2397, P2_U2398, P2_U2399, P2_U2400, P2_U2401, P2_U2402, P2_U2403, P2_U2404, P2_U2405, P2_U2406, P2_U2407, P2_U2408, P2_U2409, P2_U2410, P2_U2411, P2_U2412, P2_U2413, P2_U2414, P2_U2415, P2_U2416, P2_U2417, P2_U2418, P2_U2419, P2_U2420, P2_U2421, P2_U2422, P2_U2423, P2_U2424, P2_U2425, P2_U2426, P2_U2427, P2_U2428, P2_U2429, P2_U2430, P2_U2431, P2_U2432, P2_U2433, P2_U2434, P2_U2435, P2_U2436, P2_U2437, P2_U2438, P2_U2439, P2_U2440, P2_U2441, P2_U2442, P2_U2443, P2_U2444, P2_U2445, P2_U2446, P2_U2447, P2_U2448, P2_U2449, P2_U2450, P2_U2451, P2_U2452, P2_U2453, P2_U2454, P2_U2455, P2_U2456, P2_U2457, P2_U2458, P2_U2459, P2_U2460, P2_U2461, P2_U2462, P2_U2463, P2_U2464, P2_U2465, P2_U2466, P2_U2467, P2_U2468, P2_U2469, P2_U2470, P2_U2471, P2_U2472, P2_U2473, P2_U2474, P2_U2475, P2_U2476, P2_U2477, P2_U2478, P2_U2479, P2_U2480, P2_U2481, P2_U2482, P2_U2483, P2_U2484, P2_U2485, P2_U2486, P2_U2487, P2_U2488, P2_U2489, P2_U2490, P2_U2491, P2_U2492, P2_U2493, P2_U2494, P2_U2495, P2_U2496, P2_U2497, P2_U2498, P2_U2499, P2_U2500, P2_U2501, P2_U2502, P2_U2503, P2_U2504, P2_U2505, P2_U2506, P2_U2507, P2_U2508, P2_U2509, P2_U2510, P2_U2511, P2_U2512, P2_U2513, P2_U2514, P2_U2515, P2_U2516, P2_U2517, P2_U2518, P2_U2519, P2_U2520, P2_U2521, P2_U2522, P2_U2523, P2_U2524, P2_U2525, P2_U2526, P2_U2527, P2_U2528, P2_U2529, P2_U2530, P2_U2531, P2_U2532, P2_U2533, P2_U2534, P2_U2535, P2_U2536, P2_U2537, P2_U2538, P2_U2539, P2_U2540, P2_U2541, P2_U2542, P2_U2543, P2_U2544, P2_U2545, P2_U2546, P2_U2547, P2_U2548, P2_U2549, P2_U2550, P2_U2551, P2_U2552, P2_U2553, P2_U2554, P2_U2555, P2_U2556, P2_U2557, P2_U2558, P2_U2559, P2_U2560, P2_U2561, P2_U2562, P2_U2563, P2_U2564, P2_U2565, P2_U2566, P2_U2567, P2_U2568, P2_U2569, P2_U2570, P2_U2571, P2_U2572, P2_U2573, P2_U2574, P2_U2575, P2_U2576, P2_U2577, P2_U2578, P2_U2579, P2_U2580, P2_U2581, P2_U2582, P2_U2583, P2_U2584, P2_U2585, P2_U2586, P2_U2587, P2_U2588, P2_U2589, P2_U2590, P2_U2591, P2_U2592, P2_U2593, P2_U2594, P2_U2595, P2_U2596, P2_U2597, P2_U2598, P2_U2599, P2_U2600, P2_U2601, P2_U2602, P2_U2603, P2_U2604, P2_U2605, P2_U2606, P2_U2607, P2_U2608, P2_U2609, P2_U2610, P2_U2611, P2_U2612, P2_U2613, P2_U2614, P2_U2615, P2_U2616, P2_U2617, P2_U2618, P2_U2619, P2_U2620, P2_U2621, P2_U2622, P2_U2623, P2_U2624, P2_U2625, P2_U2626, P2_U2627, P2_U2628, P2_U2629, P2_U2630, P2_U2631, P2_U2632, P2_U2633, P2_U2634, P2_U2635, P2_U2636, P2_U2637, P2_U2638, P2_U2639, P2_U2640, P2_U2641, P2_U2642, P2_U2643, P2_U2644, P2_U2645, P2_U2646, P2_U2647, P2_U2648, P2_U2649, P2_U2650, P2_U2651, P2_U2652, P2_U2653, P2_U2654, P2_U2655, P2_U2656, P2_U2657, P2_U2658, P2_U2659, P2_U2660, P2_U2661, P2_U2662, P2_U2663, P2_U2664, P2_U2665, P2_U2666, P2_U2667, P2_U2668, P2_U2669, P2_U2670, P2_U2671, P2_U2672, P2_U2673, P2_U2674, P2_U2675, P2_U2676, P2_U2677, P2_U2678, P2_U2679, P2_U2680, P2_U2681, P2_U2682, P2_U2683, P2_U2684, P2_U2685, P2_U2686, P2_U2687, P2_U2688, P2_U2689, P2_U2690, P2_U2691, P2_U2692, P2_U2693, P2_U2694, P2_U2695, P2_U2696, P2_U2698, P2_U2699, P2_U2700, P2_U2701, P2_U2702, P2_U2703, P2_U2704, P2_U2705, P2_U2706, P2_U2707, P2_U2708, P2_U2709, P2_U2710, P2_U2711, P2_U2712, P2_U2713, P2_U2714, P2_U2715, P2_U2716, P2_U2717, P2_U2718, P2_U2719, P2_U2720, P2_U2721, P2_U2722, P2_U2723, P2_U2724, P2_U2725, P2_U2726, P2_U2727, P2_U2728, P2_U2729, P2_U2730, P2_U2731, P2_U2732, P2_U2733, P2_U2734, P2_U2735, P2_U2736, P2_U2737, P2_U2738, P2_U2739, P2_U2740, P2_U2741, P2_U2742, P2_U2743, P2_U2744, P2_U2745, P2_U2746, P2_U2747, P2_U2748, P2_U2749, P2_U2750, P2_U2751, P2_U2752, P2_U2753, P2_U2754, P2_U2755, P2_U2756, P2_U2757, P2_U2758, P2_U2759, P2_U2760, P2_U2761, P2_U2762, P2_U2763, P2_U2764, P2_U2765, P2_U2766, P2_U2767, P2_U2768, P2_U2769, P2_U2770, P2_U2771, P2_U2772, P2_U2773, P2_U2774, P2_U2775, P2_U2776, P2_U2777, P2_U2778, P2_U2779, P2_U2780, P2_U2781, P2_U2782, P2_U2783, P2_U2784, P2_U2785, P2_U2786, P2_U2787, P2_U2788, P2_U2789, P2_U2790, P2_U2791, P2_U2792, P2_U2793, P2_U2794, P2_U2795, P2_U2796, P2_U2797, P2_U2798, P2_U2799, P2_U2800, P2_U2801, P2_U2802, P2_U2803, P2_U2804, P2_U2805, P2_U2806, P2_U2807, P2_U2808, P2_U2809, P2_U2810, P2_U2811, P2_U2812, P2_U2813, P2_U3242, P2_U3243, P2_U3244, P2_U3245, P2_U3246, P2_U3247, P2_U3248, P2_U3249, P2_U3250, P2_U3251, P2_U3252, P2_U3253, P2_U3254, P2_U3255, P2_U3256, P2_U3257, P2_U3258, P2_U3259, P2_U3260, P2_U3261, P2_U3262, P2_U3263, P2_U3264, P2_U3265, P2_U3266, P2_U3267, P2_U3268, P2_U3269, P2_U3270, P2_U3271, P2_U3272, P2_U3273, P2_U3274, P2_U3275, P2_U3276, P2_U3277, P2_U3278, P2_U3279, P2_U3280, P2_U3281, P2_U3282, P2_U3283, P2_U3284, P2_U3285, P2_U3286, P2_U3287, P2_U3288, P2_U3289, P2_U3290, P2_U3291, P2_U3292, P2_U3293, P2_U3294, P2_U3295, P2_U3296, P2_U3297, P2_U3298, P2_U3299, P2_U3300, P2_U3301, P2_U3302, P2_U3303, P2_U3304, P2_U3305, P2_U3306, P2_U3307, P2_U3308, P2_U3309, P2_U3310, P2_U3311, P2_U3312, P2_U3313, P2_U3314, P2_U3315, P2_U3316, P2_U3317, P2_U3318, P2_U3319, P2_U3320, P2_U3321, P2_U3322, P2_U3323, P2_U3324, P2_U3325, P2_U3326, P2_U3327, P2_U3328, P2_U3329, P2_U3330, P2_U3331, P2_U3332, P2_U3333, P2_U3334, P2_U3335, P2_U3336, P2_U3337, P2_U3338, P2_U3339, P2_U3340, P2_U3341, P2_U3342, P2_U3343, P2_U3344, P2_U3345, P2_U3346, P2_U3347, P2_U3348, P2_U3349, P2_U3350, P2_U3351, P2_U3352, P2_U3353, P2_U3354, P2_U3355, P2_U3356, P2_U3357, P2_U3358, P2_U3359, P2_U3360, P2_U3361, P2_U3362, P2_U3363, P2_U3364, P2_U3365, P2_U3366, P2_U3367, P2_U3368, P2_U3369, P2_U3370, P2_U3371, P2_U3372, P2_U3373, P2_U3374, P2_U3375, P2_U3376, P2_U3377, P2_U3378, P2_U3379, P2_U3380, P2_U3381, P2_U3382, P2_U3383, P2_U3384, P2_U3385, P2_U3386, P2_U3387, P2_U3388, P2_U3389, P2_U3390, P2_U3391, P2_U3392, P2_U3393, P2_U3394, P2_U3395, P2_U3396, P2_U3397, P2_U3398, P2_U3399, P2_U3400, P2_U3401, P2_U3402, P2_U3403, P2_U3404, P2_U3405, P2_U3406, P2_U3407, P2_U3408, P2_U3409, P2_U3410, P2_U3411, P2_U3412, P2_U3413, P2_U3414, P2_U3415, P2_U3416, P2_U3417, P2_U3418, P2_U3419, P2_U3420, P2_U3421, P2_U3422, P2_U3423, P2_U3424, P2_U3425, P2_U3426, P2_U3427, P2_U3428, P2_U3429, P2_U3430, P2_U3431, P2_U3432, P2_U3433, P2_U3434, P2_U3435, P2_U3436, P2_U3437, P2_U3438, P2_U3439, P2_U3440, P2_U3441, P2_U3442, P2_U3443, P2_U3444, P2_U3445, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3584, P2_U3589, P2_U3590, P2_U3594, P2_U3597, P2_U3598, P2_U3606, P2_U3607, P2_U3613, P2_U3614, P2_U3615, P2_U3616, P2_U3617, P2_U3618, P2_U3619, P2_U3620, P2_U3621, P2_U3622, P2_U3623, P2_U3624, P2_U3625, P2_U3626, P2_U3627, P2_U3628, P2_U3629, P2_U3630, P2_U3631, P2_U3632, P2_U3633, P2_U3634, P2_U3635, P2_U3636, P2_U3637, P2_U3638, P2_U3639, P2_U3640, P2_U3641, P2_U3642, P2_U3643, P2_U3644, P2_U3645, P2_U3646, P2_U3647, P2_U3648, P2_U3649, P2_U3650, P2_U3651, P2_U3652, P2_U3653, P2_U3654, P2_U3655, P2_U3656, P2_U3657, P2_U3658, P2_U3659, P2_U3660, P2_U3661, P2_U3662, P2_U3663, P2_U3664, P2_U3665, P2_U3666, P2_U3667, P2_U3668, P2_U3669, P2_U3670, P2_U3671, P2_U3672, P2_U3673, P2_U3674, P2_U3675, P2_U3676, P2_U3677, P2_U3678, P2_U3679, P2_U3680, P2_U3681, P2_U3682, P2_U3683, P2_U3684, P2_U3685, P2_U3686, P2_U3687, P2_U3688, P2_U3689, P2_U3690, P2_U3691, P2_U3692, P2_U3693, P2_U3694, P2_U3695, P2_U3696, P2_U3697, P2_U3698, P2_U3699, P2_U3700, P2_U3701, P2_U3702, P2_U3703, P2_U3704, P2_U3705, P2_U3706, P2_U3707, P2_U3708, P2_U3709, P2_U3710, P2_U3711, P2_U3712, P2_U3713, P2_U3714, P2_U3715, P2_U3716, P2_U3717, P2_U3718, P2_U3719, P2_U3720, P2_U3721, P2_U3722, P2_U3723, P2_U3724, P2_U3725, P2_U3726, P2_U3727, P2_U3728, P2_U3729, P2_U3730, P2_U3731, P2_U3732, P2_U3733, P2_U3734, P2_U3735, P2_U3736, P2_U3737, P2_U3738, P2_U3739, P2_U3740, P2_U3741, P2_U3742, P2_U3743, P2_U3744, P2_U3745, P2_U3746, P2_U3747, P2_U3748, P2_U3749, P2_U3750, P2_U3751, P2_U3752, P2_U3753, P2_U3754, P2_U3755, P2_U3756, P2_U3757, P2_U3758, P2_U3759, P2_U3760, P2_U3761, P2_U3762, P2_U3763, P2_U3764, P2_U3765, P2_U3766, P2_U3767, P2_U3768, P2_U3769, P2_U3770, P2_U3771, P2_U3772, P2_U3773, P2_U3774, P2_U3775, P2_U3776, P2_U3777, P2_U3778, P2_U3779, P2_U3780, P2_U3781, P2_U3782, P2_U3783, P2_U3784, P2_U3785, P2_U3786, P2_U3787, P2_U3788, P2_U3789, P2_U3790, P2_U3791, P2_U3792, P2_U3793, P2_U3794, P2_U3795, P2_U3796, P2_U3797, P2_U3798, P2_U3799, P2_U3800, P2_U3801, P2_U3802, P2_U3803, P2_U3804, P2_U3805, P2_U3806, P2_U3807, P2_U3808, P2_U3809, P2_U3810, P2_U3811, P2_U3812, P2_U3813, P2_U3814, P2_U3815, P2_U3816, P2_U3817, P2_U3818, P2_U3819, P2_U3820, P2_U3821, P2_U3822, P2_U3823, P2_U3824, P2_U3825, P2_U3826, P2_U3827, P2_U3828, P2_U3829, P2_U3830, P2_U3831, P2_U3832, P2_U3833, P2_U3834, P2_U3835, P2_U3836, P2_U3837, P2_U3838, P2_U3839, P2_U3840, P2_U3841, P2_U3842, P2_U3843, P2_U3844, P2_U3845, P2_U3846, P2_U3847, P2_U3848, P2_U3849, P2_U3850, P2_U3851, P2_U3852, P2_U3853, P2_U3854, P2_U3855, P2_U3856, P2_U3857, P2_U3858, P2_U3859, P2_U3860, P2_U3861, P2_U3862, P2_U3863, P2_U3864, P2_U3865, P2_U3866, P2_U3867, P2_U3868, P2_U3869, P2_U3870, P2_U3871, P2_U3872, P2_U3873, P2_U3874, P2_U3875, P2_U3876, P2_U3877, P2_U3878, P2_U3879, P2_U3880, P2_U3881, P2_U3882, P2_U3883, P2_U3884, P2_U3885, P2_U3886, P2_U3887, P2_U3888, P2_U3889, P2_U3890, P2_U3891, P2_U3892, P2_U3893, P2_U3894, P2_U3895, P2_U3896, P2_U3897, P2_U3898, P2_U3899, P2_U3900, P2_U3901, P2_U3902, P2_U3903, P2_U3904, P2_U3905, P2_U3906, P2_U3907, P2_U3908, P2_U3909, P2_U3910, P2_U3911, P2_U3912, P2_U3913, P2_U3914, P2_U3915, P2_U3916, P2_U3917, P2_U3918, P2_U3919, P2_U3920, P2_U3921, P2_U3922, P2_U3923, P2_U3924, P2_U3925, P2_U3926, P2_U3927, P2_U3928, P2_U3929, P2_U3930, P2_U3931, P2_U3932, P2_U3933, P2_U3934, P2_U3935, P2_U3936, P2_U3937, P2_U3938, P2_U3939, P2_U3940, P2_U3941, P2_U3942, P2_U3943, P2_U3944, P2_U3945, P2_U3946, P2_U3947, P2_U3948, P2_U3949, P2_U3950, P2_U3951, P2_U3952, P2_U3953, P2_U3954, P2_U3955, P2_U3956, P2_U3957, P2_U3958, P2_U3959, P2_U3960, P2_U3961, P2_U3962, P2_U3963, P2_U3964, P2_U3965, P2_U3966, P2_U3967, P2_U3968, P2_U3969, P2_U3970, P2_U3971, P2_U3972, P2_U3973, P2_U3974, P2_U3975, P2_U3976, P2_U3977, P2_U3978, P2_U3979, P2_U3980, P2_U3981, P2_U3982, P2_U3983, P2_U3984, P2_U3985, P2_U3986, P2_U3987, P2_U3988, P2_U3989, P2_U3990, P2_U3991, P2_U3992, P2_U3993, P2_U3994, P2_U3995, P2_U3996, P2_U3997, P2_U3998, P2_U3999, P2_U4000, P2_U4001, P2_U4002, P2_U4003, P2_U4004, P2_U4005, P2_U4006, P2_U4007, P2_U4008, P2_U4009, P2_U4010, P2_U4011, P2_U4012, P2_U4013, P2_U4014, P2_U4015, P2_U4016, P2_U4017, P2_U4018, P2_U4019, P2_U4020, P2_U4021, P2_U4022, P2_U4023, P2_U4024, P2_U4025, P2_U4026, P2_U4027, P2_U4028, P2_U4029, P2_U4030, P2_U4031, P2_U4032, P2_U4033, P2_U4034, P2_U4035, P2_U4036, P2_U4037, P2_U4038, P2_U4039, P2_U4040, P2_U4041, P2_U4042, P2_U4043, P2_U4044, P2_U4045, P2_U4046, P2_U4047, P2_U4048, P2_U4049, P2_U4050, P2_U4051, P2_U4052, P2_U4053, P2_U4054, P2_U4055, P2_U4056, P2_U4057, P2_U4058, P2_U4059, P2_U4060, P2_U4061, P2_U4062, P2_U4063, P2_U4064, P2_U4065, P2_U4066, P2_U4067, P2_U4068, P2_U4069, P2_U4070, P2_U4071, P2_U4072, P2_U4073, P2_U4074, P2_U4075, P2_U4076, P2_U4077, P2_U4078, P2_U4079, P2_U4080, P2_U4081, P2_U4082, P2_U4083, P2_U4084, P2_U4085, P2_U4086, P2_U4087, P2_U4088, P2_U4089, P2_U4090, P2_U4091, P2_U4092, P2_U4093, P2_U4094, P2_U4095, P2_U4096, P2_U4097, P2_U4098, P2_U4099, P2_U4100, P2_U4101, P2_U4102, P2_U4103, P2_U4104, P2_U4105, P2_U4106, P2_U4107, P2_U4108, P2_U4109, P2_U4110, P2_U4111, P2_U4112, P2_U4113, P2_U4114, P2_U4115, P2_U4116, P2_U4117, P2_U4118, P2_U4119, P2_U4120, P2_U4121, P2_U4122, P2_U4123, P2_U4124, P2_U4125, P2_U4126, P2_U4127, P2_U4128, P2_U4129, P2_U4130, P2_U4131, P2_U4132, P2_U4133, P2_U4134, P2_U4135, P2_U4136, P2_U4137, P2_U4138, P2_U4139, P2_U4140, P2_U4141, P2_U4142, P2_U4143, P2_U4144, P2_U4145, P2_U4146, P2_U4147, P2_U4148, P2_U4149, P2_U4150, P2_U4151, P2_U4152, P2_U4153, P2_U4154, P2_U4155, P2_U4156, P2_U4157, P2_U4158, P2_U4159, P2_U4160, P2_U4161, P2_U4162, P2_U4163, P2_U4164, P2_U4165, P2_U4166, P2_U4167, P2_U4168, P2_U4169, P2_U4170, P2_U4171, P2_U4172, P2_U4173, P2_U4174, P2_U4175, P2_U4176, P2_U4177, P2_U4178, P2_U4179, P2_U4180, P2_U4181, P2_U4182, P2_U4183, P2_U4184, P2_U4185, P2_U4186, P2_U4187, P2_U4188, P2_U4189, P2_U4190, P2_U4191, P2_U4192, P2_U4193, P2_U4194, P2_U4195, P2_U4196, P2_U4197, P2_U4198, P2_U4199, P2_U4200, P2_U4201, P2_U4202, P2_U4203, P2_U4204, P2_U4205, P2_U4206, P2_U4207, P2_U4208, P2_U4209, P2_U4210, P2_U4211, P2_U4212, P2_U4213, P2_U4214, P2_U4215, P2_U4216, P2_U4217, P2_U4218, P2_U4219, P2_U4220, P2_U4221, P2_U4222, P2_U4223, P2_U4224, P2_U4225, P2_U4226, P2_U4227, P2_U4228, P2_U4229, P2_U4230, P2_U4231, P2_U4232, P2_U4233, P2_U4234, P2_U4235, P2_U4236, P2_U4237, P2_U4238, P2_U4239, P2_U4240, P2_U4241, P2_U4242, P2_U4243, P2_U4244, P2_U4245, P2_U4246, P2_U4247, P2_U4248, P2_U4249, P2_U4250, P2_U4251, P2_U4252, P2_U4253, P2_U4254, P2_U4255, P2_U4256, P2_U4257, P2_U4258, P2_U4259, P2_U4260, P2_U4261, P2_U4262, P2_U4263, P2_U4264, P2_U4265, P2_U4266, P2_U4267, P2_U4268, P2_U4269, P2_U4270, P2_U4271, P2_U4272, P2_U4273, P2_U4274, P2_U4275, P2_U4276, P2_U4277, P2_U4278, P2_U4279, P2_U4280, P2_U4281, P2_U4282, P2_U4283, P2_U4284, P2_U4285, P2_U4286, P2_U4287, P2_U4288, P2_U4289, P2_U4290, P2_U4291, P2_U4292, P2_U4293, P2_U4294, P2_U4295, P2_U4296, P2_U4297, P2_U4298, P2_U4299, P2_U4300, P2_U4301, P2_U4302, P2_U4303, P2_U4304, P2_U4305, P2_U4306, P2_U4307, P2_U4308, P2_U4309, P2_U4310, P2_U4311, P2_U4312, P2_U4313, P2_U4314, P2_U4315, P2_U4316, P2_U4317, P2_U4318, P2_U4319, P2_U4320, P2_U4321, P2_U4322, P2_U4323, P2_U4324, P2_U4325, P2_U4326, P2_U4327, P2_U4328, P2_U4329, P2_U4330, P2_U4331, P2_U4332, P2_U4333, P2_U4334, P2_U4335, P2_U4336, P2_U4337, P2_U4338, P2_U4339, P2_U4340, P2_U4341, P2_U4342, P2_U4343, P2_U4344, P2_U4345, P2_U4346, P2_U4347, P2_U4348, P2_U4349, P2_U4350, P2_U4351, P2_U4352, P2_U4353, P2_U4354, P2_U4355, P2_U4356, P2_U4357, P2_U4358, P2_U4359, P2_U4360, P2_U4361, P2_U4362, P2_U4363, P2_U4364, P2_U4365, P2_U4366, P2_U4367, P2_U4368, P2_U4369, P2_U4370, P2_U4371, P2_U4372, P2_U4373, P2_U4374, P2_U4375, P2_U4376, P2_U4377, P2_U4378, P2_U4379, P2_U4380, P2_U4381, P2_U4382, P2_U4383, P2_U4384, P2_U4385, P2_U4386, P2_U4387, P2_U4388, P2_U4389, P2_U4390, P2_U4391, P2_U4392, P2_U4393, P2_U4394, P2_U4395, P2_U4396, P2_U4397, P2_U4398, P2_U4399, P2_U4400, P2_U4401, P2_U4402, P2_U4403, P2_U4404, P2_U4405, P2_U4406, P2_U4407, P2_U4408, P2_U4409, P2_U4410, P2_U4411, P2_U4412, P2_U4413, P2_U4414, P2_U4415, P2_U4416, P2_U4417, P2_U4418, P2_U4419, P2_U4420, P2_U4421, P2_U4422, P2_U4423, P2_U4424, P2_U4425, P2_U4426, P2_U4427, P2_U4428, P2_U4429, P2_U4430, P2_U4431, P2_U4432, P2_U4433, P2_U4434, P2_U4435, P2_U4436, P2_U4437, P2_U4438, P2_U4439, P2_U4440, P2_U4441, P2_U4442, P2_U4443, P2_U4444, P2_U4445, P2_U4446, P2_U4447, P2_U4448, P2_U4449, P2_U4450, P2_U4451, P2_U4452, P2_U4453, P2_U4454, P2_U4455, P2_U4456, P2_U4457, P2_U4458, P2_U4459, P2_U4460, P2_U4461, P2_U4462, P2_U4463, P2_U4464, P2_U4465, P2_U4466, P2_U4467, P2_U4468, P2_U4469, P2_U4470, P2_U4471, P2_U4472, P2_U4473, P2_U4474, P2_U4475, P2_U4476, P2_U4477, P2_U4478, P2_U4479, P2_U4480, P2_U4481, P2_U4482, P2_U4483, P2_U4484, P2_U4485, P2_U4486, P2_U4487, P2_U4488, P2_U4489, P2_U4490, P2_U4491, P2_U4492, P2_U4493, P2_U4494, P2_U4495, P2_U4496, P2_U4497, P2_U4498, P2_U4499, P2_U4500, P2_U4501, P2_U4502, P2_U4503, P2_U4504, P2_U4505, P2_U4506, P2_U4507, P2_U4508, P2_U4509, P2_U4510, P2_U4511, P2_U4512, P2_U4513, P2_U4514, P2_U4515, P2_U4516, P2_U4517, P2_U4518, P2_U4519, P2_U4520, P2_U4521, P2_U4522, P2_U4523, P2_U4524, P2_U4525, P2_U4526, P2_U4527, P2_U4528, P2_U4529, P2_U4530, P2_U4531, P2_U4532, P2_U4533, P2_U4534, P2_U4535, P2_U4536, P2_U4537, P2_U4538, P2_U4539, P2_U4540, P2_U4541, P2_U4542, P2_U4543, P2_U4544, P2_U4545, P2_U4546, P2_U4547, P2_U4548, P2_U4549, P2_U4550, P2_U4551, P2_U4552, P2_U4553, P2_U4554, P2_U4555, P2_U4556, P2_U4557, P2_U4558, P2_U4559, P2_U4560, P2_U4561, P2_U4562, P2_U4563, P2_U4564, P2_U4565, P2_U4566, P2_U4567, P2_U4568, P2_U4569, P2_U4570, P2_U4571, P2_U4572, P2_U4573, P2_U4574, P2_U4575, P2_U4576, P2_U4577, P2_U4578, P2_U4579, P2_U4580, P2_U4581, P2_U4582, P2_U4583, P2_U4584, P2_U4585, P2_U4586, P2_U4587, P2_U4588, P2_U4589, P2_U4590, P2_U4591, P2_U4592, P2_U4593, P2_U4594, P2_U4595, P2_U4596, P2_U4597, P2_U4598, P2_U4599, P2_U4600, P2_U4601, P2_U4602, P2_U4603, P2_U4604, P2_U4605, P2_U4606, P2_U4607, P2_U4608, P2_U4609, P2_U4610, P2_U4611, P2_U4612, P2_U4613, P2_U4614, P2_U4615, P2_U4616, P2_U4617, P2_U4618, P2_U4619, P2_U4620, P2_U4621, P2_U4622, P2_U4623, P2_U4624, P2_U4625, P2_U4626, P2_U4627, P2_U4628, P2_U4629, P2_U4630, P2_U4631, P2_U4632, P2_U4633, P2_U4634, P2_U4635, P2_U4636, P2_U4637, P2_U4638, P2_U4639, P2_U4640, P2_U4641, P2_U4642, P2_U4643, P2_U4644, P2_U4645, P2_U4646, P2_U4647, P2_U4648, P2_U4649, P2_U4650, P2_U4651, P2_U4652, P2_U4653, P2_U4654, P2_U4655, P2_U4656, P2_U4657, P2_U4658, P2_U4659, P2_U4660, P2_U4661, P2_U4662, P2_U4663, P2_U4664, P2_U4665, P2_U4666, P2_U4667, P2_U4668, P2_U4669, P2_U4670, P2_U4671, P2_U4672, P2_U4673, P2_U4674, P2_U4675, P2_U4676, P2_U4677, P2_U4678, P2_U4679, P2_U4680, P2_U4681, P2_U4682, P2_U4683, P2_U4684, P2_U4685, P2_U4686, P2_U4687, P2_U4688, P2_U4689, P2_U4690, P2_U4691, P2_U4692, P2_U4693, P2_U4694, P2_U4695, P2_U4696, P2_U4697, P2_U4698, P2_U4699, P2_U4700, P2_U4701, P2_U4702, P2_U4703, P2_U4704, P2_U4705, P2_U4706, P2_U4707, P2_U4708, P2_U4709, P2_U4710, P2_U4711, P2_U4712, P2_U4713, P2_U4714, P2_U4715, P2_U4716, P2_U4717, P2_U4718, P2_U4719, P2_U4720, P2_U4721, P2_U4722, P2_U4723, P2_U4724, P2_U4725, P2_U4726, P2_U4727, P2_U4728, P2_U4729, P2_U4730, P2_U4731, P2_U4732, P2_U4733, P2_U4734, P2_U4735, P2_U4736, P2_U4737, P2_U4738, P2_U4739, P2_U4740, P2_U4741, P2_U4742, P2_U4743, P2_U4744, P2_U4745, P2_U4746, P2_U4747, P2_U4748, P2_U4749, P2_U4750, P2_U4751, P2_U4752, P2_U4753, P2_U4754, P2_U4755, P2_U4756, P2_U4757, P2_U4758, P2_U4759, P2_U4760, P2_U4761, P2_U4762, P2_U4763, P2_U4764, P2_U4765, P2_U4766, P2_U4767, P2_U4768, P2_U4769, P2_U4770, P2_U4771, P2_U4772, P2_U4773, P2_U4774, P2_U4775, P2_U4776, P2_U4777, P2_U4778, P2_U4779, P2_U4780, P2_U4781, P2_U4782, P2_U4783, P2_U4784, P2_U4785, P2_U4786, P2_U4787, P2_U4788, P2_U4789, P2_U4790, P2_U4791, P2_U4792, P2_U4793, P2_U4794, P2_U4795, P2_U4796, P2_U4797, P2_U4798, P2_U4799, P2_U4800, P2_U4801, P2_U4802, P2_U4803, P2_U4804, P2_U4805, P2_U4806, P2_U4807, P2_U4808, P2_U4809, P2_U4810, P2_U4811, P2_U4812, P2_U4813, P2_U4814, P2_U4815, P2_U4816, P2_U4817, P2_U4818, P2_U4819, P2_U4820, P2_U4821, P2_U4822, P2_U4823, P2_U4824, P2_U4825, P2_U4826, P2_U4827, P2_U4828, P2_U4829, P2_U4830, P2_U4831, P2_U4832, P2_U4833, P2_U4834, P2_U4835, P2_U4836, P2_U4837, P2_U4838, P2_U4839, P2_U4840, P2_U4841, P2_U4842, P2_U4843, P2_U4844, P2_U4845, P2_U4846, P2_U4847, P2_U4848, P2_U4849, P2_U4850, P2_U4851, P2_U4852, P2_U4853, P2_U4854, P2_U4855, P2_U4856, P2_U4857, P2_U4858, P2_U4859, P2_U4860, P2_U4861, P2_U4862, P2_U4863, P2_U4864, P2_U4865, P2_U4866, P2_U4867, P2_U4868, P2_U4869, P2_U4870, P2_U4871, P2_U4872, P2_U4873, P2_U4874, P2_U4875, P2_U4876, P2_U4877, P2_U4878, P2_U4879, P2_U4880, P2_U4881, P2_U4882, P2_U4883, P2_U4884, P2_U4885, P2_U4886, P2_U4887, P2_U4888, P2_U4889, P2_U4890, P2_U4891, P2_U4892, P2_U4893, P2_U4894, P2_U4895, P2_U4896, P2_U4897, P2_U4898, P2_U4899, P2_U4900, P2_U4901, P2_U4902, P2_U4903, P2_U4904, P2_U4905, P2_U4906, P2_U4907, P2_U4908, P2_U4909, P2_U4910, P2_U4911, P2_U4912, P2_U4913, P2_U4914, P2_U4915, P2_U4916, P2_U4917, P2_U4918, P2_U4919, P2_U4920, P2_U4921, P2_U4922, P2_U4923, P2_U4924, P2_U4925, P2_U4926, P2_U4927, P2_U4928, P2_U4929, P2_U4930, P2_U4931, P2_U4932, P2_U4933, P2_U4934, P2_U4935, P2_U4936, P2_U4937, P2_U4938, P2_U4939, P2_U4940, P2_U4941, P2_U4942, P2_U4943, P2_U4944, P2_U4945, P2_U4946, P2_U4947, P2_U4948, P2_U4949, P2_U4950, P2_U4951, P2_U4952, P2_U4953, P2_U4954, P2_U4955, P2_U4956, P2_U4957, P2_U4958, P2_U4959, P2_U4960, P2_U4961, P2_U4962, P2_U4963, P2_U4964, P2_U4965, P2_U4966, P2_U4967, P2_U4968, P2_U4969, P2_U4970, P2_U4971, P2_U4972, P2_U4973, P2_U4974, P2_U4975, P2_U4976, P2_U4977, P2_U4978, P2_U4979, P2_U4980, P2_U4981, P2_U4982, P2_U4983, P2_U4984, P2_U4985, P2_U4986, P2_U4987, P2_U4988, P2_U4989, P2_U4990, P2_U4991, P2_U4992, P2_U4993, P2_U4994, P2_U4995, P2_U4996, P2_U4997, P2_U4998, P2_U4999, P2_U5000, P2_U5001, P2_U5002, P2_U5003, P2_U5004, P2_U5005, P2_U5006, P2_U5007, P2_U5008, P2_U5009, P2_U5010, P2_U5011, P2_U5012, P2_U5013, P2_U5014, P2_U5015, P2_U5016, P2_U5017, P2_U5018, P2_U5019, P2_U5020, P2_U5021, P2_U5022, P2_U5023, P2_U5024, P2_U5025, P2_U5026, P2_U5027, P2_U5028, P2_U5029, P2_U5030, P2_U5031, P2_U5032, P2_U5033, P2_U5034, P2_U5035, P2_U5036, P2_U5037, P2_U5038, P2_U5039, P2_U5040, P2_U5041, P2_U5042, P2_U5043, P2_U5044, P2_U5045, P2_U5046, P2_U5047, P2_U5048, P2_U5049, P2_U5050, P2_U5051, P2_U5052, P2_U5053, P2_U5054, P2_U5055, P2_U5056, P2_U5057, P2_U5058, P2_U5059, P2_U5060, P2_U5061, P2_U5062, P2_U5063, P2_U5064, P2_U5065, P2_U5066, P2_U5067, P2_U5068, P2_U5069, P2_U5070, P2_U5071, P2_U5072, P2_U5073, P2_U5074, P2_U5075, P2_U5076, P2_U5077, P2_U5078, P2_U5079, P2_U5080, P2_U5081, P2_U5082, P2_U5083, P2_U5084, P2_U5085, P2_U5086, P2_U5087, P2_U5088, P2_U5089, P2_U5090, P2_U5091, P2_U5092, P2_U5093, P2_U5094, P2_U5095, P2_U5096, P2_U5097, P2_U5098, P2_U5099, P2_U5100, P2_U5101, P2_U5102, P2_U5103, P2_U5104, P2_U5105, P2_U5106, P2_U5107, P2_U5108, P2_U5109, P2_U5110, P2_U5111, P2_U5112, P2_U5113, P2_U5114, P2_U5115, P2_U5116, P2_U5117, P2_U5118, P2_U5119, P2_U5120, P2_U5121, P2_U5122, P2_U5123, P2_U5124, P2_U5125, P2_U5126, P2_U5127, P2_U5128, P2_U5129, P2_U5130, P2_U5131, P2_U5132, P2_U5133, P2_U5134, P2_U5135, P2_U5136, P2_U5137, P2_U5138, P2_U5139, P2_U5140, P2_U5141, P2_U5142, P2_U5143, P2_U5144, P2_U5145, P2_U5146, P2_U5147, P2_U5148, P2_U5149, P2_U5150, P2_U5151, P2_U5152, P2_U5153, P2_U5154, P2_U5155, P2_U5156, P2_U5157, P2_U5158, P2_U5159, P2_U5160, P2_U5161, P2_U5162, P2_U5163, P2_U5164, P2_U5165, P2_U5166, P2_U5167, P2_U5168, P2_U5169, P2_U5170, P2_U5171, P2_U5172, P2_U5173, P2_U5174, P2_U5175, P2_U5176, P2_U5177, P2_U5178, P2_U5179, P2_U5180, P2_U5181, P2_U5182, P2_U5183, P2_U5184, P2_U5185, P2_U5186, P2_U5187, P2_U5188, P2_U5189, P2_U5190, P2_U5191, P2_U5192, P2_U5193, P2_U5194, P2_U5195, P2_U5196, P2_U5197, P2_U5198, P2_U5199, P2_U5200, P2_U5201, P2_U5202, P2_U5203, P2_U5204, P2_U5205, P2_U5206, P2_U5207, P2_U5208, P2_U5209, P2_U5210, P2_U5211, P2_U5212, P2_U5213, P2_U5214, P2_U5215, P2_U5216, P2_U5217, P2_U5218, P2_U5219, P2_U5220, P2_U5221, P2_U5222, P2_U5223, P2_U5224, P2_U5225, P2_U5226, P2_U5227, P2_U5228, P2_U5229, P2_U5230, P2_U5231, P2_U5232, P2_U5233, P2_U5234, P2_U5235, P2_U5236, P2_U5237, P2_U5238, P2_U5239, P2_U5240, P2_U5241, P2_U5242, P2_U5243, P2_U5244, P2_U5245, P2_U5246, P2_U5247, P2_U5248, P2_U5249, P2_U5250, P2_U5251, P2_U5252, P2_U5253, P2_U5254, P2_U5255, P2_U5256, P2_U5257, P2_U5258, P2_U5259, P2_U5260, P2_U5261, P2_U5262, P2_U5263, P2_U5264, P2_U5265, P2_U5266, P2_U5267, P2_U5268, P2_U5269, P2_U5270, P2_U5271, P2_U5272, P2_U5273, P2_U5274, P2_U5275, P2_U5276, P2_U5277, P2_U5278, P2_U5279, P2_U5280, P2_U5281, P2_U5282, P2_U5283, P2_U5284, P2_U5285, P2_U5286, P2_U5287, P2_U5288, P2_U5289, P2_U5290, P2_U5291, P2_U5292, P2_U5293, P2_U5294, P2_U5295, P2_U5296, P2_U5297, P2_U5298, P2_U5299, P2_U5300, P2_U5301, P2_U5302, P2_U5303, P2_U5304, P2_U5305, P2_U5306, P2_U5307, P2_U5308, P2_U5309, P2_U5310, P2_U5311, P2_U5312, P2_U5313, P2_U5314, P2_U5315, P2_U5316, P2_U5317, P2_U5318, P2_U5319, P2_U5320, P2_U5321, P2_U5322, P2_U5323, P2_U5324, P2_U5325, P2_U5326, P2_U5327, P2_U5328, P2_U5329, P2_U5330, P2_U5331, P2_U5332, P2_U5333, P2_U5334, P2_U5335, P2_U5336, P2_U5337, P2_U5338, P2_U5339, P2_U5340, P2_U5341, P2_U5342, P2_U5343, P2_U5344, P2_U5345, P2_U5346, P2_U5347, P2_U5348, P2_U5349, P2_U5350, P2_U5351, P2_U5352, P2_U5353, P2_U5354, P2_U5355, P2_U5356, P2_U5357, P2_U5358, P2_U5359, P2_U5360, P2_U5361, P2_U5362, P2_U5363, P2_U5364, P2_U5365, P2_U5366, P2_U5367, P2_U5368, P2_U5369, P2_U5370, P2_U5371, P2_U5372, P2_U5373, P2_U5374, P2_U5375, P2_U5376, P2_U5377, P2_U5378, P2_U5379, P2_U5380, P2_U5381, P2_U5382, P2_U5383, P2_U5384, P2_U5385, P2_U5386, P2_U5387, P2_U5388, P2_U5389, P2_U5390, P2_U5391, P2_U5392, P2_U5393, P2_U5394, P2_U5395, P2_U5396, P2_U5397, P2_U5398, P2_U5399, P2_U5400, P2_U5401, P2_U5402, P2_U5403, P2_U5404, P2_U5405, P2_U5406, P2_U5407, P2_U5408, P2_U5409, P2_U5410, P2_U5411, P2_U5412, P2_U5413, P2_U5414, P2_U5415, P2_U5416, P2_U5417, P2_U5418, P2_U5419, P2_U5420, P2_U5421, P2_U5422, P2_U5423, P2_U5424, P2_U5425, P2_U5426, P2_U5427, P2_U5428, P2_U5429, P2_U5430, P2_U5431, P2_U5432, P2_U5433, P2_U5434, P2_U5435, P2_U5436, P2_U5437, P2_U5438, P2_U5439, P2_U5440, P2_U5441, P2_U5442, P2_U5443, P2_U5444, P2_U5445, P2_U5446, P2_U5447, P2_U5448, P2_U5449, P2_U5450, P2_U5451, P2_U5452, P2_U5453, P2_U5454, P2_U5455, P2_U5456, P2_U5457, P2_U5458, P2_U5459, P2_U5460, P2_U5461, P2_U5462, P2_U5463, P2_U5464, P2_U5465, P2_U5466, P2_U5467, P2_U5468, P2_U5469, P2_U5470, P2_U5471, P2_U5472, P2_U5473, P2_U5474, P2_U5475, P2_U5476, P2_U5477, P2_U5478, P2_U5479, P2_U5480, P2_U5481, P2_U5482, P2_U5483, P2_U5484, P2_U5485, P2_U5486, P2_U5487, P2_U5488, P2_U5489, P2_U5490, P2_U5491, P2_U5492, P2_U5493, P2_U5494, P2_U5495, P2_U5496, P2_U5497, P2_U5498, P2_U5499, P2_U5500, P2_U5501, P2_U5502, P2_U5503, P2_U5504, P2_U5505, P2_U5506, P2_U5507, P2_U5508, P2_U5509, P2_U5510, P2_U5511, P2_U5512, P2_U5513, P2_U5514, P2_U5515, P2_U5516, P2_U5517, P2_U5518, P2_U5519, P2_U5520, P2_U5521, P2_U5522, P2_U5523, P2_U5524, P2_U5525, P2_U5526, P2_U5527, P2_U5528, P2_U5529, P2_U5530, P2_U5531, P2_U5532, P2_U5533, P2_U5534, P2_U5535, P2_U5536, P2_U5537, P2_U5538, P2_U5539, P2_U5540, P2_U5541, P2_U5542, P2_U5543, P2_U5544, P2_U5545, P2_U5546, P2_U5547, P2_U5548, P2_U5549, P2_U5550, P2_U5551, P2_U5552, P2_U5553, P2_U5554, P2_U5555, P2_U5556, P2_U5557, P2_U5558, P2_U5559, P2_U5560, P2_U5561, P2_U5562, P2_U5563, P2_U5564, P2_U5565, P2_U5566, P2_U5567, P2_U5568, P2_U5569, P2_U5570, P2_U5571, P2_U5572, P2_U5573, P2_U5574, P2_U5575, P2_U5576, P2_U5577, P2_U5578, P2_U5579, P2_U5580, P2_U5581, P2_U5582, P2_U5583, P2_U5584, P2_U5585, P2_U5586, P2_U5587, P2_U5588, P2_U5589, P2_U5590, P2_U5591, P2_U5592, P2_U5593, P2_U5594, P2_U5595, P2_U5596, P2_U5597, P2_U5598, P2_U5599, P2_U5600, P2_U5601, P2_U5602, P2_U5603, P2_U5604, P2_U5605, P2_U5606, P2_U5607, P2_U5608, P2_U5609, P2_U5610, P2_U5611, P2_U5612, P2_U5613, P2_U5614, P2_U5615, P2_U5616, P2_U5617, P2_U5618, P2_U5619, P2_U5620, P2_U5621, P2_U5622, P2_U5623, P2_U5624, P2_U5625, P2_U5626, P2_U5627, P2_U5628, P2_U5629, P2_U5630, P2_U5631, P2_U5632, P2_U5633, P2_U5634, P2_U5635, P2_U5636, P2_U5637, P2_U5638, P2_U5639, P2_U5640, P2_U5641, P2_U5642, P2_U5643, P2_U5644, P2_U5645, P2_U5646, P2_U5647, P2_U5648, P2_U5649, P2_U5650, P2_U5651, P2_U5652, P2_U5653, P2_U5654, P2_U5655, P2_U5656, P2_U5657, P2_U5658, P2_U5659, P2_U5660, P2_U5661, P2_U5662, P2_U5663, P2_U5664, P2_U5665, P2_U5666, P2_U5667, P2_U5668, P2_U5669, P2_U5670, P2_U5671, P2_U5672, P2_U5673, P2_U5674, P2_U5675, P2_U5676, P2_U5677, P2_U5678, P2_U5679, P2_U5680, P2_U5681, P2_U5682, P2_U5683, P2_U5684, P2_U5685, P2_U5686, P2_U5687, P2_U5688, P2_U5689, P2_U5690, P2_U5691, P2_U5692, P2_U5693, P2_U5694, P2_U5695, P2_U5696, P2_U5697, P2_U5698, P2_U5699, P2_U5700, P2_U5701, P2_U5702, P2_U5703, P2_U5704, P2_U5705, P2_U5706, P2_U5707, P2_U5708, P2_U5709, P2_U5710, P2_U5711, P2_U5712, P2_U5713, P2_U5714, P2_U5715, P2_U5716, P2_U5717, P2_U5718, P2_U5719, P2_U5720, P2_U5721, P2_U5722, P2_U5723, P2_U5724, P2_U5725, P2_U5726, P2_U5727, P2_U5728, P2_U5729, P2_U5730, P2_U5731, P2_U5732, P2_U5733, P2_U5734, P2_U5735, P2_U5736, P2_U5737, P2_U5738, P2_U5739, P2_U5740, P2_U5741, P2_U5742, P2_U5743, P2_U5744, P2_U5745, P2_U5746, P2_U5747, P2_U5748, P2_U5749, P2_U5750, P2_U5751, P2_U5752, P2_U5753, P2_U5754, P2_U5755, P2_U5756, P2_U5757, P2_U5758, P2_U5759, P2_U5760, P2_U5761, P2_U5762, P2_U5763, P2_U5764, P2_U5765, P2_U5766, P2_U5767, P2_U5768, P2_U5769, P2_U5770, P2_U5771, P2_U5772, P2_U5773, P2_U5774, P2_U5775, P2_U5776, P2_U5777, P2_U5778, P2_U5779, P2_U5780, P2_U5781, P2_U5782, P2_U5783, P2_U5784, P2_U5785, P2_U5786, P2_U5787, P2_U5788, P2_U5789, P2_U5790, P2_U5791, P2_U5792, P2_U5793, P2_U5794, P2_U5795, P2_U5796, P2_U5797, P2_U5798, P2_U5799, P2_U5800, P2_U5801, P2_U5802, P2_U5803, P2_U5804, P2_U5805, P2_U5806, P2_U5807, P2_U5808, P2_U5809, P2_U5810, P2_U5811, P2_U5812, P2_U5813, P2_U5814, P2_U5815, P2_U5816, P2_U5817, P2_U5818, P2_U5819, P2_U5820, P2_U5821, P2_U5822, P2_U5823, P2_U5824, P2_U5825, P2_U5826, P2_U5827, P2_U5828, P2_U5829, P2_U5830, P2_U5831, P2_U5832, P2_U5833, P2_U5834, P2_U5835, P2_U5836, P2_U5837, P2_U5838, P2_U5839, P2_U5840, P2_U5841, P2_U5842, P2_U5843, P2_U5844, P2_U5845, P2_U5846, P2_U5847, P2_U5848, P2_U5849, P2_U5850, P2_U5851, P2_U5852, P2_U5853, P2_U5854, P2_U5855, P2_U5856, P2_U5857, P2_U5858, P2_U5859, P2_U5860, P2_U5861, P2_U5862, P2_U5863, P2_U5864, P2_U5865, P2_U5866, P2_U5867, P2_U5868, P2_U5869, P2_U5870, P2_U5871, P2_U5872, P2_U5873, P2_U5874, P2_U5875, P2_U5876, P2_U5877, P2_U5878, P2_U5879, P2_U5880, P2_U5881, P2_U5882, P2_U5883, P2_U5884, P2_U5885, P2_U5886, P2_U5887, P2_U5888, P2_U5889, P2_U5890, P2_U5891, P2_U5892, P2_U5893, P2_U5894, P2_U5895, P2_U5896, P2_U5897, P2_U5898, P2_U5899, P2_U5900, P2_U5901, P2_U5902, P2_U5903, P2_U5904, P2_U5905, P2_U5906, P2_U5907, P2_U5908, P2_U5909, P2_U5910, P2_U5911, P2_U5912, P2_U5913, P2_U5914, P2_U5915, P2_U5916, P2_U5917, P2_U5918, P2_U5919, P2_U5920, P2_U5921, P2_U5922, P2_U5923, P2_U5924, P2_U5925, P2_U5926, P2_U5927, P2_U5928, P2_U5929, P2_U5930, P2_U5931, P2_U5932, P2_U5933, P2_U5934, P2_U5935, P2_U5936, P2_U5937, P2_U5938, P2_U5939, P2_U5940, P2_U5941, P2_U5942, P2_U5943, P2_U5944, P2_U5945, P2_U5946, P2_U5947, P2_U5948, P2_U5949, P2_U5950, P2_U5951, P2_U5952, P2_U5953, P2_U5954, P2_U5955, P2_U5956, P2_U5957, P2_U5958, P2_U5959, P2_U5960, P2_U5961, P2_U5962, P2_U5963, P2_U5964, P2_U5965, P2_U5966, P2_U5967, P2_U5968, P2_U5969, P2_U5970, P2_U5971, P2_U5972, P2_U5973, P2_U5974, P2_U5975, P2_U5976, P2_U5977, P2_U5978, P2_U5979, P2_U5980, P2_U5981, P2_U5982, P2_U5983, P2_U5984, P2_U5985, P2_U5986, P2_U5987, P2_U5988, P2_U5989, P2_U5990, P2_U5991, P2_U5992, P2_U5993, P2_U5994, P2_U5995, P2_U5996, P2_U5997, P2_U5998, P2_U5999, P2_U6000, P2_U6001, P2_U6002, P2_U6003, P2_U6004, P2_U6005, P2_U6006, P2_U6007, P2_U6008, P2_U6009, P2_U6010, P2_U6011, P2_U6012, P2_U6013, P2_U6014, P2_U6015, P2_U6016, P2_U6017, P2_U6018, P2_U6019, P2_U6020, P2_U6021, P2_U6022, P2_U6023, P2_U6024, P2_U6025, P2_U6026, P2_U6027, P2_U6028, P2_U6029, P2_U6030, P2_U6031, P2_U6032, P2_U6033, P2_U6034, P2_U6035, P2_U6036, P2_U6037, P2_U6038, P2_U6039, P2_U6040, P2_U6041, P2_U6042, P2_U6043, P2_U6044, P2_U6045, P2_U6046, P2_U6047, P2_U6048, P2_U6049, P2_U6050, P2_U6051, P2_U6052, P2_U6053, P2_U6054, P2_U6055, P2_U6056, P2_U6057, P2_U6058, P2_U6059, P2_U6060, P2_U6061, P2_U6062, P2_U6063, P2_U6064, P2_U6065, P2_U6066, P2_U6067, P2_U6068, P2_U6069, P2_U6070, P2_U6071, P2_U6072, P2_U6073, P2_U6074, P2_U6075, P2_U6076, P2_U6077, P2_U6078, P2_U6079, P2_U6080, P2_U6081, P2_U6082, P2_U6083, P2_U6084, P2_U6085, P2_U6086, P2_U6087, P2_U6088, P2_U6089, P2_U6090, P2_U6091, P2_U6092, P2_U6093, P2_U6094, P2_U6095, P2_U6096, P2_U6097, P2_U6098, P2_U6099, P2_U6100, P2_U6101, P2_U6102, P2_U6103, P2_U6104, P2_U6105, P2_U6106, P2_U6107, P2_U6108, P2_U6109, P2_U6110, P2_U6111, P2_U6112, P2_U6113, P2_U6114, P2_U6115, P2_U6116, P2_U6117, P2_U6118, P2_U6119, P2_U6120, P2_U6121, P2_U6122, P2_U6123, P2_U6124, P2_U6125, P2_U6126, P2_U6127, P2_U6128, P2_U6129, P2_U6130, P2_U6131, P2_U6132, P2_U6133, P2_U6134, P2_U6135, P2_U6136, P2_U6137, P2_U6138, P2_U6139, P2_U6140, P2_U6141, P2_U6142, P2_U6143, P2_U6144, P2_U6145, P2_U6146, P2_U6147, P2_U6148, P2_U6149, P2_U6150, P2_U6151, P2_U6152, P2_U6153, P2_U6154, P2_U6155, P2_U6156, P2_U6157, P2_U6158, P2_U6159, P2_U6160, P2_U6161, P2_U6162, P2_U6163, P2_U6164, P2_U6165, P2_U6166, P2_U6167, P2_U6168, P2_U6169, P2_U6170, P2_U6171, P2_U6172, P2_U6173, P2_U6174, P2_U6175, P2_U6176, P2_U6177, P2_U6178, P2_U6179, P2_U6180, P2_U6181, P2_U6182, P2_U6183, P2_U6184, P2_U6185, P2_U6186, P2_U6187, P2_U6188, P2_U6189, P2_U6190, P2_U6191, P2_U6192, P2_U6193, P2_U6194, P2_U6195, P2_U6196, P2_U6197, P2_U6198, P2_U6199, P2_U6200, P2_U6201, P2_U6202, P2_U6203, P2_U6204, P2_U6205, P2_U6206, P2_U6207, P2_U6208, P2_U6209, P2_U6210, P2_U6211, P2_U6212, P2_U6213, P2_U6214, P2_U6215, P2_U6216, P2_U6217, P2_U6218, P2_U6219, P2_U6220, P2_U6221, P2_U6222, P2_U6223, P2_U6224, P2_U6225, P2_U6226, P2_U6227, P2_U6228, P2_U6229, P2_U6230, P2_U6231, P2_U6232, P2_U6233, P2_U6234, P2_U6235, P2_U6236, P2_U6237, P2_U6238, P2_U6239, P2_U6240, P2_U6241, P2_U6242, P2_U6243, P2_U6244, P2_U6245, P2_U6246, P2_U6247, P2_U6248, P2_U6249, P2_U6250, P2_U6251, P2_U6252, P2_U6253, P2_U6254, P2_U6255, P2_U6256, P2_U6257, P2_U6258, P2_U6259, P2_U6260, P2_U6261, P2_U6262, P2_U6263, P2_U6264, P2_U6265, P2_U6266, P2_U6267, P2_U6268, P2_U6269, P2_U6270, P2_U6271, P2_U6272, P2_U6273, P2_U6274, P2_U6275, P2_U6276, P2_U6277, P2_U6278, P2_U6279, P2_U6280, P2_U6281, P2_U6282, P2_U6283, P2_U6284, P2_U6285, P2_U6286, P2_U6287, P2_U6288, P2_U6289, P2_U6290, P2_U6291, P2_U6292, P2_U6293, P2_U6294, P2_U6295, P2_U6296, P2_U6297, P2_U6298, P2_U6299, P2_U6300, P2_U6301, P2_U6302, P2_U6303, P2_U6304, P2_U6305, P2_U6306, P2_U6307, P2_U6308, P2_U6309, P2_U6310, P2_U6311, P2_U6312, P2_U6313, P2_U6314, P2_U6315, P2_U6316, P2_U6317, P2_U6318, P2_U6319, P2_U6320, P2_U6321, P2_U6322, P2_U6323, P2_U6324, P2_U6325, P2_U6326, P2_U6327, P2_U6328, P2_U6329, P2_U6330, P2_U6331, P2_U6332, P2_U6333, P2_U6334, P2_U6335, P2_U6336, P2_U6337, P2_U6338, P2_U6339, P2_U6340, P2_U6341, P2_U6342, P2_U6343, P2_U6344, P2_U6345, P2_U6346, P2_U6347, P2_U6348, P2_U6349, P2_U6350, P2_U6351, P2_U6352, P2_U6353, P2_U6354, P2_U6355, P2_U6356, P2_U6357, P2_U6358, P2_U6359, P2_U6360, P2_U6361, P2_U6362, P2_U6363, P2_U6364, P2_U6365, P2_U6366, P2_U6367, P2_U6368, P2_U6369, P2_U6370, P2_U6371, P2_U6372, P2_U6373, P2_U6374, P2_U6375, P2_U6376, P2_U6377, P2_U6378, P2_U6379, P2_U6380, P2_U6381, P2_U6382, P2_U6383, P2_U6384, P2_U6385, P2_U6386, P2_U6387, P2_U6388, P2_U6389, P2_U6390, P2_U6391, P2_U6392, P2_U6393, P2_U6394, P2_U6395, P2_U6396, P2_U6397, P2_U6398, P2_U6399, P2_U6400, P2_U6401, P2_U6402, P2_U6403, P2_U6404, P2_U6405, P2_U6406, P2_U6407, P2_U6408, P2_U6409, P2_U6410, P2_U6411, P2_U6412, P2_U6413, P2_U6414, P2_U6415, P2_U6416, P2_U6417, P2_U6418, P2_U6419, P2_U6420, P2_U6421, P2_U6422, P2_U6423, P2_U6424, P2_U6425, P2_U6426, P2_U6427, P2_U6428, P2_U6429, P2_U6430, P2_U6431, P2_U6432, P2_U6433, P2_U6434, P2_U6435, P2_U6436, P2_U6437, P2_U6438, P2_U6439, P2_U6440, P2_U6441, P2_U6442, P2_U6443, P2_U6444, P2_U6445, P2_U6446, P2_U6447, P2_U6448, P2_U6449, P2_U6450, P2_U6451, P2_U6452, P2_U6453, P2_U6454, P2_U6455, P2_U6456, P2_U6457, P2_U6458, P2_U6459, P2_U6460, P2_U6461, P2_U6462, P2_U6463, P2_U6464, P2_U6465, P2_U6466, P2_U6467, P2_U6468, P2_U6469, P2_U6470, P2_U6471, P2_U6472, P2_U6473, P2_U6474, P2_U6475, P2_U6476, P2_U6477, P2_U6478, P2_U6479, P2_U6480, P2_U6481, P2_U6482, P2_U6483, P2_U6484, P2_U6485, P2_U6486, P2_U6487, P2_U6488, P2_U6489, P2_U6490, P2_U6491, P2_U6492, P2_U6493, P2_U6494, P2_U6495, P2_U6496, P2_U6497, P2_U6498, P2_U6499, P2_U6500, P2_U6501, P2_U6502, P2_U6503, P2_U6504, P2_U6505, P2_U6506, P2_U6507, P2_U6508, P2_U6509, P2_U6510, P2_U6511, P2_U6512, P2_U6513, P2_U6514, P2_U6515, P2_U6516, P2_U6517, P2_U6518, P2_U6519, P2_U6520, P2_U6521, P2_U6522, P2_U6523, P2_U6524, P2_U6525, P2_U6526, P2_U6527, P2_U6528, P2_U6529, P2_U6530, P2_U6531, P2_U6532, P2_U6533, P2_U6534, P2_U6535, P2_U6536, P2_U6537, P2_U6538, P2_U6539, P2_U6540, P2_U6541, P2_U6542, P2_U6543, P2_U6544, P2_U6545, P2_U6546, P2_U6547, P2_U6548, P2_U6549, P2_U6550, P2_U6551, P2_U6552, P2_U6553, P2_U6554, P2_U6555, P2_U6556, P2_U6557, P2_U6558, P2_U6559, P2_U6560, P2_U6561, P2_U6562, P2_U6563, P2_U6564, P2_U6565, P2_U6566, P2_U6567, P2_U6568, P2_U6569, P2_U6570, P2_U6571, P2_U6572, P2_U6573, P2_U6574, P2_U6575, P2_U6576, P2_U6577, P2_U6578, P2_U6579, P2_U6580, P2_U6581, P2_U6582, P2_U6583, P2_U6584, P2_U6585, P2_U6586, P2_U6587, P2_U6588, P2_U6589, P2_U6590, P2_U6591, P2_U6592, P2_U6593, P2_U6594, P2_U6595, P2_U6596, P2_U6597, P2_U6598, P2_U6599, P2_U6600, P2_U6601, P2_U6602, P2_U6603, P2_U6604, P2_U6605, P2_U6606, P2_U6607, P2_U6608, P2_U6609, P2_U6610, P2_U6611, P2_U6612, P2_U6613, P2_U6614, P2_U6615, P2_U6616, P2_U6617, P2_U6618, P2_U6619, P2_U6620, P2_U6621, P2_U6622, P2_U6623, P2_U6624, P2_U6625, P2_U6626, P2_U6627, P2_U6628, P2_U6629, P2_U6630, P2_U6631, P2_U6632, P2_U6633, P2_U6634, P2_U6635, P2_U6636, P2_U6637, P2_U6638, P2_U6639, P2_U6640, P2_U6641, P2_U6642, P2_U6643, P2_U6644, P2_U6645, P2_U6646, P2_U6647, P2_U6648, P2_U6649, P2_U6650, P2_U6651, P2_U6652, P2_U6653, P2_U6654, P2_U6655, P2_U6656, P2_U6657, P2_U6658, P2_U6659, P2_U6660, P2_U6661, P2_U6662, P2_U6663, P2_U6664, P2_U6665, P2_U6666, P2_U6667, P2_U6668, P2_U6669, P2_U6670, P2_U6671, P2_U6672, P2_U6673, P2_U6674, P2_U6675, P2_U6676, P2_U6677, P2_U6678, P2_U6679, P2_U6680, P2_U6681, P2_U6682, P2_U6683, P2_U6684, P2_U6685, P2_U6686, P2_U6687, P2_U6688, P2_U6689, P2_U6690, P2_U6691, P2_U6692, P2_U6693, P2_U6694, P2_U6695, P2_U6696, P2_U6697, P2_U6698, P2_U6699, P2_U6700, P2_U6701, P2_U6702, P2_U6703, P2_U6704, P2_U6705, P2_U6706, P2_U6707, P2_U6708, P2_U6709, P2_U6710, P2_U6711, P2_U6712, P2_U6713, P2_U6714, P2_U6715, P2_U6716, P2_U6717, P2_U6718, P2_U6719, P2_U6720, P2_U6721, P2_U6722, P2_U6723, P2_U6724, P2_U6725, P2_U6726, P2_U6727, P2_U6728, P2_U6729, P2_U6730, P2_U6731, P2_U6732, P2_U6733, P2_U6734, P2_U6735, P2_U6736, P2_U6737, P2_U6738, P2_U6739, P2_U6740, P2_U6741, P2_U6742, P2_U6743, P2_U6744, P2_U6745, P2_U6746, P2_U6747, P2_U6748, P2_U6749, P2_U6750, P2_U6751, P2_U6752, P2_U6753, P2_U6754, P2_U6755, P2_U6756, P2_U6757, P2_U6758, P2_U6759, P2_U6760, P2_U6761, P2_U6762, P2_U6763, P2_U6764, P2_U6765, P2_U6766, P2_U6767, P2_U6768, P2_U6769, P2_U6770, P2_U6771, P2_U6772, P2_U6773, P2_U6774, P2_U6775, P2_U6776, P2_U6777, P2_U6778, P2_U6779, P2_U6780, P2_U6781, P2_U6782, P2_U6783, P2_U6784, P2_U6785, P2_U6786, P2_U6787, P2_U6788, P2_U6789, P2_U6790, P2_U6791, P2_U6792, P2_U6793, P2_U6794, P2_U6795, P2_U6796, P2_U6797, P2_U6798, P2_U6799, P2_U6800, P2_U6801, P2_U6802, P2_U6803, P2_U6804, P2_U6805, P2_U6806, P2_U6807, P2_U6808, P2_U6809, P2_U6810, P2_U6811, P2_U6812, P2_U6813, P2_U6814, P2_U6815, P2_U6816, P2_U6817, P2_U6818, P2_U6819, P2_U6820, P2_U6821, P2_U6822, P2_U6823, P2_U6824, P2_U6825, P2_U6826, P2_U6827, P2_U6828, P2_U6829, P2_U6830, P2_U6831, P2_U6832, P2_U6833, P2_U6834, P2_U6835, P2_U6836, P2_U6837, P2_U6838, P2_U6839, P2_U6840, P2_U6841, P2_U6842, P2_U6843, P2_U6844, P2_U6845, P2_U6846, P2_U6847, P2_U6848, P2_U6849, P2_U6850, P2_U6851, P2_U6852, P2_U6853, P2_U6854, P2_U6855, P2_U6856, P2_U6857, P2_U6858, P2_U6859, P2_U6860, P2_U6861, P2_U6862, P2_U6863, P2_U6864, P2_U6865, P2_U6866, P2_U6867, P2_U6868, P2_U6869, P2_U6870, P2_U6871, P2_U6872, P2_U6873, P2_U6874, P2_U6875, P2_U6876, P2_U6877, P2_U6878, P2_U6879, P2_U6880, P2_U6881, P2_U6882, P2_U6883, P2_U6884, P2_U6885, P2_U6886, P2_U6887, P2_U6888, P2_U6889, P2_U6890, P2_U6891, P2_U6892, P2_U6893, P2_U6894, P2_U6895, P2_U6896, P2_U6897, P2_U6898, P2_U6899, P2_U6900, P2_U6901, P2_U6902, P2_U6903, P2_U6904, P2_U6905, P2_U6906, P2_U6907, P2_U6908, P2_U6909, P2_U6910, P2_U6911, P2_U6912, P2_U6913, P2_U6914, P2_U6915, P2_U6916, P2_U6917, P2_U6918, P2_U6919, P2_U6920, P2_U6921, P2_U6922, P2_U6923, P2_U6924, P2_U6925, P2_U6926, P2_U6927, P2_U6928, P2_U6929, P2_U6930, P2_U6931, P2_U6932, P2_U6933, P2_U6934, P2_U6935, P2_U6936, P2_U6937, P2_U6938, P2_U6939, P2_U6940, P2_U6941, P2_U6942, P2_U6943, P2_U6944, P2_U6945, P2_U6946, P2_U6947, P2_U6948, P2_U6949, P2_U6950, P2_U6951, P2_U6952, P2_U6953, P2_U6954, P2_U6955, P2_U6956, P2_U6957, P2_U6958, P2_U6959, P2_U6960, P2_U6961, P2_U6962, P2_U6963, P2_U6964, P2_U6965, P2_U6966, P2_U6967, P2_U6968, P2_U6969, P2_U6970, P2_U6971, P2_U6972, P2_U6973, P2_U6974, P2_U6975, P2_U6976, P2_U6977, P2_U6978, P2_U6979, P2_U6980, P2_U6981, P2_U6982, P2_U6983, P2_U6984, P2_U6985, P2_U6986, P2_U6987, P2_U6988, P2_U6989, P2_U6990, P2_U6991, P2_U6992, P2_U6993, P2_U6994, P2_U6995, P2_U6996, P2_U6997, P2_U6998, P2_U6999, P2_U7000, P2_U7001, P2_U7002, P2_U7003, P2_U7004, P2_U7005, P2_U7006, P2_U7007, P2_U7008, P2_U7009, P2_U7010, P2_U7011, P2_U7012, P2_U7013, P2_U7014, P2_U7015, P2_U7016, P2_U7017, P2_U7018, P2_U7019, P2_U7020, P2_U7021, P2_U7022, P2_U7023, P2_U7024, P2_U7025, P2_U7026, P2_U7027, P2_U7028, P2_U7029, P2_U7030, P2_U7031, P2_U7032, P2_U7033, P2_U7034, P2_U7035, P2_U7036, P2_U7037, P2_U7038, P2_U7039, P2_U7040, P2_U7041, P2_U7042, P2_U7043, P2_U7044, P2_U7045, P2_U7046, P2_U7047, P2_U7048, P2_U7049, P2_U7050, P2_U7051, P2_U7052, P2_U7053, P2_U7054, P2_U7055, P2_U7056, P2_U7057, P2_U7058, P2_U7059, P2_U7060, P2_U7061, P2_U7062, P2_U7063, P2_U7064, P2_U7065, P2_U7066, P2_U7067, P2_U7068, P2_U7069, P2_U7070, P2_U7071, P2_U7072, P2_U7073, P2_U7074, P2_U7075, P2_U7076, P2_U7077, P2_U7078, P2_U7079, P2_U7080, P2_U7081, P2_U7082, P2_U7083, P2_U7084, P2_U7085, P2_U7086, P2_U7087, P2_U7088, P2_U7089, P2_U7090, P2_U7091, P2_U7092, P2_U7093, P2_U7094, P2_U7095, P2_U7096, P2_U7097, P2_U7098, P2_U7099, P2_U7100, P2_U7101, P2_U7102, P2_U7103, P2_U7104, P2_U7105, P2_U7106, P2_U7107, P2_U7108, P2_U7109, P2_U7110, P2_U7111, P2_U7112, P2_U7113, P2_U7114, P2_U7115, P2_U7116, P2_U7117, P2_U7118, P2_U7119, P2_U7120, P2_U7121, P2_U7122, P2_U7123, P2_U7124, P2_U7125, P2_U7126, P2_U7127, P2_U7128, P2_U7129, P2_U7130, P2_U7131, P2_U7132, P2_U7133, P2_U7134, P2_U7135, P2_U7136, P2_U7137, P2_U7138, P2_U7139, P2_U7140, P2_U7141, P2_U7142, P2_U7143, P2_U7144, P2_U7145, P2_U7146, P2_U7147, P2_U7148, P2_U7149, P2_U7150, P2_U7151, P2_U7152, P2_U7153, P2_U7154, P2_U7155, P2_U7156, P2_U7157, P2_U7158, P2_U7159, P2_U7160, P2_U7161, P2_U7162, P2_U7163, P2_U7164, P2_U7165, P2_U7166, P2_U7167, P2_U7168, P2_U7169, P2_U7170, P2_U7171, P2_U7172, P2_U7173, P2_U7174, P2_U7175, P2_U7176, P2_U7177, P2_U7178, P2_U7179, P2_U7180, P2_U7181, P2_U7182, P2_U7183, P2_U7184, P2_U7185, P2_U7186, P2_U7187, P2_U7188, P2_U7189, P2_U7190, P2_U7191, P2_U7192, P2_U7193, P2_U7194, P2_U7195, P2_U7196, P2_U7197, P2_U7198, P2_U7199, P2_U7200, P2_U7201, P2_U7202, P2_U7203, P2_U7204, P2_U7205, P2_U7206, P2_U7207, P2_U7208, P2_U7209, P2_U7210, P2_U7211, P2_U7212, P2_U7213, P2_U7214, P2_U7215, P2_U7216, P2_U7217, P2_U7218, P2_U7219, P2_U7220, P2_U7221, P2_U7222, P2_U7223, P2_U7224, P2_U7225, P2_U7226, P2_U7227, P2_U7228, P2_U7229, P2_U7230, P2_U7231, P2_U7232, P2_U7233, P2_U7234, P2_U7235, P2_U7236, P2_U7237, P2_U7238, P2_U7239, P2_U7240, P2_U7241, P2_U7242, P2_U7243, P2_U7244, P2_U7245, P2_U7246, P2_U7247, P2_U7248, P2_U7249, P2_U7250, P2_U7251, P2_U7252, P2_U7253, P2_U7254, P2_U7255, P2_U7256, P2_U7257, P2_U7258, P2_U7259, P2_U7260, P2_U7261, P2_U7262, P2_U7263, P2_U7264, P2_U7265, P2_U7266, P2_U7267, P2_U7268, P2_U7269, P2_U7270, P2_U7271, P2_U7272, P2_U7273, P2_U7274, P2_U7275, P2_U7276, P2_U7277, P2_U7278, P2_U7279, P2_U7280, P2_U7281, P2_U7282, P2_U7283, P2_U7284, P2_U7285, P2_U7286, P2_U7287, P2_U7288, P2_U7289, P2_U7290, P2_U7291, P2_U7292, P2_U7293, P2_U7294, P2_U7295, P2_U7296, P2_U7297, P2_U7298, P2_U7299, P2_U7300, P2_U7301, P2_U7302, P2_U7303, P2_U7304, P2_U7305, P2_U7306, P2_U7307, P2_U7308, P2_U7309, P2_U7310, P2_U7311, P2_U7312, P2_U7313, P2_U7314, P2_U7315, P2_U7316, P2_U7317, P2_U7318, P2_U7319, P2_U7320, P2_U7321, P2_U7322, P2_U7323, P2_U7324, P2_U7325, P2_U7326, P2_U7327, P2_U7328, P2_U7329, P2_U7330, P2_U7331, P2_U7332, P2_U7333, P2_U7334, P2_U7335, P2_U7336, P2_U7337, P2_U7338, P2_U7339, P2_U7340, P2_U7341, P2_U7342, P2_U7343, P2_U7344, P2_U7345, P2_U7346, P2_U7347, P2_U7348, P2_U7349, P2_U7350, P2_U7351, P2_U7352, P2_U7353, P2_U7354, P2_U7355, P2_U7356, P2_U7357, P2_U7358, P2_U7359, P2_U7360, P2_U7361, P2_U7362, P2_U7363, P2_U7364, P2_U7365, P2_U7366, P2_U7367, P2_U7368, P2_U7369, P2_U7370, P2_U7371, P2_U7372, P2_U7373, P2_U7374, P2_U7375, P2_U7376, P2_U7377, P2_U7378, P2_U7379, P2_U7380, P2_U7381, P2_U7382, P2_U7383, P2_U7384, P2_U7385, P2_U7386, P2_U7387, P2_U7388, P2_U7389, P2_U7390, P2_U7391, P2_U7392, P2_U7393, P2_U7394, P2_U7395, P2_U7396, P2_U7397, P2_U7398, P2_U7399, P2_U7400, P2_U7401, P2_U7402, P2_U7403, P2_U7404, P2_U7405, P2_U7406, P2_U7407, P2_U7408, P2_U7409, P2_U7410, P2_U7411, P2_U7412, P2_U7413, P2_U7414, P2_U7415, P2_U7416, P2_U7417, P2_U7418, P2_U7419, P2_U7420, P2_U7421, P2_U7422, P2_U7423, P2_U7424, P2_U7425, P2_U7426, P2_U7427, P2_U7428, P2_U7429, P2_U7430, P2_U7431, P2_U7432, P2_U7433, P2_U7434, P2_U7435, P2_U7436, P2_U7437, P2_U7438, P2_U7439, P2_U7440, P2_U7441, P2_U7442, P2_U7443, P2_U7444, P2_U7445, P2_U7446, P2_U7447, P2_U7448, P2_U7449, P2_U7450, P2_U7451, P2_U7452, P2_U7453, P2_U7454, P2_U7455, P2_U7456, P2_U7457, P2_U7458, P2_U7459, P2_U7460, P2_U7461, P2_U7462, P2_U7463, P2_U7464, P2_U7465, P2_U7466, P2_U7467, P2_U7468, P2_U7469, P2_U7470, P2_U7471, P2_U7472, P2_U7473, P2_U7474, P2_U7475, P2_U7476, P2_U7477, P2_U7478, P2_U7479, P2_U7480, P2_U7481, P2_U7482, P2_U7483, P2_U7484, P2_U7485, P2_U7486, P2_U7487, P2_U7488, P2_U7489, P2_U7490, P2_U7491, P2_U7492, P2_U7493, P2_U7494, P2_U7495, P2_U7496, P2_U7497, P2_U7498, P2_U7499, P2_U7500, P2_U7501, P2_U7502, P2_U7503, P2_U7504, P2_U7505, P2_U7506, P2_U7507, P2_U7508, P2_U7509, P2_U7510, P2_U7511, P2_U7512, P2_U7513, P2_U7514, P2_U7515, P2_U7516, P2_U7517, P2_U7518, P2_U7519, P2_U7520, P2_U7521, P2_U7522, P2_U7523, P2_U7524, P2_U7525, P2_U7526, P2_U7527, P2_U7528, P2_U7529, P2_U7530, P2_U7531, P2_U7532, P2_U7533, P2_U7534, P2_U7535, P2_U7536, P2_U7537, P2_U7538, P2_U7539, P2_U7540, P2_U7541, P2_U7542, P2_U7543, P2_U7544, P2_U7545, P2_U7546, P2_U7547, P2_U7548, P2_U7549, P2_U7550, P2_U7551, P2_U7552, P2_U7553, P2_U7554, P2_U7555, P2_U7556, P2_U7557, P2_U7558, P2_U7559, P2_U7560, P2_U7561, P2_U7562, P2_U7563, P2_U7564, P2_U7565, P2_U7566, P2_U7567, P2_U7568, P2_U7569, P2_U7570, P2_U7571, P2_U7572, P2_U7573, P2_U7574, P2_U7575, P2_U7576, P2_U7577, P2_U7578, P2_U7579, P2_U7580, P2_U7581, P2_U7582, P2_U7583, P2_U7584, P2_U7585, P2_U7586, P2_U7587, P2_U7588, P2_U7589, P2_U7590, P2_U7591, P2_U7592, P2_U7593, P2_U7594, P2_U7595, P2_U7596, P2_U7597, P2_U7598, P2_U7599, P2_U7600, P2_U7601, P2_U7602, P2_U7603, P2_U7604, P2_U7605, P2_U7606, P2_U7607, P2_U7608, P2_U7609, P2_U7610, P2_U7611, P2_U7612, P2_U7613, P2_U7614, P2_U7615, P2_U7616, P2_U7617, P2_U7618, P2_U7619, P2_U7620, P2_U7621, P2_U7622, P2_U7623, P2_U7624, P2_U7625, P2_U7626, P2_U7627, P2_U7628, P2_U7629, P2_U7630, P2_U7631, P2_U7632, P2_U7633, P2_U7634, P2_U7635, P2_U7636, P2_U7637, P2_U7638, P2_U7639, P2_U7640, P2_U7641, P2_U7642, P2_U7643, P2_U7644, P2_U7645, P2_U7646, P2_U7647, P2_U7648, P2_U7649, P2_U7650, P2_U7651, P2_U7652, P2_U7653, P2_U7654, P2_U7655, P2_U7656, P2_U7657, P2_U7658, P2_U7659, P2_U7660, P2_U7661, P2_U7662, P2_U7663, P2_U7664, P2_U7665, P2_U7666, P2_U7667, P2_U7668, P2_U7669, P2_U7670, P2_U7671, P2_U7672, P2_U7673, P2_U7674, P2_U7675, P2_U7676, P2_U7677, P2_U7678, P2_U7679, P2_U7680, P2_U7681, P2_U7682, P2_U7683, P2_U7684, P2_U7685, P2_U7686, P2_U7687, P2_U7688, P2_U7689, P2_U7690, P2_U7691, P2_U7692, P2_U7693, P2_U7694, P2_U7695, P2_U7696, P2_U7697, P2_U7698, P2_U7699, P2_U7700, P2_U7701, P2_U7702, P2_U7703, P2_U7704, P2_U7705, P2_U7706, P2_U7707, P2_U7708, P2_U7709, P2_U7710, P2_U7711, P2_U7712, P2_U7713, P2_U7714, P2_U7715, P2_U7716, P2_U7717, P2_U7718, P2_U7719, P2_U7720, P2_U7721, P2_U7722, P2_U7723, P2_U7724, P2_U7725, P2_U7726, P2_U7727, P2_U7728, P2_U7729, P2_U7730, P2_U7731, P2_U7732, P2_U7733, P2_U7734, P2_U7735, P2_U7736, P2_U7737, P2_U7738, P2_U7739, P2_U7740, P2_U7741, P2_U7742, P2_U7743, P2_U7744, P2_U7745, P2_U7746, P2_U7747, P2_U7748, P2_U7749, P2_U7750, P2_U7751, P2_U7752, P2_U7753, P2_U7754, P2_U7755, P2_U7756, P2_U7757, P2_U7758, P2_U7759, P2_U7760, P2_U7761, P2_U7762, P2_U7763, P2_U7764, P2_U7765, P2_U7766, P2_U7767, P2_U7768, P2_U7769, P2_U7770, P2_U7771, P2_U7772, P2_U7773, P2_U7774, P2_U7775, P2_U7776, P2_U7777, P2_U7778, P2_U7779, P2_U7780, P2_U7781, P2_U7782, P2_U7783, P2_U7784, P2_U7785, P2_U7786, P2_U7787, P2_U7788, P2_U7789, P2_U7790, P2_U7791, P2_U7792, P2_U7793, P2_U7794, P2_U7795, P2_U7796, P2_U7797, P2_U7798, P2_U7799, P2_U7800, P2_U7801, P2_U7802, P2_U7803, P2_U7804, P2_U7805, P2_U7806, P2_U7807, P2_U7808, P2_U7809, P2_U7810, P2_U7811, P2_U7812, P2_U7813, P2_U7814, P2_U7815, P2_U7816, P2_U7817, P2_U7818, P2_U7819, P2_U7820, P2_U7821, P2_U7822, P2_U7823, P2_U7824, P2_U7825, P2_U7826, P2_U7827, P2_U7828, P2_U7829, P2_U7830, P2_U7831, P2_U7832, P2_U7833, P2_U7834, P2_U7835, P2_U7836, P2_U7837, P2_U7838, P2_U7839, P2_U7840, P2_U7841, P2_U7842, P2_U7843, P2_U7844, P2_U7845, P2_U7846, P2_U7847, P2_U7848, P2_U7849, P2_U7850, P2_U7851, P2_U7852, P2_U7853, P2_U7854, P2_U7855, P2_U7856, P2_U7857, P2_U7858, P2_U7859, P2_U7860, P2_U7861, P2_U7862, P2_U7863, P2_U7864, P2_U7865, P2_U7866, P2_U7867, P2_U7868, P2_U7869, P2_U7870, P2_U7871, P2_U7872, P2_U7873, P2_U7874, P2_U7875, P2_U7876, P2_U7877, P2_U7878, P2_U7879, P2_U7880, P2_U7881, P2_U7882, P2_U7883, P2_U7884, P2_U7885, P2_U7886, P2_U7887, P2_U7888, P2_U7889, P2_U7890, P2_U7891, P2_U7892, P2_U7893, P2_U7894, P2_U7895, P2_U7896, P2_U7897, P2_U7898, P2_U7899, P2_U7900, P2_U7901, P2_U7902, P2_U7903, P2_U7904, P2_U7905, P2_U7906, P2_U7907, P2_U7908, P2_U7909, P2_U7910, P2_U7911, P2_U7912, P2_U7913, P2_U7914, P2_U7915, P2_U7916, P2_U7917, P2_U7918, P2_U7919, P2_U7920, P2_U7921, P2_U7922, P2_U7923, P2_U7924, P2_U7925, P2_U7926, P2_U7927, P2_U7928, P2_U7929, P2_U7930, P2_U7931, P2_U7932, P2_U7933, P2_U7934, P2_U7935, P2_U7936, P2_U7937, P2_U7938, P2_U7939, P2_U7940, P2_U7941, P2_U7942, P2_U7943, P2_U7944, P2_U7945, P2_U7946, P2_U7947, P2_U7948, P2_U7949, P2_U7950, P2_U7951, P2_U7952, P2_U7953, P2_U7954, P2_U7955, P2_U7956, P2_U7957, P2_U7958, P2_U7959, P2_U7960, P2_U7961, P2_U7962, P2_U7963, P2_U7964, P2_U7965, P2_U7966, P2_U7967, P2_U7968, P2_U7969, P2_U7970, P2_U7971, P2_U7972, P2_U7973, P2_U7974, P2_U7975, P2_U7976, P2_U7977, P2_U7978, P2_U7979, P2_U7980, P2_U7981, P2_U7982, P2_U7983, P2_U7984, P2_U7985, P2_U7986, P2_U7987, P2_U7988, P2_U7989, P2_U7990, P2_U7991, P2_U7992, P2_U7993, P2_U7994, P2_U7995, P2_U7996, P2_U7997, P2_U7998, P2_U7999, P2_U8000, P2_U8001, P2_U8002, P2_U8003, P2_U8004, P2_U8005, P2_U8006, P2_U8007, P2_U8008, P2_U8009, P2_U8010, P2_U8011, P2_U8012, P2_U8013, P2_U8014, P2_U8015, P2_U8016, P2_U8017, P2_U8018, P2_U8019, P2_U8020, P2_U8021, P2_U8022, P2_U8023, P2_U8024, P2_U8025, P2_U8026, P2_U8027, P2_U8028, P2_U8029, P2_U8030, P2_U8031, P2_U8032, P2_U8033, P2_U8034, P2_U8035, P2_U8036, P2_U8037, P2_U8038, P2_U8039, P2_U8040, P2_U8041, P2_U8042, P2_U8043, P2_U8044, P2_U8045, P2_U8046, P2_U8047, P2_U8048, P2_U8049, P2_U8050, P2_U8051, P2_U8052, P2_U8053, P2_U8054, P2_U8055, P2_U8056, P2_U8057, P2_U8058, P2_U8059, P2_U8060, P2_U8061, P2_U8062, P2_U8063, P2_U8064, P2_U8065, P2_U8066, P2_U8067, P2_U8068, P2_U8069, P2_U8070, P2_U8071, P2_U8072, P2_U8073, P2_U8074, P2_U8075, P2_U8076, P2_U8077, P2_U8078, P2_U8079, P2_U8080, P2_U8081, P2_U8082, P2_U8083, P2_U8084, P2_U8085, P2_U8086, P2_U8087, P2_U8088, P2_U8089, P2_U8090, P2_U8091, P2_U8092, P2_U8093, P2_U8094, P2_U8095, P2_U8096, P2_U8097, P2_U8098, P2_U8099, P2_U8100, P2_U8101, P2_U8102, P2_U8103, P2_U8104, P2_U8105, P2_U8106, P2_U8107, P2_U8108, P2_U8109, P2_U8110, P2_U8111, P2_U8112, P2_U8113, P2_U8114, P2_U8115, P2_U8116, P2_U8117, P2_U8118, P2_U8119, P2_U8120, P2_U8121, P2_U8122, P2_U8123, P2_U8124, P2_U8125, P2_U8126, P2_U8127, P2_U8128, P2_U8129, P2_U8130, P2_U8131, P2_U8132, P2_U8133, P2_U8134, P2_U8135, P2_U8136, P2_U8137, P2_U8138, P2_U8139, P2_U8140, P2_U8141, P2_U8142, P2_U8143, P2_U8144, P2_U8145, P2_U8146, P2_U8147, P2_U8148, P2_U8149, P2_U8150, P2_U8151, P2_U8152, P2_U8153, P2_U8154, P2_U8155, P2_U8156, P2_U8157, P2_U8158, P2_U8159, P2_U8160, P2_U8161, P2_U8162, P2_U8163, P2_U8164, P2_U8165, P2_U8166, P2_U8167, P2_U8168, P2_U8169, P2_U8170, P2_U8171, P2_U8172, P2_U8173, P2_U8174, P2_U8175, P2_U8176, P2_U8177, P2_U8178, P2_U8179, P2_U8180, P2_U8181, P2_U8182, P2_U8183, P2_U8184, P2_U8185, P2_U8186, P2_U8187, P2_U8188, P2_U8189, P2_U8190, P2_U8191, P2_U8192, P2_U8193, P2_U8194, P2_U8195, P2_U8196, P2_U8197, P2_U8198, P2_U8199, P2_U8200, P2_U8201, P2_U8202, P2_U8203, P2_U8204, P2_U8205, P2_U8206, P2_U8207, P2_U8208, P2_U8209, P2_U8210, P2_U8211, P2_U8212, P2_U8213, P2_U8214, P2_U8215, P2_U8216, P2_U8217, P2_U8218, P2_U8219, P2_U8220, P2_U8221, P2_U8222, P2_U8223, P2_U8224, P2_U8225, P2_U8226, P2_U8227, P2_U8228, P2_U8229, P2_U8230, P2_U8231, P2_U8232, P2_U8233, P2_U8234, P2_U8235, P2_U8236, P2_U8237, P2_U8238, P2_U8239, P2_U8240, P2_U8241, P2_U8242, P2_U8243, P2_U8244, P2_U8245, P2_U8246, P2_U8247, P2_U8248, P2_U8249, P2_U8250, P2_U8251, P2_U8252, P2_U8253, P2_U8254, P2_U8255, P2_U8256, P2_U8257, P2_U8258, P2_U8259, P2_U8260, P2_U8261, P2_U8262, P2_U8263, P2_U8264, P2_U8265, P2_U8266, P2_U8267, P2_U8268, P2_U8269, P2_U8270, P2_U8271, P2_U8272, P2_U8273, P2_U8274, P2_U8275, P2_U8276, P2_U8277, P2_U8278, P2_U8279, P2_U8280, P2_U8281, P2_U8282, P2_U8283, P2_U8284, P2_U8285, P2_U8286, P2_U8287, P2_U8288, P2_U8289, P2_U8290, P2_U8291, P2_U8292, P2_U8293, P2_U8294, P2_U8295, P2_U8296, P2_U8297, P2_U8298, P2_U8299, P2_U8300, P2_U8301, P2_U8302, P2_U8303, P2_U8304, P2_U8305, P2_U8306, P2_U8307, P2_U8308, P2_U8309, P2_U8310, P2_U8311, P2_U8312, P2_U8313, P2_U8314, P2_U8315, P2_U8316, P2_U8317, P2_U8318, P2_U8319, P2_U8320, P2_U8321, P2_U8322, P2_U8323, P2_U8324, P2_U8325, P2_U8326, P2_U8327, P2_U8328, P2_U8329, P2_U8330, P2_U8331, P2_U8332, P2_U8333, P2_U8334, P2_U8335, P2_U8336, P2_U8337, P2_U8338, P2_U8339, P2_U8340, P2_U8341, P2_U8342, P2_U8343, P2_U8344, P2_U8345, P2_U8346, P2_U8347, P2_U8348, P2_U8349, P2_U8350, P2_U8351, P2_U8352, P2_U8353, P2_U8354, P2_U8355, P2_U8356, P2_U8357, P2_U8358, P2_U8359, P2_U8360, P2_U8361, P2_U8362, P2_U8363, P2_U8364, P2_U8365, P2_U8366, P2_U8367, P2_U8368, P2_U8369, P2_U8370, P2_U8371, P2_U8372, P2_U8373, P2_U8374, P2_U8375, P2_U8376, P2_U8377, P2_U8378, P2_U8379, P2_U8380, P2_U8381, P2_U8382, P2_U8383, P2_U8384, P2_U8385, P2_U8386, P2_U8387, P2_U8388, P2_U8389, P2_U8390, P2_U8391, P2_U8392, P2_U8393, P2_U8394, P2_U8395, P2_U8396, P2_U8397, P2_U8398, P2_U8399, P2_U8400, P2_U8401, P2_U8402, P2_U8403, P2_U8404, P2_U8405, P2_U8406, P2_U8407, P2_U8408, P2_U8409, P2_U8410, P2_U8411, P2_U8412, P2_U8413, P2_U8414, P2_U8415, P2_U8416, P2_U8417, P2_U8418, P2_U8419, P2_U8420, P2_U8421, P2_U8422, P2_U8423, P2_U8424, P2_U8425, P2_U8426, P2_U8427, P2_U8428, P2_U8429, P2_U8430, P2_U8431, P2_U8432, P2_U8433, P2_U8434, P1_U2352, P1_U2353, P1_U2354, P1_U2355, P1_U2356, P1_U2357, P1_U2358, P1_U2359, P1_U2360, P1_U2361, P1_U2362, P1_U2363, P1_U2364, P1_U2365, P1_U2366, P1_U2367, P1_U2368, P1_U2369, P1_U2370, P1_U2371, P1_U2372, P1_U2373, P1_U2374, P1_U2375, P1_U2376, P1_U2377, P1_U2378, P1_U2379, P1_U2380, P1_U2381, P1_U2382, P1_U2383, P1_U2384, P1_U2385, P1_U2386, P1_U2387, P1_U2388, P1_U2389, P1_U2390, P1_U2391, P1_U2392, P1_U2393, P1_U2394, P1_U2395, P1_U2396, P1_U2397, P1_U2398, P1_U2399, P1_U2400, P1_U2401, P1_U2402, P1_U2403, P1_U2404, P1_U2405, P1_U2406, P1_U2407, P1_U2408, P1_U2409, P1_U2410, P1_U2411, P1_U2412, P1_U2413, P1_U2414, P1_U2415, P1_U2416, P1_U2417, P1_U2418, P1_U2419, P1_U2420, P1_U2421, P1_U2422, P1_U2423, P1_U2424, P1_U2425, P1_U2426, P1_U2427, P1_U2428, P1_U2429, P1_U2430, P1_U2431, P1_U2432, P1_U2433, P1_U2434, P1_U2435, P1_U2436, P1_U2437, P1_U2438, P1_U2439, P1_U2440, P1_U2441, P1_U2442, P1_U2443, P1_U2444, P1_U2445, P1_U2446, P1_U2447, P1_U2448, P1_U2449, P1_U2450, P1_U2451, P1_U2452, P1_U2453, P1_U2454, P1_U2455, P1_U2456, P1_U2457, P1_U2458, P1_U2459, P1_U2460, P1_U2461, P1_U2462, P1_U2463, P1_U2464, P1_U2465, P1_U2466, P1_U2467, P1_U2468, P1_U2469, P1_U2470, P1_U2471, P1_U2472, P1_U2473, P1_U2474, P1_U2475, P1_U2476, P1_U2477, P1_U2478, P1_U2479, P1_U2480, P1_U2481, P1_U2482, P1_U2483, P1_U2484, P1_U2485, P1_U2486, P1_U2487, P1_U2488, P1_U2489, P1_U2490, P1_U2491, P1_U2492, P1_U2493, P1_U2494, P1_U2495, P1_U2496, P1_U2497, P1_U2498, P1_U2499, P1_U2500, P1_U2501, P1_U2502, P1_U2503, P1_U2504, P1_U2505, P1_U2506, P1_U2507, P1_U2508, P1_U2509, P1_U2510, P1_U2511, P1_U2512, P1_U2513, P1_U2514, P1_U2515, P1_U2516, P1_U2517, P1_U2518, P1_U2519, P1_U2520, P1_U2521, P1_U2522, P1_U2523, P1_U2524, P1_U2525, P1_U2526, P1_U2527, P1_U2528, P1_U2529, P1_U2530, P1_U2531, P1_U2532, P1_U2533, P1_U2534, P1_U2535, P1_U2536, P1_U2537, P1_U2538, P1_U2539, P1_U2540, P1_U2541, P1_U2542, P1_U2543, P1_U2544, P1_U2545, P1_U2546, P1_U2547, P1_U2548, P1_U2549, P1_U2550, P1_U2551, P1_U2552, P1_U2553, P1_U2554, P1_U2555, P1_U2556, P1_U2557, P1_U2558, P1_U2559, P1_U2560, P1_U2561, P1_U2562, P1_U2563, P1_U2564, P1_U2565, P1_U2566, P1_U2567, P1_U2568, P1_U2569, P1_U2570, P1_U2571, P1_U2572, P1_U2573, P1_U2574, P1_U2575, P1_U2576, P1_U2577, P1_U2578, P1_U2579, P1_U2580, P1_U2581, P1_U2582, P1_U2583, P1_U2584, P1_U2585, P1_U2586, P1_U2587, P1_U2588, P1_U2589, P1_U2590, P1_U2591, P1_U2592, P1_U2593, P1_U2594, P1_U2595, P1_U2596, P1_U2597, P1_U2598, P1_U2599, P1_U2600, P1_U2601, P1_U2602, P1_U2603, P1_U2604, P1_U2605, P1_U2606, P1_U2607, P1_U2608, P1_U2609, P1_U2610, P1_U2611, P1_U2612, P1_U2613, P1_U2614, P1_U2615, P1_U2616, P1_U2617, P1_U2618, P1_U2620, P1_U2621, P1_U2622, P1_U2623, P1_U2624, P1_U2625, P1_U2626, P1_U2627, P1_U2628, P1_U2629, P1_U2630, P1_U2631, P1_U2632, P1_U2633, P1_U2634, P1_U2635, P1_U2636, P1_U2637, P1_U2638, P1_U2639, P1_U2640, P1_U2641, P1_U2642, P1_U2643, P1_U2644, P1_U2645, P1_U2646, P1_U2647, P1_U2648, P1_U2649, P1_U2650, P1_U2651, P1_U2652, P1_U2653, P1_U2654, P1_U2655, P1_U2656, P1_U2657, P1_U2658, P1_U2659, P1_U2660, P1_U2661, P1_U2662, P1_U2663, P1_U2664, P1_U2665, P1_U2666, P1_U2667, P1_U2668, P1_U2669, P1_U2670, P1_U2671, P1_U2672, P1_U2673, P1_U2674, P1_U2675, P1_U2676, P1_U2677, P1_U2678, P1_U2679, P1_U2680, P1_U2681, P1_U2682, P1_U2683, P1_U2684, P1_U2685, P1_U2686, P1_U2687, P1_U2688, P1_U2689, P1_U2690, P1_U2691, P1_U2692, P1_U2693, P1_U2694, P1_U2695, P1_U2696, P1_U2697, P1_U2698, P1_U2699, P1_U2700, P1_U2701, P1_U2702, P1_U2703, P1_U2704, P1_U2705, P1_U2706, P1_U2707, P1_U2708, P1_U2709, P1_U2710, P1_U2711, P1_U2712, P1_U2713, P1_U2714, P1_U2715, P1_U2716, P1_U2717, P1_U2718, P1_U2719, P1_U2720, P1_U2721, P1_U2722, P1_U2723, P1_U2724, P1_U2725, P1_U2726, P1_U2727, P1_U2728, P1_U2729, P1_U2730, P1_U2731, P1_U2732, P1_U2733, P1_U2734, P1_U2735, P1_U2736, P1_U2737, P1_U2738, P1_U2739, P1_U2740, P1_U2741, P1_U2742, P1_U2743, P1_U2744, P1_U2745, P1_U2746, P1_U2747, P1_U2748, P1_U2749, P1_U2750, P1_U2751, P1_U2752, P1_U2753, P1_U2754, P1_U2755, P1_U2756, P1_U2757, P1_U2758, P1_U2759, P1_U2760, P1_U2761, P1_U2762, P1_U2763, P1_U2764, P1_U2765, P1_U2766, P1_U2767, P1_U2768, P1_U2769, P1_U2770, P1_U2771, P1_U2772, P1_U2773, P1_U2774, P1_U2775, P1_U2776, P1_U2777, P1_U2778, P1_U2779, P1_U2780, P1_U2781, P1_U2782, P1_U2783, P1_U2784, P1_U2785, P1_U2786, P1_U2787, P1_U2788, P1_U2789, P1_U2790, P1_U2791, P1_U2792, P1_U2793, P1_U2794, P1_U2795, P1_U2796, P1_U2797, P1_U2798, P1_U2799, P1_U2800, P1_U3227, P1_U3228, P1_U3229, P1_U3230, P1_U3231, P1_U3232, P1_U3233, P1_U3234, P1_U3235, P1_U3236, P1_U3237, P1_U3238, P1_U3239, P1_U3240, P1_U3241, P1_U3242, P1_U3243, P1_U3244, P1_U3245, P1_U3246, P1_U3247, P1_U3248, P1_U3249, P1_U3250, P1_U3251, P1_U3252, P1_U3253, P1_U3254, P1_U3255, P1_U3256, P1_U3257, P1_U3258, P1_U3259, P1_U3260, P1_U3261, P1_U3262, P1_U3263, P1_U3264, P1_U3265, P1_U3266, P1_U3267, P1_U3268, P1_U3269, P1_U3270, P1_U3271, P1_U3272, P1_U3273, P1_U3274, P1_U3275, P1_U3276, P1_U3277, P1_U3278, P1_U3279, P1_U3280, P1_U3281, P1_U3282, P1_U3283, P1_U3284, P1_U3285, P1_U3286, P1_U3287, P1_U3288, P1_U3289, P1_U3290, P1_U3291, P1_U3292, P1_U3293, P1_U3294, P1_U3295, P1_U3296, P1_U3297, P1_U3298, P1_U3299, P1_U3300, P1_U3301, P1_U3302, P1_U3303, P1_U3304, P1_U3305, P1_U3306, P1_U3307, P1_U3308, P1_U3309, P1_U3310, P1_U3311, P1_U3312, P1_U3313, P1_U3314, P1_U3315, P1_U3316, P1_U3317, P1_U3318, P1_U3319, P1_U3320, P1_U3321, P1_U3322, P1_U3323, P1_U3324, P1_U3325, P1_U3326, P1_U3327, P1_U3328, P1_U3329, P1_U3330, P1_U3331, P1_U3332, P1_U3333, P1_U3334, P1_U3335, P1_U3336, P1_U3337, P1_U3338, P1_U3339, P1_U3340, P1_U3341, P1_U3342, P1_U3343, P1_U3344, P1_U3345, P1_U3346, P1_U3347, P1_U3348, P1_U3349, P1_U3350, P1_U3351, P1_U3352, P1_U3353, P1_U3354, P1_U3355, P1_U3356, P1_U3357, P1_U3358, P1_U3359, P1_U3360, P1_U3361, P1_U3362, P1_U3363, P1_U3364, P1_U3365, P1_U3366, P1_U3367, P1_U3368, P1_U3369, P1_U3370, P1_U3371, P1_U3372, P1_U3373, P1_U3374, P1_U3375, P1_U3376, P1_U3377, P1_U3378, P1_U3379, P1_U3380, P1_U3381, P1_U3382, P1_U3383, P1_U3384, P1_U3385, P1_U3386, P1_U3387, P1_U3388, P1_U3389, P1_U3390, P1_U3391, P1_U3392, P1_U3393, P1_U3394, P1_U3395, P1_U3396, P1_U3397, P1_U3398, P1_U3399, P1_U3400, P1_U3401, P1_U3402, P1_U3403, P1_U3404, P1_U3405, P1_U3406, P1_U3407, P1_U3408, P1_U3409, P1_U3410, P1_U3411, P1_U3412, P1_U3413, P1_U3414, P1_U3415, P1_U3416, P1_U3417, P1_U3418, P1_U3419, P1_U3420, P1_U3421, P1_U3422, P1_U3423, P1_U3424, P1_U3425, P1_U3426, P1_U3427, P1_U3428, P1_U3429, P1_U3430, P1_U3431, P1_U3432, P1_U3433, P1_U3434, P1_U3435, P1_U3436, P1_U3437, P1_U3438, P1_U3439, P1_U3440, P1_U3441, P1_U3442, P1_U3443, P1_U3444, P1_U3445, P1_U3446, P1_U3447, P1_U3448, P1_U3449, P1_U3450, P1_U3451, P1_U3452, P1_U3453, P1_U3454, P1_U3455, P1_U3456, P1_U3457, P1_U3462, P1_U3463, P1_U3467, P1_U3470, P1_U3471, P1_U3479, P1_U3480, P1_U3488, P1_U3489, P1_U3490, P1_U3491, P1_U3492, P1_U3493, P1_U3494, P1_U3495, P1_U3496, P1_U3497, P1_U3498, P1_U3499, P1_U3500, P1_U3501, P1_U3502, P1_U3503, P1_U3504, P1_U3505, P1_U3506, P1_U3507, P1_U3508, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3592, P1_U3593, P1_U3594, P1_U3595, P1_U3596, P1_U3597, P1_U3598, P1_U3599, P1_U3600, P1_U3601, P1_U3602, P1_U3603, P1_U3604, P1_U3605, P1_U3606, P1_U3607, P1_U3608, P1_U3609, P1_U3610, P1_U3611, P1_U3612, P1_U3613, P1_U3614, P1_U3615, P1_U3616, P1_U3617, P1_U3618, P1_U3619, P1_U3620, P1_U3621, P1_U3622, P1_U3623, P1_U3624, P1_U3625, P1_U3626, P1_U3627, P1_U3628, P1_U3629, P1_U3630, P1_U3631, P1_U3632, P1_U3633, P1_U3634, P1_U3635, P1_U3636, P1_U3637, P1_U3638, P1_U3639, P1_U3640, P1_U3641, P1_U3642, P1_U3643, P1_U3644, P1_U3645, P1_U3646, P1_U3647, P1_U3648, P1_U3649, P1_U3650, P1_U3651, P1_U3652, P1_U3653, P1_U3654, P1_U3655, P1_U3656, P1_U3657, P1_U3658, P1_U3659, P1_U3660, P1_U3661, P1_U3662, P1_U3663, P1_U3664, P1_U3665, P1_U3666, P1_U3667, P1_U3668, P1_U3669, P1_U3670, P1_U3671, P1_U3672, P1_U3673, P1_U3674, P1_U3675, P1_U3676, P1_U3677, P1_U3678, P1_U3679, P1_U3680, P1_U3681, P1_U3682, P1_U3683, P1_U3684, P1_U3685, P1_U3686, P1_U3687, P1_U3688, P1_U3689, P1_U3690, P1_U3691, P1_U3692, P1_U3693, P1_U3694, P1_U3695, P1_U3696, P1_U3697, P1_U3698, P1_U3699, P1_U3700, P1_U3701, P1_U3702, P1_U3703, P1_U3704, P1_U3705, P1_U3706, P1_U3707, P1_U3708, P1_U3709, P1_U3710, P1_U3711, P1_U3712, P1_U3713, P1_U3714, P1_U3715, P1_U3716, P1_U3717, P1_U3718, P1_U3719, P1_U3720, P1_U3721, P1_U3722, P1_U3723, P1_U3724, P1_U3725, P1_U3726, P1_U3727, P1_U3728, P1_U3729, P1_U3730, P1_U3731, P1_U3732, P1_U3733, P1_U3734, P1_U3735, P1_U3736, P1_U3737, P1_U3738, P1_U3739, P1_U3740, P1_U3741, P1_U3742, P1_U3743, P1_U3744, P1_U3745, P1_U3746, P1_U3747, P1_U3748, P1_U3749, P1_U3750, P1_U3751, P1_U3752, P1_U3753, P1_U3754, P1_U3755, P1_U3756, P1_U3757, P1_U3758, P1_U3759, P1_U3760, P1_U3761, P1_U3762, P1_U3763, P1_U3764, P1_U3765, P1_U3766, P1_U3767, P1_U3768, P1_U3769, P1_U3770, P1_U3771, P1_U3772, P1_U3773, P1_U3774, P1_U3775, P1_U3776, P1_U3777, P1_U3778, P1_U3779, P1_U3780, P1_U3781, P1_U3782, P1_U3783, P1_U3784, P1_U3785, P1_U3786, P1_U3787, P1_U3788, P1_U3789, P1_U3790, P1_U3791, P1_U3792, P1_U3793, P1_U3794, P1_U3795, P1_U3796, P1_U3797, P1_U3798, P1_U3799, P1_U3800, P1_U3801, P1_U3802, P1_U3803, P1_U3804, P1_U3805, P1_U3806, P1_U3807, P1_U3808, P1_U3809, P1_U3810, P1_U3811, P1_U3812, P1_U3813, P1_U3814, P1_U3815, P1_U3816, P1_U3817, P1_U3818, P1_U3819, P1_U3820, P1_U3821, P1_U3822, P1_U3823, P1_U3824, P1_U3825, P1_U3826, P1_U3827, P1_U3828, P1_U3829, P1_U3830, P1_U3831, P1_U3832, P1_U3833, P1_U3834, P1_U3835, P1_U3836, P1_U3837, P1_U3838, P1_U3839, P1_U3840, P1_U3841, P1_U3842, P1_U3843, P1_U3844, P1_U3845, P1_U3846, P1_U3847, P1_U3848, P1_U3849, P1_U3850, P1_U3851, P1_U3852, P1_U3853, P1_U3854, P1_U3855, P1_U3856, P1_U3857, P1_U3858, P1_U3859, P1_U3860, P1_U3861, P1_U3862, P1_U3863, P1_U3864, P1_U3865, P1_U3866, P1_U3867, P1_U3868, P1_U3869, P1_U3870, P1_U3871, P1_U3872, P1_U3873, P1_U3874, P1_U3875, P1_U3876, P1_U3877, P1_U3878, P1_U3879, P1_U3880, P1_U3881, P1_U3882, P1_U3883, P1_U3884, P1_U3885, P1_U3886, P1_U3887, P1_U3888, P1_U3889, P1_U3890, P1_U3891, P1_U3892, P1_U3893, P1_U3894, P1_U3895, P1_U3896, P1_U3897, P1_U3898, P1_U3899, P1_U3900, P1_U3901, P1_U3902, P1_U3903, P1_U3904, P1_U3905, P1_U3906, P1_U3907, P1_U3908, P1_U3909, P1_U3910, P1_U3911, P1_U3912, P1_U3913, P1_U3914, P1_U3915, P1_U3916, P1_U3917, P1_U3918, P1_U3919, P1_U3920, P1_U3921, P1_U3922, P1_U3923, P1_U3924, P1_U3925, P1_U3926, P1_U3927, P1_U3928, P1_U3929, P1_U3930, P1_U3931, P1_U3932, P1_U3933, P1_U3934, P1_U3935, P1_U3936, P1_U3937, P1_U3938, P1_U3939, P1_U3940, P1_U3941, P1_U3942, P1_U3943, P1_U3944, P1_U3945, P1_U3946, P1_U3947, P1_U3948, P1_U3949, P1_U3950, P1_U3951, P1_U3952, P1_U3953, P1_U3954, P1_U3955, P1_U3956, P1_U3957, P1_U3958, P1_U3959, P1_U3960, P1_U3961, P1_U3962, P1_U3963, P1_U3964, P1_U3965, P1_U3966, P1_U3967, P1_U3968, P1_U3969, P1_U3970, P1_U3971, P1_U3972, P1_U3973, P1_U3974, P1_U3975, P1_U3976, P1_U3977, P1_U3978, P1_U3979, P1_U3980, P1_U3981, P1_U3982, P1_U3983, P1_U3984, P1_U3985, P1_U3986, P1_U3987, P1_U3988, P1_U3989, P1_U3990, P1_U3991, P1_U3992, P1_U3993, P1_U3994, P1_U3995, P1_U3996, P1_U3997, P1_U3998, P1_U3999, P1_U4000, P1_U4001, P1_U4002, P1_U4003, P1_U4004, P1_U4005, P1_U4006, P1_U4007, P1_U4008, P1_U4009, P1_U4010, P1_U4011, P1_U4012, P1_U4013, P1_U4014, P1_U4015, P1_U4016, P1_U4017, P1_U4018, P1_U4019, P1_U4020, P1_U4021, P1_U4022, P1_U4023, P1_U4024, P1_U4025, P1_U4026, P1_U4027, P1_U4028, P1_U4029, P1_U4030, P1_U4031, P1_U4032, P1_U4033, P1_U4034, P1_U4035, P1_U4036, P1_U4037, P1_U4038, P1_U4039, P1_U4040, P1_U4041, P1_U4042, P1_U4043, P1_U4044, P1_U4045, P1_U4046, P1_U4047, P1_U4048, P1_U4049, P1_U4050, P1_U4051, P1_U4052, P1_U4053, P1_U4054, P1_U4055, P1_U4056, P1_U4057, P1_U4058, P1_U4059, P1_U4060, P1_U4061, P1_U4062, P1_U4063, P1_U4064, P1_U4065, P1_U4066, P1_U4067, P1_U4068, P1_U4069, P1_U4070, P1_U4071, P1_U4072, P1_U4073, P1_U4074, P1_U4075, P1_U4076, P1_U4077, P1_U4078, P1_U4079, P1_U4080, P1_U4081, P1_U4082, P1_U4083, P1_U4084, P1_U4085, P1_U4086, P1_U4087, P1_U4088, P1_U4089, P1_U4090, P1_U4091, P1_U4092, P1_U4093, P1_U4094, P1_U4095, P1_U4096, P1_U4097, P1_U4098, P1_U4099, P1_U4100, P1_U4101, P1_U4102, P1_U4103, P1_U4104, P1_U4105, P1_U4106, P1_U4107, P1_U4108, P1_U4109, P1_U4110, P1_U4111, P1_U4112, P1_U4113, P1_U4114, P1_U4115, P1_U4116, P1_U4117, P1_U4118, P1_U4119, P1_U4120, P1_U4121, P1_U4122, P1_U4123, P1_U4124, P1_U4125, P1_U4126, P1_U4127, P1_U4128, P1_U4129, P1_U4130, P1_U4131, P1_U4132, P1_U4133, P1_U4134, P1_U4135, P1_U4136, P1_U4137, P1_U4138, P1_U4139, P1_U4140, P1_U4141, P1_U4142, P1_U4143, P1_U4144, P1_U4145, P1_U4146, P1_U4147, P1_U4148, P1_U4149, P1_U4150, P1_U4151, P1_U4152, P1_U4153, P1_U4154, P1_U4155, P1_U4156, P1_U4157, P1_U4158, P1_U4159, P1_U4160, P1_U4161, P1_U4162, P1_U4163, P1_U4164, P1_U4165, P1_U4166, P1_U4167, P1_U4168, P1_U4169, P1_U4170, P1_U4171, P1_U4172, P1_U4173, P1_U4174, P1_U4175, P1_U4176, P1_U4177, P1_U4178, P1_U4179, P1_U4180, P1_U4181, P1_U4182, P1_U4183, P1_U4184, P1_U4185, P1_U4186, P1_U4187, P1_U4188, P1_U4189, P1_U4190, P1_U4191, P1_U4192, P1_U4193, P1_U4194, P1_U4195, P1_U4196, P1_U4197, P1_U4198, P1_U4199, P1_U4200, P1_U4201, P1_U4202, P1_U4203, P1_U4204, P1_U4205, P1_U4206, P1_U4207, P1_U4208, P1_U4209, P1_U4210, P1_U4211, P1_U4212, P1_U4213, P1_U4214, P1_U4215, P1_U4216, P1_U4217, P1_U4218, P1_U4219, P1_U4220, P1_U4221, P1_U4222, P1_U4223, P1_U4224, P1_U4225, P1_U4226, P1_U4227, P1_U4228, P1_U4229, P1_U4230, P1_U4231, P1_U4232, P1_U4233, P1_U4234, P1_U4235, P1_U4236, P1_U4237, P1_U4238, P1_U4239, P1_U4240, P1_U4241, P1_U4242, P1_U4243, P1_U4244, P1_U4245, P1_U4246, P1_U4247, P1_U4248, P1_U4249, P1_U4250, P1_U4251, P1_U4252, P1_U4253, P1_U4254, P1_U4255, P1_U4256, P1_U4257, P1_U4258, P1_U4259, P1_U4260, P1_U4261, P1_U4262, P1_U4263, P1_U4264, P1_U4265, P1_U4266, P1_U4267, P1_U4268, P1_U4269, P1_U4270, P1_U4271, P1_U4272, P1_U4273, P1_U4274, P1_U4275, P1_U4276, P1_U4277, P1_U4278, P1_U4279, P1_U4280, P1_U4281, P1_U4282, P1_U4283, P1_U4284, P1_U4285, P1_U4286, P1_U4287, P1_U4288, P1_U4289, P1_U4290, P1_U4291, P1_U4292, P1_U4293, P1_U4294, P1_U4295, P1_U4296, P1_U4297, P1_U4298, P1_U4299, P1_U4300, P1_U4301, P1_U4302, P1_U4303, P1_U4304, P1_U4305, P1_U4306, P1_U4307, P1_U4308, P1_U4309, P1_U4310, P1_U4311, P1_U4312, P1_U4313, P1_U4314, P1_U4315, P1_U4316, P1_U4317, P1_U4318, P1_U4319, P1_U4320, P1_U4321, P1_U4322, P1_U4323, P1_U4324, P1_U4325, P1_U4326, P1_U4327, P1_U4328, P1_U4329, P1_U4330, P1_U4331, P1_U4332, P1_U4333, P1_U4334, P1_U4335, P1_U4336, P1_U4337, P1_U4338, P1_U4339, P1_U4340, P1_U4341, P1_U4342, P1_U4343, P1_U4344, P1_U4345, P1_U4346, P1_U4347, P1_U4348, P1_U4349, P1_U4350, P1_U4351, P1_U4352, P1_U4353, P1_U4354, P1_U4355, P1_U4356, P1_U4357, P1_U4358, P1_U4359, P1_U4360, P1_U4361, P1_U4362, P1_U4363, P1_U4364, P1_U4365, P1_U4366, P1_U4367, P1_U4368, P1_U4369, P1_U4370, P1_U4371, P1_U4372, P1_U4373, P1_U4374, P1_U4375, P1_U4376, P1_U4377, P1_U4378, P1_U4379, P1_U4380, P1_U4381, P1_U4382, P1_U4383, P1_U4384, P1_U4385, P1_U4386, P1_U4387, P1_U4388, P1_U4389, P1_U4390, P1_U4391, P1_U4392, P1_U4393, P1_U4394, P1_U4395, P1_U4396, P1_U4397, P1_U4398, P1_U4399, P1_U4400, P1_U4401, P1_U4402, P1_U4403, P1_U4404, P1_U4405, P1_U4406, P1_U4407, P1_U4408, P1_U4409, P1_U4410, P1_U4411, P1_U4412, P1_U4413, P1_U4414, P1_U4415, P1_U4416, P1_U4417, P1_U4418, P1_U4419, P1_U4420, P1_U4421, P1_U4422, P1_U4423, P1_U4424, P1_U4425, P1_U4426, P1_U4427, P1_U4428, P1_U4429, P1_U4430, P1_U4431, P1_U4432, P1_U4433, P1_U4434, P1_U4435, P1_U4436, P1_U4437, P1_U4438, P1_U4439, P1_U4440, P1_U4441, P1_U4442, P1_U4443, P1_U4444, P1_U4445, P1_U4446, P1_U4447, P1_U4448, P1_U4449, P1_U4450, P1_U4451, P1_U4452, P1_U4453, P1_U4454, P1_U4455, P1_U4456, P1_U4457, P1_U4458, P1_U4459, P1_U4460, P1_U4461, P1_U4462, P1_U4463, P1_U4464, P1_U4465, P1_U4466, P1_U4467, P1_U4468, P1_U4469, P1_U4470, P1_U4471, P1_U4472, P1_U4473, P1_U4474, P1_U4475, P1_U4476, P1_U4477, P1_U4478, P1_U4479, P1_U4480, P1_U4481, P1_U4482, P1_U4483, P1_U4484, P1_U4485, P1_U4486, P1_U4487, P1_U4488, P1_U4489, P1_U4490, P1_U4491, P1_U4492, P1_U4493, P1_U4494, P1_U4495, P1_U4496, P1_U4497, P1_U4498, P1_U4499, P1_U4500, P1_U4501, P1_U4502, P1_U4503, P1_U4504, P1_U4505, P1_U4506, P1_U4507, P1_U4508, P1_U4509, P1_U4510, P1_U4511, P1_U4512, P1_U4513, P1_U4514, P1_U4515, P1_U4516, P1_U4517, P1_U4518, P1_U4519, P1_U4520, P1_U4521, P1_U4522, P1_U4523, P1_U4524, P1_U4525, P1_U4526, P1_U4527, P1_U4528, P1_U4529, P1_U4530, P1_U4531, P1_U4532, P1_U4533, P1_U4534, P1_U4535, P1_U4536, P1_U4537, P1_U4538, P1_U4539, P1_U4540, P1_U4541, P1_U4542, P1_U4543, P1_U4544, P1_U4545, P1_U4546, P1_U4547, P1_U4548, P1_U4549, P1_U4550, P1_U4551, P1_U4552, P1_U4553, P1_U4554, P1_U4555, P1_U4556, P1_U4557, P1_U4558, P1_U4559, P1_U4560, P1_U4561, P1_U4562, P1_U4563, P1_U4564, P1_U4565, P1_U4566, P1_U4567, P1_U4568, P1_U4569, P1_U4570, P1_U4571, P1_U4572, P1_U4573, P1_U4574, P1_U4575, P1_U4576, P1_U4577, P1_U4578, P1_U4579, P1_U4580, P1_U4581, P1_U4582, P1_U4583, P1_U4584, P1_U4585, P1_U4586, P1_U4587, P1_U4588, P1_U4589, P1_U4590, P1_U4591, P1_U4592, P1_U4593, P1_U4594, P1_U4595, P1_U4596, P1_U4597, P1_U4598, P1_U4599, P1_U4600, P1_U4601, P1_U4602, P1_U4603, P1_U4604, P1_U4605, P1_U4606, P1_U4607, P1_U4608, P1_U4609, P1_U4610, P1_U4611, P1_U4612, P1_U4613, P1_U4614, P1_U4615, P1_U4616, P1_U4617, P1_U4618, P1_U4619, P1_U4620, P1_U4621, P1_U4622, P1_U4623, P1_U4624, P1_U4625, P1_U4626, P1_U4627, P1_U4628, P1_U4629, P1_U4630, P1_U4631, P1_U4632, P1_U4633, P1_U4634, P1_U4635, P1_U4636, P1_U4637, P1_U4638, P1_U4639, P1_U4640, P1_U4641, P1_U4642, P1_U4643, P1_U4644, P1_U4645, P1_U4646, P1_U4647, P1_U4648, P1_U4649, P1_U4650, P1_U4651, P1_U4652, P1_U4653, P1_U4654, P1_U4655, P1_U4656, P1_U4657, P1_U4658, P1_U4659, P1_U4660, P1_U4661, P1_U4662, P1_U4663, P1_U4664, P1_U4665, P1_U4666, P1_U4667, P1_U4668, P1_U4669, P1_U4670, P1_U4671, P1_U4672, P1_U4673, P1_U4674, P1_U4675, P1_U4676, P1_U4677, P1_U4678, P1_U4679, P1_U4680, P1_U4681, P1_U4682, P1_U4683, P1_U4684, P1_U4685, P1_U4686, P1_U4687, P1_U4688, P1_U4689, P1_U4690, P1_U4691, P1_U4692, P1_U4693, P1_U4694, P1_U4695, P1_U4696, P1_U4697, P1_U4698, P1_U4699, P1_U4700, P1_U4701, P1_U4702, P1_U4703, P1_U4704, P1_U4705, P1_U4706, P1_U4707, P1_U4708, P1_U4709, P1_U4710, P1_U4711, P1_U4712, P1_U4713, P1_U4714, P1_U4715, P1_U4716, P1_U4717, P1_U4718, P1_U4719, P1_U4720, P1_U4721, P1_U4722, P1_U4723, P1_U4724, P1_U4725, P1_U4726, P1_U4727, P1_U4728, P1_U4729, P1_U4730, P1_U4731, P1_U4732, P1_U4733, P1_U4734, P1_U4735, P1_U4736, P1_U4737, P1_U4738, P1_U4739, P1_U4740, P1_U4741, P1_U4742, P1_U4743, P1_U4744, P1_U4745, P1_U4746, P1_U4747, P1_U4748, P1_U4749, P1_U4750, P1_U4751, P1_U4752, P1_U4753, P1_U4754, P1_U4755, P1_U4756, P1_U4757, P1_U4758, P1_U4759, P1_U4760, P1_U4761, P1_U4762, P1_U4763, P1_U4764, P1_U4765, P1_U4766, P1_U4767, P1_U4768, P1_U4769, P1_U4770, P1_U4771, P1_U4772, P1_U4773, P1_U4774, P1_U4775, P1_U4776, P1_U4777, P1_U4778, P1_U4779, P1_U4780, P1_U4781, P1_U4782, P1_U4783, P1_U4784, P1_U4785, P1_U4786, P1_U4787, P1_U4788, P1_U4789, P1_U4790, P1_U4791, P1_U4792, P1_U4793, P1_U4794, P1_U4795, P1_U4796, P1_U4797, P1_U4798, P1_U4799, P1_U4800, P1_U4801, P1_U4802, P1_U4803, P1_U4804, P1_U4805, P1_U4806, P1_U4807, P1_U4808, P1_U4809, P1_U4810, P1_U4811, P1_U4812, P1_U4813, P1_U4814, P1_U4815, P1_U4816, P1_U4817, P1_U4818, P1_U4819, P1_U4820, P1_U4821, P1_U4822, P1_U4823, P1_U4824, P1_U4825, P1_U4826, P1_U4827, P1_U4828, P1_U4829, P1_U4830, P1_U4831, P1_U4832, P1_U4833, P1_U4834, P1_U4835, P1_U4836, P1_U4837, P1_U4838, P1_U4839, P1_U4840, P1_U4841, P1_U4842, P1_U4843, P1_U4844, P1_U4845, P1_U4846, P1_U4847, P1_U4848, P1_U4849, P1_U4850, P1_U4851, P1_U4852, P1_U4853, P1_U4854, P1_U4855, P1_U4856, P1_U4857, P1_U4858, P1_U4859, P1_U4860, P1_U4861, P1_U4862, P1_U4863, P1_U4864, P1_U4865, P1_U4866, P1_U4867, P1_U4868, P1_U4869, P1_U4870, P1_U4871, P1_U4872, P1_U4873, P1_U4874, P1_U4875, P1_U4876, P1_U4877, P1_U4878, P1_U4879, P1_U4880, P1_U4881, P1_U4882, P1_U4883, P1_U4884, P1_U4885, P1_U4886, P1_U4887, P1_U4888, P1_U4889, P1_U4890, P1_U4891, P1_U4892, P1_U4893, P1_U4894, P1_U4895, P1_U4896, P1_U4897, P1_U4898, P1_U4899, P1_U4900, P1_U4901, P1_U4902, P1_U4903, P1_U4904, P1_U4905, P1_U4906, P1_U4907, P1_U4908, P1_U4909, P1_U4910, P1_U4911, P1_U4912, P1_U4913, P1_U4914, P1_U4915, P1_U4916, P1_U4917, P1_U4918, P1_U4919, P1_U4920, P1_U4921, P1_U4922, P1_U4923, P1_U4924, P1_U4925, P1_U4926, P1_U4927, P1_U4928, P1_U4929, P1_U4930, P1_U4931, P1_U4932, P1_U4933, P1_U4934, P1_U4935, P1_U4936, P1_U4937, P1_U4938, P1_U4939, P1_U4940, P1_U4941, P1_U4942, P1_U4943, P1_U4944, P1_U4945, P1_U4946, P1_U4947, P1_U4948, P1_U4949, P1_U4950, P1_U4951, P1_U4952, P1_U4953, P1_U4954, P1_U4955, P1_U4956, P1_U4957, P1_U4958, P1_U4959, P1_U4960, P1_U4961, P1_U4962, P1_U4963, P1_U4964, P1_U4965, P1_U4966, P1_U4967, P1_U4968, P1_U4969, P1_U4970, P1_U4971, P1_U4972, P1_U4973, P1_U4974, P1_U4975, P1_U4976, P1_U4977, P1_U4978, P1_U4979, P1_U4980, P1_U4981, P1_U4982, P1_U4983, P1_U4984, P1_U4985, P1_U4986, P1_U4987, P1_U4988, P1_U4989, P1_U4990, P1_U4991, P1_U4992, P1_U4993, P1_U4994, P1_U4995, P1_U4996, P1_U4997, P1_U4998, P1_U4999, P1_U5000, P1_U5001, P1_U5002, P1_U5003, P1_U5004, P1_U5005, P1_U5006, P1_U5007, P1_U5008, P1_U5009, P1_U5010, P1_U5011, P1_U5012, P1_U5013, P1_U5014, P1_U5015, P1_U5016, P1_U5017, P1_U5018, P1_U5019, P1_U5020, P1_U5021, P1_U5022, P1_U5023, P1_U5024, P1_U5025, P1_U5026, P1_U5027, P1_U5028, P1_U5029, P1_U5030, P1_U5031, P1_U5032, P1_U5033, P1_U5034, P1_U5035, P1_U5036, P1_U5037, P1_U5038, P1_U5039, P1_U5040, P1_U5041, P1_U5042, P1_U5043, P1_U5044, P1_U5045, P1_U5046, P1_U5047, P1_U5048, P1_U5049, P1_U5050, P1_U5051, P1_U5052, P1_U5053, P1_U5054, P1_U5055, P1_U5056, P1_U5057, P1_U5058, P1_U5059, P1_U5060, P1_U5061, P1_U5062, P1_U5063, P1_U5064, P1_U5065, P1_U5066, P1_U5067, P1_U5068, P1_U5069, P1_U5070, P1_U5071, P1_U5072, P1_U5073, P1_U5074, P1_U5075, P1_U5076, P1_U5077, P1_U5078, P1_U5079, P1_U5080, P1_U5081, P1_U5082, P1_U5083, P1_U5084, P1_U5085, P1_U5086, P1_U5087, P1_U5088, P1_U5089, P1_U5090, P1_U5091, P1_U5092, P1_U5093, P1_U5094, P1_U5095, P1_U5096, P1_U5097, P1_U5098, P1_U5099, P1_U5100, P1_U5101, P1_U5102, P1_U5103, P1_U5104, P1_U5105, P1_U5106, P1_U5107, P1_U5108, P1_U5109, P1_U5110, P1_U5111, P1_U5112, P1_U5113, P1_U5114, P1_U5115, P1_U5116, P1_U5117, P1_U5118, P1_U5119, P1_U5120, P1_U5121, P1_U5122, P1_U5123, P1_U5124, P1_U5125, P1_U5126, P1_U5127, P1_U5128, P1_U5129, P1_U5130, P1_U5131, P1_U5132, P1_U5133, P1_U5134, P1_U5135, P1_U5136, P1_U5137, P1_U5138, P1_U5139, P1_U5140, P1_U5141, P1_U5142, P1_U5143, P1_U5144, P1_U5145, P1_U5146, P1_U5147, P1_U5148, P1_U5149, P1_U5150, P1_U5151, P1_U5152, P1_U5153, P1_U5154, P1_U5155, P1_U5156, P1_U5157, P1_U5158, P1_U5159, P1_U5160, P1_U5161, P1_U5162, P1_U5163, P1_U5164, P1_U5165, P1_U5166, P1_U5167, P1_U5168, P1_U5169, P1_U5170, P1_U5171, P1_U5172, P1_U5173, P1_U5174, P1_U5175, P1_U5176, P1_U5177, P1_U5178, P1_U5179, P1_U5180, P1_U5181, P1_U5182, P1_U5183, P1_U5184, P1_U5185, P1_U5186, P1_U5187, P1_U5188, P1_U5189, P1_U5190, P1_U5191, P1_U5192, P1_U5193, P1_U5194, P1_U5195, P1_U5196, P1_U5197, P1_U5198, P1_U5199, P1_U5200, P1_U5201, P1_U5202, P1_U5203, P1_U5204, P1_U5205, P1_U5206, P1_U5207, P1_U5208, P1_U5209, P1_U5210, P1_U5211, P1_U5212, P1_U5213, P1_U5214, P1_U5215, P1_U5216, P1_U5217, P1_U5218, P1_U5219, P1_U5220, P1_U5221, P1_U5222, P1_U5223, P1_U5224, P1_U5225, P1_U5226, P1_U5227, P1_U5228, P1_U5229, P1_U5230, P1_U5231, P1_U5232, P1_U5233, P1_U5234, P1_U5235, P1_U5236, P1_U5237, P1_U5238, P1_U5239, P1_U5240, P1_U5241, P1_U5242, P1_U5243, P1_U5244, P1_U5245, P1_U5246, P1_U5247, P1_U5248, P1_U5249, P1_U5250, P1_U5251, P1_U5252, P1_U5253, P1_U5254, P1_U5255, P1_U5256, P1_U5257, P1_U5258, P1_U5259, P1_U5260, P1_U5261, P1_U5262, P1_U5263, P1_U5264, P1_U5265, P1_U5266, P1_U5267, P1_U5268, P1_U5269, P1_U5270, P1_U5271, P1_U5272, P1_U5273, P1_U5274, P1_U5275, P1_U5276, P1_U5277, P1_U5278, P1_U5279, P1_U5280, P1_U5281, P1_U5282, P1_U5283, P1_U5284, P1_U5285, P1_U5286, P1_U5287, P1_U5288, P1_U5289, P1_U5290, P1_U5291, P1_U5292, P1_U5293, P1_U5294, P1_U5295, P1_U5296, P1_U5297, P1_U5298, P1_U5299, P1_U5300, P1_U5301, P1_U5302, P1_U5303, P1_U5304, P1_U5305, P1_U5306, P1_U5307, P1_U5308, P1_U5309, P1_U5310, P1_U5311, P1_U5312, P1_U5313, P1_U5314, P1_U5315, P1_U5316, P1_U5317, P1_U5318, P1_U5319, P1_U5320, P1_U5321, P1_U5322, P1_U5323, P1_U5324, P1_U5325, P1_U5326, P1_U5327, P1_U5328, P1_U5329, P1_U5330, P1_U5331, P1_U5332, P1_U5333, P1_U5334, P1_U5335, P1_U5336, P1_U5337, P1_U5338, P1_U5339, P1_U5340, P1_U5341, P1_U5342, P1_U5343, P1_U5344, P1_U5345, P1_U5346, P1_U5347, P1_U5348, P1_U5349, P1_U5350, P1_U5351, P1_U5352, P1_U5353, P1_U5354, P1_U5355, P1_U5356, P1_U5357, P1_U5358, P1_U5359, P1_U5360, P1_U5361, P1_U5362, P1_U5363, P1_U5364, P1_U5365, P1_U5366, P1_U5367, P1_U5368, P1_U5369, P1_U5370, P1_U5371, P1_U5372, P1_U5373, P1_U5374, P1_U5375, P1_U5376, P1_U5377, P1_U5378, P1_U5379, P1_U5380, P1_U5381, P1_U5382, P1_U5383, P1_U5384, P1_U5385, P1_U5386, P1_U5387, P1_U5388, P1_U5389, P1_U5390, P1_U5391, P1_U5392, P1_U5393, P1_U5394, P1_U5395, P1_U5396, P1_U5397, P1_U5398, P1_U5399, P1_U5400, P1_U5401, P1_U5402, P1_U5403, P1_U5404, P1_U5405, P1_U5406, P1_U5407, P1_U5408, P1_U5409, P1_U5410, P1_U5411, P1_U5412, P1_U5413, P1_U5414, P1_U5415, P1_U5416, P1_U5417, P1_U5418, P1_U5419, P1_U5420, P1_U5421, P1_U5422, P1_U5423, P1_U5424, P1_U5425, P1_U5426, P1_U5427, P1_U5428, P1_U5429, P1_U5430, P1_U5431, P1_U5432, P1_U5433, P1_U5434, P1_U5435, P1_U5436, P1_U5437, P1_U5438, P1_U5439, P1_U5440, P1_U5441, P1_U5442, P1_U5443, P1_U5444, P1_U5445, P1_U5446, P1_U5447, P1_U5448, P1_U5449, P1_U5450, P1_U5451, P1_U5452, P1_U5453, P1_U5454, P1_U5455, P1_U5456, P1_U5457, P1_U5458, P1_U5459, P1_U5460, P1_U5461, P1_U5462, P1_U5463, P1_U5464, P1_U5465, P1_U5466, P1_U5467, P1_U5468, P1_U5469, P1_U5470, P1_U5471, P1_U5472, P1_U5473, P1_U5474, P1_U5475, P1_U5476, P1_U5477, P1_U5478, P1_U5479, P1_U5480, P1_U5481, P1_U5482, P1_U5483, P1_U5484, P1_U5485, P1_U5486, P1_U5487, P1_U5488, P1_U5489, P1_U5490, P1_U5491, P1_U5492, P1_U5493, P1_U5494, P1_U5495, P1_U5496, P1_U5497, P1_U5498, P1_U5499, P1_U5500, P1_U5501, P1_U5502, P1_U5503, P1_U5504, P1_U5505, P1_U5506, P1_U5507, P1_U5508, P1_U5509, P1_U5510, P1_U5511, P1_U5512, P1_U5513, P1_U5514, P1_U5515, P1_U5516, P1_U5517, P1_U5518, P1_U5519, P1_U5520, P1_U5521, P1_U5522, P1_U5523, P1_U5524, P1_U5525, P1_U5526, P1_U5527, P1_U5528, P1_U5529, P1_U5530, P1_U5531, P1_U5532, P1_U5533, P1_U5534, P1_U5535, P1_U5536, P1_U5537, P1_U5538, P1_U5539, P1_U5540, P1_U5541, P1_U5542, P1_U5543, P1_U5544, P1_U5545, P1_U5546, P1_U5547, P1_U5548, P1_U5549, P1_U5550, P1_U5551, P1_U5552, P1_U5553, P1_U5554, P1_U5555, P1_U5556, P1_U5557, P1_U5558, P1_U5559, P1_U5560, P1_U5561, P1_U5562, P1_U5563, P1_U5564, P1_U5565, P1_U5566, P1_U5567, P1_U5568, P1_U5569, P1_U5570, P1_U5571, P1_U5572, P1_U5573, P1_U5574, P1_U5575, P1_U5576, P1_U5577, P1_U5578, P1_U5579, P1_U5580, P1_U5581, P1_U5582, P1_U5583, P1_U5584, P1_U5585, P1_U5586, P1_U5587, P1_U5588, P1_U5589, P1_U5590, P1_U5591, P1_U5592, P1_U5593, P1_U5594, P1_U5595, P1_U5596, P1_U5597, P1_U5598, P1_U5599, P1_U5600, P1_U5601, P1_U5602, P1_U5603, P1_U5604, P1_U5605, P1_U5606, P1_U5607, P1_U5608, P1_U5609, P1_U5610, P1_U5611, P1_U5612, P1_U5613, P1_U5614, P1_U5615, P1_U5616, P1_U5617, P1_U5618, P1_U5619, P1_U5620, P1_U5621, P1_U5622, P1_U5623, P1_U5624, P1_U5625, P1_U5626, P1_U5627, P1_U5628, P1_U5629, P1_U5630, P1_U5631, P1_U5632, P1_U5633, P1_U5634, P1_U5635, P1_U5636, P1_U5637, P1_U5638, P1_U5639, P1_U5640, P1_U5641, P1_U5642, P1_U5643, P1_U5644, P1_U5645, P1_U5646, P1_U5647, P1_U5648, P1_U5649, P1_U5650, P1_U5651, P1_U5652, P1_U5653, P1_U5654, P1_U5655, P1_U5656, P1_U5657, P1_U5658, P1_U5659, P1_U5660, P1_U5661, P1_U5662, P1_U5663, P1_U5664, P1_U5665, P1_U5666, P1_U5667, P1_U5668, P1_U5669, P1_U5670, P1_U5671, P1_U5672, P1_U5673, P1_U5674, P1_U5675, P1_U5676, P1_U5677, P1_U5678, P1_U5679, P1_U5680, P1_U5681, P1_U5682, P1_U5683, P1_U5684, P1_U5685, P1_U5686, P1_U5687, P1_U5688, P1_U5689, P1_U5690, P1_U5691, P1_U5692, P1_U5693, P1_U5694, P1_U5695, P1_U5696, P1_U5697, P1_U5698, P1_U5699, P1_U5700, P1_U5701, P1_U5702, P1_U5703, P1_U5704, P1_U5705, P1_U5706, P1_U5707, P1_U5708, P1_U5709, P1_U5710, P1_U5711, P1_U5712, P1_U5713, P1_U5714, P1_U5715, P1_U5716, P1_U5717, P1_U5718, P1_U5719, P1_U5720, P1_U5721, P1_U5722, P1_U5723, P1_U5724, P1_U5725, P1_U5726, P1_U5727, P1_U5728, P1_U5729, P1_U5730, P1_U5731, P1_U5732, P1_U5733, P1_U5734, P1_U5735, P1_U5736, P1_U5737, P1_U5738, P1_U5739, P1_U5740, P1_U5741, P1_U5742, P1_U5743, P1_U5744, P1_U5745, P1_U5746, P1_U5747, P1_U5748, P1_U5749, P1_U5750, P1_U5751, P1_U5752, P1_U5753, P1_U5754, P1_U5755, P1_U5756, P1_U5757, P1_U5758, P1_U5759, P1_U5760, P1_U5761, P1_U5762, P1_U5763, P1_U5764, P1_U5765, P1_U5766, P1_U5767, P1_U5768, P1_U5769, P1_U5770, P1_U5771, P1_U5772, P1_U5773, P1_U5774, P1_U5775, P1_U5776, P1_U5777, P1_U5778, P1_U5779, P1_U5780, P1_U5781, P1_U5782, P1_U5783, P1_U5784, P1_U5785, P1_U5786, P1_U5787, P1_U5788, P1_U5789, P1_U5790, P1_U5791, P1_U5792, P1_U5793, P1_U5794, P1_U5795, P1_U5796, P1_U5797, P1_U5798, P1_U5799, P1_U5800, P1_U5801, P1_U5802, P1_U5803, P1_U5804, P1_U5805, P1_U5806, P1_U5807, P1_U5808, P1_U5809, P1_U5810, P1_U5811, P1_U5812, P1_U5813, P1_U5814, P1_U5815, P1_U5816, P1_U5817, P1_U5818, P1_U5819, P1_U5820, P1_U5821, P1_U5822, P1_U5823, P1_U5824, P1_U5825, P1_U5826, P1_U5827, P1_U5828, P1_U5829, P1_U5830, P1_U5831, P1_U5832, P1_U5833, P1_U5834, P1_U5835, P1_U5836, P1_U5837, P1_U5838, P1_U5839, P1_U5840, P1_U5841, P1_U5842, P1_U5843, P1_U5844, P1_U5845, P1_U5846, P1_U5847, P1_U5848, P1_U5849, P1_U5850, P1_U5851, P1_U5852, P1_U5853, P1_U5854, P1_U5855, P1_U5856, P1_U5857, P1_U5858, P1_U5859, P1_U5860, P1_U5861, P1_U5862, P1_U5863, P1_U5864, P1_U5865, P1_U5866, P1_U5867, P1_U5868, P1_U5869, P1_U5870, P1_U5871, P1_U5872, P1_U5873, P1_U5874, P1_U5875, P1_U5876, P1_U5877, P1_U5878, P1_U5879, P1_U5880, P1_U5881, P1_U5882, P1_U5883, P1_U5884, P1_U5885, P1_U5886, P1_U5887, P1_U5888, P1_U5889, P1_U5890, P1_U5891, P1_U5892, P1_U5893, P1_U5894, P1_U5895, P1_U5896, P1_U5897, P1_U5898, P1_U5899, P1_U5900, P1_U5901, P1_U5902, P1_U5903, P1_U5904, P1_U5905, P1_U5906, P1_U5907, P1_U5908, P1_U5909, P1_U5910, P1_U5911, P1_U5912, P1_U5913, P1_U5914, P1_U5915, P1_U5916, P1_U5917, P1_U5918, P1_U5919, P1_U5920, P1_U5921, P1_U5922, P1_U5923, P1_U5924, P1_U5925, P1_U5926, P1_U5927, P1_U5928, P1_U5929, P1_U5930, P1_U5931, P1_U5932, P1_U5933, P1_U5934, P1_U5935, P1_U5936, P1_U5937, P1_U5938, P1_U5939, P1_U5940, P1_U5941, P1_U5942, P1_U5943, P1_U5944, P1_U5945, P1_U5946, P1_U5947, P1_U5948, P1_U5949, P1_U5950, P1_U5951, P1_U5952, P1_U5953, P1_U5954, P1_U5955, P1_U5956, P1_U5957, P1_U5958, P1_U5959, P1_U5960, P1_U5961, P1_U5962, P1_U5963, P1_U5964, P1_U5965, P1_U5966, P1_U5967, P1_U5968, P1_U5969, P1_U5970, P1_U5971, P1_U5972, P1_U5973, P1_U5974, P1_U5975, P1_U5976, P1_U5977, P1_U5978, P1_U5979, P1_U5980, P1_U5981, P1_U5982, P1_U5983, P1_U5984, P1_U5985, P1_U5986, P1_U5987, P1_U5988, P1_U5989, P1_U5990, P1_U5991, P1_U5992, P1_U5993, P1_U5994, P1_U5995, P1_U5996, P1_U5997, P1_U5998, P1_U5999, P1_U6000, P1_U6001, P1_U6002, P1_U6003, P1_U6004, P1_U6005, P1_U6006, P1_U6007, P1_U6008, P1_U6009, P1_U6010, P1_U6011, P1_U6012, P1_U6013, P1_U6014, P1_U6015, P1_U6016, P1_U6017, P1_U6018, P1_U6019, P1_U6020, P1_U6021, P1_U6022, P1_U6023, P1_U6024, P1_U6025, P1_U6026, P1_U6027, P1_U6028, P1_U6029, P1_U6030, P1_U6031, P1_U6032, P1_U6033, P1_U6034, P1_U6035, P1_U6036, P1_U6037, P1_U6038, P1_U6039, P1_U6040, P1_U6041, P1_U6042, P1_U6043, P1_U6044, P1_U6045, P1_U6046, P1_U6047, P1_U6048, P1_U6049, P1_U6050, P1_U6051, P1_U6052, P1_U6053, P1_U6054, P1_U6055, P1_U6056, P1_U6057, P1_U6058, P1_U6059, P1_U6060, P1_U6061, P1_U6062, P1_U6063, P1_U6064, P1_U6065, P1_U6066, P1_U6067, P1_U6068, P1_U6069, P1_U6070, P1_U6071, P1_U6072, P1_U6073, P1_U6074, P1_U6075, P1_U6076, P1_U6077, P1_U6078, P1_U6079, P1_U6080, P1_U6081, P1_U6082, P1_U6083, P1_U6084, P1_U6085, P1_U6086, P1_U6087, P1_U6088, P1_U6089, P1_U6090, P1_U6091, P1_U6092, P1_U6093, P1_U6094, P1_U6095, P1_U6096, P1_U6097, P1_U6098, P1_U6099, P1_U6100, P1_U6101, P1_U6102, P1_U6103, P1_U6104, P1_U6105, P1_U6106, P1_U6107, P1_U6108, P1_U6109, P1_U6110, P1_U6111, P1_U6112, P1_U6113, P1_U6114, P1_U6115, P1_U6116, P1_U6117, P1_U6118, P1_U6119, P1_U6120, P1_U6121, P1_U6122, P1_U6123, P1_U6124, P1_U6125, P1_U6126, P1_U6127, P1_U6128, P1_U6129, P1_U6130, P1_U6131, P1_U6132, P1_U6133, P1_U6134, P1_U6135, P1_U6136, P1_U6137, P1_U6138, P1_U6139, P1_U6140, P1_U6141, P1_U6142, P1_U6143, P1_U6144, P1_U6145, P1_U6146, P1_U6147, P1_U6148, P1_U6149, P1_U6150, P1_U6151, P1_U6152, P1_U6153, P1_U6154, P1_U6155, P1_U6156, P1_U6157, P1_U6158, P1_U6159, P1_U6160, P1_U6161, P1_U6162, P1_U6163, P1_U6164, P1_U6165, P1_U6166, P1_U6167, P1_U6168, P1_U6169, P1_U6170, P1_U6171, P1_U6172, P1_U6173, P1_U6174, P1_U6175, P1_U6176, P1_U6177, P1_U6178, P1_U6179, P1_U6180, P1_U6181, P1_U6182, P1_U6183, P1_U6184, P1_U6185, P1_U6186, P1_U6187, P1_U6188, P1_U6189, P1_U6190, P1_U6191, P1_U6192, P1_U6193, P1_U6194, P1_U6195, P1_U6196, P1_U6197, P1_U6198, P1_U6199, P1_U6200, P1_U6201, P1_U6202, P1_U6203, P1_U6204, P1_U6205, P1_U6206, P1_U6207, P1_U6208, P1_U6209, P1_U6210, P1_U6211, P1_U6212, P1_U6213, P1_U6214, P1_U6215, P1_U6216, P1_U6217, P1_U6218, P1_U6219, P1_U6220, P1_U6221, P1_U6222, P1_U6223, P1_U6224, P1_U6225, P1_U6226, P1_U6227, P1_U6228, P1_U6229, P1_U6230, P1_U6231, P1_U6232, P1_U6233, P1_U6234, P1_U6235, P1_U6236, P1_U6237, P1_U6238, P1_U6239, P1_U6240, P1_U6241, P1_U6242, P1_U6243, P1_U6244, P1_U6245, P1_U6246, P1_U6247, P1_U6248, P1_U6249, P1_U6250, P1_U6251, P1_U6252, P1_U6253, P1_U6254, P1_U6255, P1_U6256, P1_U6257, P1_U6258, P1_U6259, P1_U6260, P1_U6261, P1_U6262, P1_U6263, P1_U6264, P1_U6265, P1_U6266, P1_U6267, P1_U6268, P1_U6269, P1_U6270, P1_U6271, P1_U6272, P1_U6273, P1_U6274, P1_U6275, P1_U6276, P1_U6277, P1_U6278, P1_U6279, P1_U6280, P1_U6281, P1_U6282, P1_U6283, P1_U6284, P1_U6285, P1_U6286, P1_U6287, P1_U6288, P1_U6289, P1_U6290, P1_U6291, P1_U6292, P1_U6293, P1_U6294, P1_U6295, P1_U6296, P1_U6297, P1_U6298, P1_U6299, P1_U6300, P1_U6301, P1_U6302, P1_U6303, P1_U6304, P1_U6305, P1_U6306, P1_U6307, P1_U6308, P1_U6309, P1_U6310, P1_U6311, P1_U6312, P1_U6313, P1_U6314, P1_U6315, P1_U6316, P1_U6317, P1_U6318, P1_U6319, P1_U6320, P1_U6321, P1_U6322, P1_U6323, P1_U6324, P1_U6325, P1_U6326, P1_U6327, P1_U6328, P1_U6329, P1_U6330, P1_U6331, P1_U6332, P1_U6333, P1_U6334, P1_U6335, P1_U6336, P1_U6337, P1_U6338, P1_U6339, P1_U6340, P1_U6341, P1_U6342, P1_U6343, P1_U6344, P1_U6345, P1_U6346, P1_U6347, P1_U6348, P1_U6349, P1_U6350, P1_U6351, P1_U6352, P1_U6353, P1_U6354, P1_U6355, P1_U6356, P1_U6357, P1_U6358, P1_U6359, P1_U6360, P1_U6361, P1_U6362, P1_U6363, P1_U6364, P1_U6365, P1_U6366, P1_U6367, P1_U6368, P1_U6369, P1_U6370, P1_U6371, P1_U6372, P1_U6373, P1_U6374, P1_U6375, P1_U6376, P1_U6377, P1_U6378, P1_U6379, P1_U6380, P1_U6381, P1_U6382, P1_U6383, P1_U6384, P1_U6385, P1_U6386, P1_U6387, P1_U6388, P1_U6389, P1_U6390, P1_U6391, P1_U6392, P1_U6393, P1_U6394, P1_U6395, P1_U6396, P1_U6397, P1_U6398, P1_U6399, P1_U6400, P1_U6401, P1_U6402, P1_U6403, P1_U6404, P1_U6405, P1_U6406, P1_U6407, P1_U6408, P1_U6409, P1_U6410, P1_U6411, P1_U6412, P1_U6413, P1_U6414, P1_U6415, P1_U6416, P1_U6417, P1_U6418, P1_U6419, P1_U6420, P1_U6421, P1_U6422, P1_U6423, P1_U6424, P1_U6425, P1_U6426, P1_U6427, P1_U6428, P1_U6429, P1_U6430, P1_U6431, P1_U6432, P1_U6433, P1_U6434, P1_U6435, P1_U6436, P1_U6437, P1_U6438, P1_U6439, P1_U6440, P1_U6441, P1_U6442, P1_U6443, P1_U6444, P1_U6445, P1_U6446, P1_U6447, P1_U6448, P1_U6449, P1_U6450, P1_U6451, P1_U6452, P1_U6453, P1_U6454, P1_U6455, P1_U6456, P1_U6457, P1_U6458, P1_U6459, P1_U6460, P1_U6461, P1_U6462, P1_U6463, P1_U6464, P1_U6465, P1_U6466, P1_U6467, P1_U6468, P1_U6469, P1_U6470, P1_U6471, P1_U6472, P1_U6473, P1_U6474, P1_U6475, P1_U6476, P1_U6477, P1_U6478, P1_U6479, P1_U6480, P1_U6481, P1_U6482, P1_U6483, P1_U6484, P1_U6485, P1_U6486, P1_U6487, P1_U6488, P1_U6489, P1_U6490, P1_U6491, P1_U6492, P1_U6493, P1_U6494, P1_U6495, P1_U6496, P1_U6497, P1_U6498, P1_U6499, P1_U6500, P1_U6501, P1_U6502, P1_U6503, P1_U6504, P1_U6505, P1_U6506, P1_U6507, P1_U6508, P1_U6509, P1_U6510, P1_U6511, P1_U6512, P1_U6513, P1_U6514, P1_U6515, P1_U6516, P1_U6517, P1_U6518, P1_U6519, P1_U6520, P1_U6521, P1_U6522, P1_U6523, P1_U6524, P1_U6525, P1_U6526, P1_U6527, P1_U6528, P1_U6529, P1_U6530, P1_U6531, P1_U6532, P1_U6533, P1_U6534, P1_U6535, P1_U6536, P1_U6537, P1_U6538, P1_U6539, P1_U6540, P1_U6541, P1_U6542, P1_U6543, P1_U6544, P1_U6545, P1_U6546, P1_U6547, P1_U6548, P1_U6549, P1_U6550, P1_U6551, P1_U6552, P1_U6553, P1_U6554, P1_U6555, P1_U6556, P1_U6557, P1_U6558, P1_U6559, P1_U6560, P1_U6561, P1_U6562, P1_U6563, P1_U6564, P1_U6565, P1_U6566, P1_U6567, P1_U6568, P1_U6569, P1_U6570, P1_U6571, P1_U6572, P1_U6573, P1_U6574, P1_U6575, P1_U6576, P1_U6577, P1_U6578, P1_U6579, P1_U6580, P1_U6581, P1_U6582, P1_U6583, P1_U6584, P1_U6585, P1_U6586, P1_U6587, P1_U6588, P1_U6589, P1_U6590, P1_U6591, P1_U6592, P1_U6593, P1_U6594, P1_U6595, P1_U6596, P1_U6597, P1_U6598, P1_U6599, P1_U6600, P1_U6601, P1_U6602, P1_U6603, P1_U6604, P1_U6605, P1_U6606, P1_U6607, P1_U6608, P1_U6609, P1_U6610, P1_U6611, P1_U6612, P1_U6613, P1_U6614, P1_U6615, P1_U6616, P1_U6617, P1_U6618, P1_U6619, P1_U6620, P1_U6621, P1_U6622, P1_U6623, P1_U6624, P1_U6625, P1_U6626, P1_U6627, P1_U6628, P1_U6629, P1_U6630, P1_U6631, P1_U6632, P1_U6633, P1_U6634, P1_U6635, P1_U6636, P1_U6637, P1_U6638, P1_U6639, P1_U6640, P1_U6641, P1_U6642, P1_U6643, P1_U6644, P1_U6645, P1_U6646, P1_U6647, P1_U6648, P1_U6649, P1_U6650, P1_U6651, P1_U6652, P1_U6653, P1_U6654, P1_U6655, P1_U6656, P1_U6657, P1_U6658, P1_U6659, P1_U6660, P1_U6661, P1_U6662, P1_U6663, P1_U6664, P1_U6665, P1_U6666, P1_U6667, P1_U6668, P1_U6669, P1_U6670, P1_U6671, P1_U6672, P1_U6673, P1_U6674, P1_U6675, P1_U6676, P1_U6677, P1_U6678, P1_U6679, P1_U6680, P1_U6681, P1_U6682, P1_U6683, P1_U6684, P1_U6685, P1_U6686, P1_U6687, P1_U6688, P1_U6689, P1_U6690, P1_U6691, P1_U6692, P1_U6693, P1_U6694, P1_U6695, P1_U6696, P1_U6697, P1_U6698, P1_U6699, P1_U6700, P1_U6701, P1_U6702, P1_U6703, P1_U6704, P1_U6705, P1_U6706, P1_U6707, P1_U6708, P1_U6709, P1_U6710, P1_U6711, P1_U6712, P1_U6713, P1_U6714, P1_U6715, P1_U6716, P1_U6717, P1_U6718, P1_U6719, P1_U6720, P1_U6721, P1_U6722, P1_U6723, P1_U6724, P1_U6725, P1_U6726, P1_U6727, P1_U6728, P1_U6729, P1_U6730, P1_U6731, P1_U6732, P1_U6733, P1_U6734, P1_U6735, P1_U6736, P1_U6737, P1_U6738, P1_U6739, P1_U6740, P1_U6741, P1_U6742, P1_U6743, P1_U6744, P1_U6745, P1_U6746, P1_U6747, P1_U6748, P1_U6749, P1_U6750, P1_U6751, P1_U6752, P1_U6753, P1_U6754, P1_U6755, P1_U6756, P1_U6757, P1_U6758, P1_U6759, P1_U6760, P1_U6761, P1_U6762, P1_U6763, P1_U6764, P1_U6765, P1_U6766, P1_U6767, P1_U6768, P1_U6769, P1_U6770, P1_U6771, P1_U6772, P1_U6773, P1_U6774, P1_U6775, P1_U6776, P1_U6777, P1_U6778, P1_U6779, P1_U6780, P1_U6781, P1_U6782, P1_U6783, P1_U6784, P1_U6785, P1_U6786, P1_U6787, P1_U6788, P1_U6789, P1_U6790, P1_U6791, P1_U6792, P1_U6793, P1_U6794, P1_U6795, P1_U6796, P1_U6797, P1_U6798, P1_U6799, P1_U6800, P1_U6801, P1_U6802, P1_U6803, P1_U6804, P1_U6805, P1_U6806, P1_U6807, P1_U6808, P1_U6809, P1_U6810, P1_U6811, P1_U6812, P1_U6813, P1_U6814, P1_U6815, P1_U6816, P1_U6817, P1_U6818, P1_U6819, P1_U6820, P1_U6821, P1_U6822, P1_U6823, P1_U6824, P1_U6825, P1_U6826, P1_U6827, P1_U6828, P1_U6829, P1_U6830, P1_U6831, P1_U6832, P1_U6833, P1_U6834, P1_U6835, P1_U6836, P1_U6837, P1_U6838, P1_U6839, P1_U6840, P1_U6841, P1_U6842, P1_U6843, P1_U6844, P1_U6845, P1_U6846, P1_U6847, P1_U6848, P1_U6849, P1_U6850, P1_U6851, P1_U6852, P1_U6853, P1_U6854, P1_U6855, P1_U6856, P1_U6857, P1_U6858, P1_U6859, P1_U6860, P1_U6861, P1_U6862, P1_U6863, P1_U6864, P1_U6865, P1_U6866, P1_U6867, P1_U6868, P1_U6869, P1_U6870, P1_U6871, P1_U6872, P1_U6873, P1_U6874, P1_U6875, P1_U6876, P1_U6877, P1_U6878, P1_U6879, P1_U6880, P1_U6881, P1_U6882, P1_U6883, P1_U6884, P1_U6885, P1_U6886, P1_U6887, P1_U6888, P1_U6889, P1_U6890, P1_U6891, P1_U6892, P1_U6893, P1_U6894, P1_U6895, P1_U6896, P1_U6897, P1_U6898, P1_U6899, P1_U6900, P1_U6901, P1_U6902, P1_U6903, P1_U6904, P1_U6905, P1_U6906, P1_U6907, P1_U6908, P1_U6909, P1_U6910, P1_U6911, P1_U6912, P1_U6913, P1_U6914, P1_U6915, P1_U6916, P1_U6917, P1_U6918, P1_U6919, P1_U6920, P1_U6921, P1_U6922, P1_U6923, P1_U6924, P1_U6925, P1_U6926, P1_U6927, P1_U6928, P1_U6929, P1_U6930, P1_U6931, P1_U6932, P1_U6933, P1_U6934, P1_U6935, P1_U6936, P1_U6937, P1_U6938, P1_U6939, P1_U6940, P1_U6941, P1_U6942, P1_U6943, P1_U6944, P1_U6945, P1_U6946, P1_U6947, P1_U6948, P1_U6949, P1_U6950, P1_U6951, P1_U6952, P1_U6953, P1_U6954, P1_U6955, P1_U6956, P1_U6957, P1_U6958, P1_U6959, P1_U6960, P1_U6961, P1_U6962, P1_U6963, P1_U6964, P1_U6965, P1_U6966, P1_U6967, P1_U6968, P1_U6969, P1_U6970, P1_U6971, P1_U6972, P1_U6973, P1_U6974, P1_U6975, P1_U6976, P1_U6977, P1_U6978, P1_U6979, P1_U6980, P1_U6981, P1_U6982, P1_U6983, P1_U6984, P1_U6985, P1_U6986, P1_U6987, P1_U6988, P1_U6989, P1_U6990, P1_U6991, P1_U6992, P1_U6993, P1_U6994, P1_U6995, P1_U6996, P1_U6997, P1_U6998, P1_U6999, P1_U7000, P1_U7001, P1_U7002, P1_U7003, P1_U7004, P1_U7005, P1_U7006, P1_U7007, P1_U7008, P1_U7009, P1_U7010, P1_U7011, P1_U7012, P1_U7013, P1_U7014, P1_U7015, P1_U7016, P1_U7017, P1_U7018, P1_U7019, P1_U7020, P1_U7021, P1_U7022, P1_U7023, P1_U7024, P1_U7025, P1_U7026, P1_U7027, P1_U7028, P1_U7029, P1_U7030, P1_U7031, P1_U7032, P1_U7033, P1_U7034, P1_U7035, P1_U7036, P1_U7037, P1_U7038, P1_U7039, P1_U7040, P1_U7041, P1_U7042, P1_U7043, P1_U7044, P1_U7045, P1_U7046, P1_U7047, P1_U7048, P1_U7049, P1_U7050, P1_U7051, P1_U7052, P1_U7053, P1_U7054, P1_U7055, P1_U7056, P1_U7057, P1_U7058, P1_U7059, P1_U7060, P1_U7061, P1_U7062, P1_U7063, P1_U7064, P1_U7065, P1_U7066, P1_U7067, P1_U7068, P1_U7069, P1_U7070, P1_U7071, P1_U7072, P1_U7073, P1_U7074, P1_U7075, P1_U7076, P1_U7077, P1_U7078, P1_U7079, P1_U7080, P1_U7081, P1_U7082, P1_U7083, P1_U7084, P1_U7085, P1_U7086, P1_U7087, P1_U7088, P1_U7089, P1_U7090, P1_U7091, P1_U7092, P1_U7093, P1_U7094, P1_U7095, P1_U7096, P1_U7097, P1_U7098, P1_U7099, P1_U7100, P1_U7101, P1_U7102, P1_U7103, P1_U7104, P1_U7105, P1_U7106, P1_U7107, P1_U7108, P1_U7109, P1_U7110, P1_U7111, P1_U7112, P1_U7113, P1_U7114, P1_U7115, P1_U7116, P1_U7117, P1_U7118, P1_U7119, P1_U7120, P1_U7121, P1_U7122, P1_U7123, P1_U7124, P1_U7125, P1_U7126, P1_U7127, P1_U7128, P1_U7129, P1_U7130, P1_U7131, P1_U7132, P1_U7133, P1_U7134, P1_U7135, P1_U7136, P1_U7137, P1_U7138, P1_U7139, P1_U7140, P1_U7141, P1_U7142, P1_U7143, P1_U7144, P1_U7145, P1_U7146, P1_U7147, P1_U7148, P1_U7149, P1_U7150, P1_U7151, P1_U7152, P1_U7153, P1_U7154, P1_U7155, P1_U7156, P1_U7157, P1_U7158, P1_U7159, P1_U7160, P1_U7161, P1_U7162, P1_U7163, P1_U7164, P1_U7165, P1_U7166, P1_U7167, P1_U7168, P1_U7169, P1_U7170, P1_U7171, P1_U7172, P1_U7173, P1_U7174, P1_U7175, P1_U7176, P1_U7177, P1_U7178, P1_U7179, P1_U7180, P1_U7181, P1_U7182, P1_U7183, P1_U7184, P1_U7185, P1_U7186, P1_U7187, P1_U7188, P1_U7189, P1_U7190, P1_U7191, P1_U7192, P1_U7193, P1_U7194, P1_U7195, P1_U7196, P1_U7197, P1_U7198, P1_U7199, P1_U7200, P1_U7201, P1_U7202, P1_U7203, P1_U7204, P1_U7205, P1_U7206, P1_U7207, P1_U7208, P1_U7209, P1_U7210, P1_U7211, P1_U7212, P1_U7213, P1_U7214, P1_U7215, P1_U7216, P1_U7217, P1_U7218, P1_U7219, P1_U7220, P1_U7221, P1_U7222, P1_U7223, P1_U7224, P1_U7225, P1_U7226, P1_U7227, P1_U7228, P1_U7229, P1_U7230, P1_U7231, P1_U7232, P1_U7233, P1_U7234, P1_U7235, P1_U7236, P1_U7237, P1_U7238, P1_U7239, P1_U7240, P1_U7241, P1_U7242, P1_U7243, P1_U7244, P1_U7245, P1_U7246, P1_U7247, P1_U7248, P1_U7249, P1_U7250, P1_U7251, P1_U7252, P1_U7253, P1_U7254, P1_U7255, P1_U7256, P1_U7257, P1_U7258, P1_U7259, P1_U7260, P1_U7261, P1_U7262, P1_U7263, P1_U7264, P1_U7265, P1_U7266, P1_U7267, P1_U7268, P1_U7269, P1_U7270, P1_U7271, P1_U7272, P1_U7273, P1_U7274, P1_U7275, P1_U7276, P1_U7277, P1_U7278, P1_U7279, P1_U7280, P1_U7281, P1_U7282, P1_U7283, P1_U7284, P1_U7285, P1_U7286, P1_U7287, P1_U7288, P1_U7289, P1_U7290, P1_U7291, P1_U7292, P1_U7293, P1_U7294, P1_U7295, P1_U7296, P1_U7297, P1_U7298, P1_U7299, P1_U7300, P1_U7301, P1_U7302, P1_U7303, P1_U7304, P1_U7305, P1_U7306, P1_U7307, P1_U7308, P1_U7309, P1_U7310, P1_U7311, P1_U7312, P1_U7313, P1_U7314, P1_U7315, P1_U7316, P1_U7317, P1_U7318, P1_U7319, P1_U7320, P1_U7321, P1_U7322, P1_U7323, P1_U7324, P1_U7325, P1_U7326, P1_U7327, P1_U7328, P1_U7329, P1_U7330, P1_U7331, P1_U7332, P1_U7333, P1_U7334, P1_U7335, P1_U7336, P1_U7337, P1_U7338, P1_U7339, P1_U7340, P1_U7341, P1_U7342, P1_U7343, P1_U7344, P1_U7345, P1_U7346, P1_U7347, P1_U7348, P1_U7349, P1_U7350, P1_U7351, P1_U7352, P1_U7353, P1_U7354, P1_U7355, P1_U7356, P1_U7357, P1_U7358, P1_U7359, P1_U7360, P1_U7361, P1_U7362, P1_U7363, P1_U7364, P1_U7365, P1_U7366, P1_U7367, P1_U7368, P1_U7369, P1_U7370, P1_U7371, P1_U7372, P1_U7373, P1_U7374, P1_U7375, P1_U7376, P1_U7377, P1_U7378, P1_U7379, P1_U7380, P1_U7381, P1_U7382, P1_U7383, P1_U7384, P1_U7385, P1_U7386, P1_U7387, P1_U7388, P1_U7389, P1_U7390, P1_U7391, P1_U7392, P1_U7393, P1_U7394, P1_U7395, P1_U7396, P1_U7397, P1_U7398, P1_U7399, P1_U7400, P1_U7401, P1_U7402, P1_U7403, P1_U7404, P1_U7405, P1_U7406, P1_U7407, P1_U7408, P1_U7409, P1_U7410, P1_U7411, P1_U7412, P1_U7413, P1_U7414, P1_U7415, P1_U7416, P1_U7417, P1_U7418, P1_U7419, P1_U7420, P1_U7421, P1_U7422, P1_U7423, P1_U7424, P1_U7425, P1_U7426, P1_U7427, P1_U7428, P1_U7429, P1_U7430, P1_U7431, P1_U7432, P1_U7433, P1_U7434, P1_U7435, P1_U7436, P1_U7437, P1_U7438, P1_U7439, P1_U7440, P1_U7441, P1_U7442, P1_U7443, P1_U7444, P1_U7445, P1_U7446, P1_U7447, P1_U7448, P1_U7449, P1_U7450, P1_U7451, P1_U7452, P1_U7453, P1_U7454, P1_U7455, P1_U7456, P1_U7457, P1_U7458, P1_U7459, P1_U7460, P1_U7461, P1_U7462, P1_U7463, P1_U7464, P1_U7465, P1_U7466, P1_U7467, P1_U7468, P1_U7469, P1_U7470, P1_U7471, P1_U7472, P1_U7473, P1_U7474, P1_U7475, P1_U7476, P1_U7477, P1_U7478, P1_U7479, P1_U7480, P1_U7481, P1_U7482, P1_U7483, P1_U7484, P1_U7485, P1_U7486, P1_U7487, P1_U7488, P1_U7489, P1_U7490, P1_U7491, P1_U7492, P1_U7493, P1_U7494, P1_U7495, P1_U7496, P1_U7497, P1_U7498, P1_U7499, P1_U7500, P1_U7501, P1_U7502, P1_U7503, P1_U7504, P1_U7505, P1_U7506, P1_U7507, P1_U7508, P1_U7509, P1_U7510, P1_U7511, P1_U7512, P1_U7513, P1_U7514, P1_U7515, P1_U7516, P1_U7517, P1_U7518, P1_U7519, P1_U7520, P1_U7521, P1_U7522, P1_U7523, P1_U7524, P1_U7525, P1_U7526, P1_U7527, P1_U7528, P1_U7529, P1_U7530, P1_U7531, P1_U7532, P1_U7533, P1_U7534, P1_U7535, P1_U7536, P1_U7537, P1_U7538, P1_U7539, P1_U7540, P1_U7541, P1_U7542, P1_U7543, P1_U7544, P1_U7545, P1_U7546, P1_U7547, P1_U7548, P1_U7549, P1_U7550, P1_U7551, P1_U7552, P1_U7553, P1_U7554, P1_U7555, P1_U7556, P1_U7557, P1_U7558, P1_U7559, P1_U7560, P1_U7561, P1_U7562, P1_U7563, P1_U7564, P1_U7565, P1_U7566, P1_U7567, P1_U7568, P1_U7569, P1_U7570, P1_U7571, P1_U7572, P1_U7573, P1_U7574, P1_U7575, P1_U7576, P1_U7577, P1_U7578, P1_U7579, P1_U7580, P1_U7581, P1_U7582, P1_U7583, P1_U7584, P1_U7585, P1_U7586, P1_U7587, P1_U7588, P1_U7589, P1_U7590, P1_U7591, P1_U7592, P1_U7593, P1_U7594, P1_U7595, P1_U7596, P1_U7597, P1_U7598, P1_U7599, P1_U7600, P1_U7601, P1_U7602, P1_U7603, P1_U7604, P1_U7605, P1_U7606, P1_U7607, P1_U7608, P1_U7609, P1_U7610, P1_U7611, P1_U7612, P1_U7613, P1_U7614, P1_U7615, P1_U7616, P1_U7617, P1_U7618, P1_U7619, P1_U7620, P1_U7621, P1_U7622, P1_U7623, P1_U7624, P1_U7625, P1_U7626, P1_U7627, P1_U7628, P1_U7629, P1_U7630, P1_U7631, P1_U7632, P1_U7633, P1_U7634, P1_U7635, P1_U7636, P1_U7637, P1_U7638, P1_U7639, P1_U7640, P1_U7641, P1_U7642, P1_U7643, P1_U7644, P1_U7645, P1_U7646, P1_U7647, P1_U7648, P1_U7649, P1_U7650, P1_U7651, P1_U7652, P1_U7653, P1_U7654, P1_U7655, P1_U7656, P1_U7657, P1_U7658, P1_U7659, P1_U7660, P1_U7661, P1_U7662, P1_U7663, P1_U7664, P1_U7665, P1_U7666, P1_U7667, P1_U7668, P1_U7669, P1_U7670, P1_U7671, P1_U7672, P1_U7673, P1_U7674, P1_U7675, P1_U7676, P1_U7677, P1_U7678, P1_U7679, P1_U7680, P1_U7681, P1_U7682, P1_U7683, P1_U7684, P1_U7685, P1_U7686, P1_U7687, P1_U7688, P1_U7689, P1_U7690, P1_U7691, P1_U7692, P1_U7693, P1_U7694, P1_U7695, P1_U7696, P1_U7697, P1_U7698, P1_U7699, P1_U7700, P1_U7701, P1_U7702, P1_U7703, P1_U7704, P1_U7705, P1_U7706, P1_U7707, P1_U7708, P1_U7709, P1_U7710, P1_U7711, P1_U7712, P1_U7713, P1_U7714, P1_U7715, P1_U7716, P1_U7717, P1_U7718, P1_U7719, P1_U7720, P1_U7721, P1_U7722, P1_U7723, P1_U7724, P1_U7725, P1_U7726, P1_U7727, P1_U7728, P1_U7729, P1_U7730, P1_U7731, P1_U7732, P1_U7733, P1_U7734, P1_U7735, P1_U7736, P1_U7737, P1_U7738, P1_U7739, P1_U7740, P1_U7741, P1_U7742, P1_U7743, P1_U7744, P1_U7745, P1_U7746, P1_U7747, P1_U7748, P1_U7749, P1_U7750, P1_U7751, P1_U7752, P1_U7753, P1_U7754, P1_U7755, P1_U7756, P1_U7757, P1_U7758, P1_U7759, P1_U7760, P1_U7761, P1_U7762, P1_U7763, P1_U7764, P1_U7765, P1_U7766, P1_U7767, P1_U7768, P1_U7769, P1_U7770, P1_U7771, P1_U7772, P1_U7773, P1_U7774, P1_U7775, P1_U7776, P1_U7777, P1_U7778, P1_U7779, P1_U7780, P1_U7781, P1_U7782, P1_U7783, P1_U7784, P1_U7785, P1_U7786, P1_U7787, P1_U7788, P1_U7789, P1_U7790, P1_U7791, P1_U7792, P1_U7793, P1_U7794, LT_782_120_U6, LT_782_120_U7, LT_782_U6, LT_782_U7, LT_748_U6, R170_U6, R170_U7, R170_U8, R170_U9, R170_U10, R170_U11, R170_U12, R170_U13, R170_U14, R170_U15, R165_U6, R165_U7, R165_U8, R165_U9, R165_U10, R165_U11, R165_U12, R165_U13, R165_U14, R165_U15, LT_782_119_U6, LT_782_119_U7, P3_ADD_526_U5, P3_ADD_526_U6, P3_ADD_526_U7, P3_ADD_526_U8, P3_ADD_526_U9, P3_ADD_526_U10, P3_ADD_526_U11, P3_ADD_526_U12, P3_ADD_526_U13, P3_ADD_526_U14, P3_ADD_526_U15, P3_ADD_526_U16, P3_ADD_526_U17, P3_ADD_526_U18, P3_ADD_526_U19, P3_ADD_526_U20, P3_ADD_526_U21, P3_ADD_526_U22, P3_ADD_526_U23, P3_ADD_526_U24, P3_ADD_526_U25, P3_ADD_526_U26, P3_ADD_526_U27, P3_ADD_526_U28, P3_ADD_526_U29, P3_ADD_526_U30, P3_ADD_526_U31, P3_ADD_526_U32, P3_ADD_526_U33, P3_ADD_526_U34, P3_ADD_526_U35, P3_ADD_526_U36, P3_ADD_526_U37, P3_ADD_526_U38, P3_ADD_526_U39, P3_ADD_526_U40, P3_ADD_526_U41, P3_ADD_526_U42, P3_ADD_526_U43, P3_ADD_526_U44, P3_ADD_526_U45, P3_ADD_526_U46, P3_ADD_526_U47, P3_ADD_526_U48, P3_ADD_526_U49, P3_ADD_526_U50, P3_ADD_526_U51, P3_ADD_526_U52, P3_ADD_526_U53, P3_ADD_526_U54, P3_ADD_526_U55, P3_ADD_526_U56, P3_ADD_526_U57, P3_ADD_526_U58, P3_ADD_526_U59, P3_ADD_526_U60, P3_ADD_526_U61, P3_ADD_526_U62, P3_ADD_526_U63, P3_ADD_526_U64, P3_ADD_526_U65, P3_ADD_526_U66, P3_ADD_526_U67, P3_ADD_526_U68, P3_ADD_526_U69, P3_ADD_526_U70, P3_ADD_526_U71, P3_ADD_526_U72, P3_ADD_526_U73, P3_ADD_526_U74, P3_ADD_526_U75, P3_ADD_526_U76, P3_ADD_526_U77, P3_ADD_526_U78, P3_ADD_526_U79, P3_ADD_526_U80, P3_ADD_526_U81, P3_ADD_526_U82, P3_ADD_526_U83, P3_ADD_526_U84, P3_ADD_526_U85, P3_ADD_526_U86, P3_ADD_526_U87, P3_ADD_526_U88, P3_ADD_526_U89, P3_ADD_526_U90, P3_ADD_526_U91, P3_ADD_526_U92, P3_ADD_526_U93, P3_ADD_526_U94, P3_ADD_526_U95, P3_ADD_526_U96, P3_ADD_526_U97, P3_ADD_526_U98, P3_ADD_526_U99, P3_ADD_526_U100, P3_ADD_526_U101, P3_ADD_526_U102, P3_ADD_526_U103, P3_ADD_526_U104, P3_ADD_526_U105, P3_ADD_526_U106, P3_ADD_526_U107, P3_ADD_526_U108, P3_ADD_526_U109, P3_ADD_526_U110, P3_ADD_526_U111, P3_ADD_526_U112, P3_ADD_526_U113, P3_ADD_526_U114, P3_ADD_526_U115, P3_ADD_526_U116, P3_ADD_526_U117, P3_ADD_526_U118, P3_ADD_526_U119, P3_ADD_526_U120, P3_ADD_526_U121, P3_ADD_526_U122, P3_ADD_526_U123, P3_ADD_526_U124, P3_ADD_526_U125, P3_ADD_526_U126, P3_ADD_526_U127, P3_ADD_526_U128, P3_ADD_526_U129, P3_ADD_526_U130, P3_ADD_526_U131, P3_ADD_526_U132, P3_ADD_526_U133, P3_ADD_526_U134, P3_ADD_526_U135, P3_ADD_526_U136, P3_ADD_526_U137, P3_ADD_526_U138, P3_ADD_526_U139, P3_ADD_526_U140, P3_ADD_526_U141, P3_ADD_526_U142, P3_ADD_526_U143, P3_ADD_526_U144, P3_ADD_526_U145, P3_ADD_526_U146, P3_ADD_526_U147, P3_ADD_526_U148, P3_ADD_526_U149, P3_ADD_526_U150, P3_ADD_526_U151, P3_ADD_526_U152, P3_ADD_526_U153, P3_ADD_526_U154, P3_ADD_526_U155, P3_ADD_526_U156, P3_ADD_526_U157, P3_ADD_526_U158, P3_ADD_526_U159, P3_ADD_526_U160, P3_ADD_526_U161, P3_ADD_526_U162, P3_ADD_526_U163, P3_ADD_526_U164, P3_ADD_526_U165, P3_ADD_526_U166, P3_ADD_526_U167, P3_ADD_526_U168, P3_ADD_526_U169, P3_ADD_526_U170, P3_ADD_526_U171, P3_ADD_526_U172, P3_ADD_526_U173, P3_ADD_526_U174, P3_ADD_526_U175, P3_ADD_526_U176, P3_ADD_526_U177, P3_ADD_526_U178, P3_ADD_526_U179, P3_ADD_526_U180, P3_ADD_526_U181, P3_ADD_526_U182, P3_ADD_526_U183, P3_ADD_526_U184, P3_ADD_526_U185, P3_ADD_526_U186, P3_ADD_526_U187, P3_ADD_526_U188, P3_ADD_526_U189, P3_ADD_526_U190, P3_ADD_526_U191, P3_ADD_526_U192, P3_ADD_526_U193, P3_ADD_526_U194, P3_ADD_526_U195, P3_ADD_526_U196, P3_ADD_526_U197, P3_ADD_526_U198, P3_ADD_526_U199, P3_ADD_526_U200, P3_ADD_526_U201, P3_ADD_526_U202, P3_ADD_552_U5, P3_ADD_552_U6, P3_ADD_552_U7, P3_ADD_552_U8, P3_ADD_552_U9, P3_ADD_552_U10, P3_ADD_552_U11, P3_ADD_552_U12, P3_ADD_552_U13, P3_ADD_552_U14, P3_ADD_552_U15, P3_ADD_552_U16, P3_ADD_552_U17, P3_ADD_552_U18, P3_ADD_552_U19, P3_ADD_552_U20, P3_ADD_552_U21, P3_ADD_552_U22, P3_ADD_552_U23, P3_ADD_552_U24, P3_ADD_552_U25, P3_ADD_552_U26, P3_ADD_552_U27, P3_ADD_552_U28, P3_ADD_552_U29, P3_ADD_552_U30, P3_ADD_552_U31, P3_ADD_552_U32, P3_ADD_552_U33, P3_ADD_552_U34, P3_ADD_552_U35, P3_ADD_552_U36, P3_ADD_552_U37, P3_ADD_552_U38, P3_ADD_552_U39, P3_ADD_552_U40, P3_ADD_552_U41, P3_ADD_552_U42, P3_ADD_552_U43, P3_ADD_552_U44, P3_ADD_552_U45, P3_ADD_552_U46, P3_ADD_552_U47, P3_ADD_552_U48, P3_ADD_552_U49, P3_ADD_552_U50, P3_ADD_552_U51, P3_ADD_552_U52, P3_ADD_552_U53, P3_ADD_552_U54, P3_ADD_552_U55, P3_ADD_552_U56, P3_ADD_552_U57, P3_ADD_552_U58, P3_ADD_552_U59, P3_ADD_552_U60, P3_ADD_552_U61, P3_ADD_552_U62, P3_ADD_552_U63, P3_ADD_552_U64, P3_ADD_552_U65, P3_ADD_552_U66, P3_ADD_552_U67, P3_ADD_552_U68, P3_ADD_552_U69, P3_ADD_552_U70, P3_ADD_552_U71, P3_ADD_552_U72, P3_ADD_552_U73, P3_ADD_552_U74, P3_ADD_552_U75, P3_ADD_552_U76, P3_ADD_552_U77, P3_ADD_552_U78, P3_ADD_552_U79, P3_ADD_552_U80, P3_ADD_552_U81, P3_ADD_552_U82, P3_ADD_552_U83, P3_ADD_552_U84, P3_ADD_552_U85, P3_ADD_552_U86, P3_ADD_552_U87, P3_ADD_552_U88, P3_ADD_552_U89, P3_ADD_552_U90, P3_ADD_552_U91, P3_ADD_552_U92, P3_ADD_552_U93, P3_ADD_552_U94, P3_ADD_552_U95, P3_ADD_552_U96, P3_ADD_552_U97, P3_ADD_552_U98, P3_ADD_552_U99, P3_ADD_552_U100, P3_ADD_552_U101, P3_ADD_552_U102, P3_ADD_552_U103, P3_ADD_552_U104, P3_ADD_552_U105, P3_ADD_552_U106, P3_ADD_552_U107, P3_ADD_552_U108, P3_ADD_552_U109, P3_ADD_552_U110, P3_ADD_552_U111, P3_ADD_552_U112, P3_ADD_552_U113, P3_ADD_552_U114, P3_ADD_552_U115, P3_ADD_552_U116, P3_ADD_552_U117, P3_ADD_552_U118, P3_ADD_552_U119, P3_ADD_552_U120, P3_ADD_552_U121, P3_ADD_552_U122, P3_ADD_552_U123, P3_ADD_552_U124, P3_ADD_552_U125, P3_ADD_552_U126, P3_ADD_552_U127, P3_ADD_552_U128, P3_ADD_552_U129, P3_ADD_552_U130, P3_ADD_552_U131, P3_ADD_552_U132, P3_ADD_552_U133, P3_ADD_552_U134, P3_ADD_552_U135, P3_ADD_552_U136, P3_ADD_552_U137, P3_ADD_552_U138, P3_ADD_552_U139, P3_ADD_552_U140, P3_ADD_552_U141, P3_ADD_552_U142, P3_ADD_552_U143, P3_ADD_552_U144, P3_ADD_552_U145, P3_ADD_552_U146, P3_ADD_552_U147, P3_ADD_552_U148, P3_ADD_552_U149, P3_ADD_552_U150, P3_ADD_552_U151, P3_ADD_552_U152, P3_ADD_552_U153, P3_ADD_552_U154, P3_ADD_552_U155, P3_ADD_552_U156, P3_ADD_552_U157, P3_ADD_552_U158, P3_ADD_552_U159, P3_ADD_552_U160, P3_ADD_552_U161, P3_ADD_552_U162, P3_ADD_552_U163, P3_ADD_552_U164, P3_ADD_552_U165, P3_ADD_552_U166, P3_ADD_552_U167, P3_ADD_552_U168, P3_ADD_552_U169, P3_ADD_552_U170, P3_ADD_552_U171, P3_ADD_552_U172, P3_ADD_552_U173, P3_ADD_552_U174, P3_ADD_552_U175, P3_ADD_552_U176, P3_ADD_552_U177, P3_ADD_552_U178, P3_ADD_552_U179, P3_ADD_552_U180, P3_ADD_552_U181, P3_ADD_552_U182, P3_ADD_552_U183, P3_ADD_552_U184, P3_ADD_552_U185, P3_ADD_552_U186, P3_ADD_552_U187, P3_ADD_552_U188, P3_ADD_552_U189, P3_ADD_552_U190, P3_ADD_552_U191, P3_ADD_552_U192, P3_ADD_552_U193, P3_ADD_552_U194, P3_ADD_552_U195, P3_ADD_552_U196, P3_ADD_552_U197, P3_ADD_552_U198, P3_ADD_552_U199, P3_ADD_552_U200, P3_ADD_552_U201, P3_ADD_552_U202, P3_ADD_546_U5, P3_ADD_546_U6, P3_ADD_546_U7, P3_ADD_546_U8, P3_ADD_546_U9, P3_ADD_546_U10, P3_ADD_546_U11, P3_ADD_546_U12, P3_ADD_546_U13, P3_ADD_546_U14, P3_ADD_546_U15, P3_ADD_546_U16, P3_ADD_546_U17, P3_ADD_546_U18, P3_ADD_546_U19, P3_ADD_546_U20, P3_ADD_546_U21, P3_ADD_546_U22, P3_ADD_546_U23, P3_ADD_546_U24, P3_ADD_546_U25, P3_ADD_546_U26, P3_ADD_546_U27, P3_ADD_546_U28, P3_ADD_546_U29, P3_ADD_546_U30, P3_ADD_546_U31, P3_ADD_546_U32, P3_ADD_546_U33, P3_ADD_546_U34, P3_ADD_546_U35, P3_ADD_546_U36, P3_ADD_546_U37, P3_ADD_546_U38, P3_ADD_546_U39, P3_ADD_546_U40, P3_ADD_546_U41, P3_ADD_546_U42, P3_ADD_546_U43, P3_ADD_546_U44, P3_ADD_546_U45, P3_ADD_546_U46, P3_ADD_546_U47, P3_ADD_546_U48, P3_ADD_546_U49, P3_ADD_546_U50, P3_ADD_546_U51, P3_ADD_546_U52, P3_ADD_546_U53, P3_ADD_546_U54, P3_ADD_546_U55, P3_ADD_546_U56, P3_ADD_546_U57, P3_ADD_546_U58, P3_ADD_546_U59, P3_ADD_546_U60, P3_ADD_546_U61, P3_ADD_546_U62, P3_ADD_546_U63, P3_ADD_546_U64, P3_ADD_546_U65, P3_ADD_546_U66, P3_ADD_546_U67, P3_ADD_546_U68, P3_ADD_546_U69, P3_ADD_546_U70, P3_ADD_546_U71, P3_ADD_546_U72, P3_ADD_546_U73, P3_ADD_546_U74, P3_ADD_546_U75, P3_ADD_546_U76, P3_ADD_546_U77, P3_ADD_546_U78, P3_ADD_546_U79, P3_ADD_546_U80, P3_ADD_546_U81, P3_ADD_546_U82, P3_ADD_546_U83, P3_ADD_546_U84, P3_ADD_546_U85, P3_ADD_546_U86, P3_ADD_546_U87, P3_ADD_546_U88, P3_ADD_546_U89, P3_ADD_546_U90, P3_ADD_546_U91, P3_ADD_546_U92, P3_ADD_546_U93, P3_ADD_546_U94, P3_ADD_546_U95, P3_ADD_546_U96, P3_ADD_546_U97, P3_ADD_546_U98, P3_ADD_546_U99, P3_ADD_546_U100, P3_ADD_546_U101, P3_ADD_546_U102, P3_ADD_546_U103, P3_ADD_546_U104, P3_ADD_546_U105, P3_ADD_546_U106, P3_ADD_546_U107, P3_ADD_546_U108, P3_ADD_546_U109, P3_ADD_546_U110, P3_ADD_546_U111, P3_ADD_546_U112, P3_ADD_546_U113, P3_ADD_546_U114, P3_ADD_546_U115, P3_ADD_546_U116, P3_ADD_546_U117, P3_ADD_546_U118, P3_ADD_546_U119, P3_ADD_546_U120, P3_ADD_546_U121, P3_ADD_546_U122, P3_ADD_546_U123, P3_ADD_546_U124, P3_ADD_546_U125, P3_ADD_546_U126, P3_ADD_546_U127, P3_ADD_546_U128, P3_ADD_546_U129, P3_ADD_546_U130, P3_ADD_546_U131, P3_ADD_546_U132, P3_ADD_546_U133, P3_ADD_546_U134, P3_ADD_546_U135, P3_ADD_546_U136, P3_ADD_546_U137, P3_ADD_546_U138, P3_ADD_546_U139, P3_ADD_546_U140, P3_ADD_546_U141, P3_ADD_546_U142, P3_ADD_546_U143, P3_ADD_546_U144, P3_ADD_546_U145, P3_ADD_546_U146, P3_ADD_546_U147, P3_ADD_546_U148, P3_ADD_546_U149, P3_ADD_546_U150, P3_ADD_546_U151, P3_ADD_546_U152, P3_ADD_546_U153, P3_ADD_546_U154, P3_ADD_546_U155, P3_ADD_546_U156, P3_ADD_546_U157, P3_ADD_546_U158, P3_ADD_546_U159, P3_ADD_546_U160, P3_ADD_546_U161, P3_ADD_546_U162, P3_ADD_546_U163, P3_ADD_546_U164, P3_ADD_546_U165, P3_ADD_546_U166, P3_ADD_546_U167, P3_ADD_546_U168, P3_ADD_546_U169, P3_ADD_546_U170, P3_ADD_546_U171, P3_ADD_546_U172, P3_ADD_546_U173, P3_ADD_546_U174, P3_ADD_546_U175, P3_ADD_546_U176, P3_ADD_546_U177, P3_ADD_546_U178, P3_ADD_546_U179, P3_ADD_546_U180, P3_ADD_546_U181, P3_ADD_546_U182, P3_ADD_546_U183, P3_ADD_546_U184, P3_ADD_546_U185, P3_ADD_546_U186, P3_ADD_546_U187, P3_ADD_546_U188, P3_ADD_546_U189, P3_ADD_546_U190, P3_ADD_546_U191, P3_ADD_546_U192, P3_ADD_546_U193, P3_ADD_546_U194, P3_ADD_546_U195, P3_ADD_546_U196, P3_ADD_546_U197, P3_ADD_546_U198, P3_ADD_546_U199, P3_ADD_546_U200, P3_ADD_546_U201, P3_ADD_546_U202, P3_GTE_401_U6, P3_GTE_401_U7, P3_GTE_401_U8, P3_GTE_401_U9, P3_ADD_391_1180_U4, P3_ADD_391_1180_U5, P3_ADD_391_1180_U6, P3_ADD_391_1180_U7, P3_ADD_391_1180_U8, P3_ADD_391_1180_U9, P3_ADD_391_1180_U10, P3_ADD_391_1180_U11, P3_ADD_391_1180_U12, P3_ADD_391_1180_U13, P3_ADD_391_1180_U14, P3_ADD_391_1180_U15, P3_ADD_391_1180_U16, P3_ADD_391_1180_U17, P3_ADD_391_1180_U18, P3_ADD_391_1180_U19, P3_ADD_391_1180_U20, P3_ADD_391_1180_U21, P3_ADD_391_1180_U22, P3_ADD_391_1180_U23, P3_ADD_391_1180_U24, P3_ADD_391_1180_U25, P3_ADD_391_1180_U26, P3_ADD_391_1180_U27, P3_ADD_391_1180_U28, P3_ADD_391_1180_U29, P3_ADD_391_1180_U30, P3_ADD_391_1180_U31, P3_ADD_391_1180_U32, P3_ADD_391_1180_U33, P3_ADD_391_1180_U34, P3_ADD_391_1180_U35, P3_ADD_391_1180_U36, P3_ADD_391_1180_U37, P3_ADD_391_1180_U38, P3_ADD_391_1180_U39, P3_ADD_391_1180_U40, P3_ADD_391_1180_U41, P3_ADD_391_1180_U42, P3_ADD_391_1180_U43, P3_ADD_391_1180_U44, P3_ADD_391_1180_U45, P3_ADD_391_1180_U46, P3_ADD_391_1180_U47, P3_ADD_391_1180_U48, P3_ADD_391_1180_U49, P3_ADD_391_1180_U50, P3_ADD_476_U4, P3_ADD_476_U5, P3_ADD_476_U6, P3_ADD_476_U7, P3_ADD_476_U8, P3_ADD_476_U9, P3_ADD_476_U10, P3_ADD_476_U11, P3_ADD_476_U12, P3_ADD_476_U13, P3_ADD_476_U14, P3_ADD_476_U15, P3_ADD_476_U16, P3_ADD_476_U17, P3_ADD_476_U18, P3_ADD_476_U19, P3_ADD_476_U20, P3_ADD_476_U21, P3_ADD_476_U22, P3_ADD_476_U23, P3_ADD_476_U24, P3_ADD_476_U25, P3_ADD_476_U26, P3_ADD_476_U27, P3_ADD_476_U28, P3_ADD_476_U29, P3_ADD_476_U30, P3_ADD_476_U31, P3_ADD_476_U32, P3_ADD_476_U33, P3_ADD_476_U34, P3_ADD_476_U35, P3_ADD_476_U36, P3_ADD_476_U37, P3_ADD_476_U38, P3_ADD_476_U39, P3_ADD_476_U40, P3_ADD_476_U41, P3_ADD_476_U42, P3_ADD_476_U43, P3_ADD_476_U44, P3_ADD_476_U45, P3_ADD_476_U46, P3_ADD_476_U47, P3_ADD_476_U48, P3_ADD_476_U49, P3_ADD_476_U50, P3_ADD_476_U51, P3_ADD_476_U52, P3_ADD_476_U53, P3_ADD_476_U54, P3_ADD_476_U55, P3_ADD_476_U56, P3_ADD_476_U57, P3_ADD_476_U58, P3_ADD_476_U59, P3_ADD_476_U60, P3_ADD_476_U61, P3_ADD_476_U62, P3_ADD_476_U63, P3_ADD_476_U64, P3_ADD_476_U65, P3_ADD_476_U66, P3_ADD_476_U67, P3_ADD_476_U68, P3_ADD_476_U69, P3_ADD_476_U70, P3_ADD_476_U71, P3_ADD_476_U72, P3_ADD_476_U73, P3_ADD_476_U74, P3_ADD_476_U75, P3_ADD_476_U76, P3_ADD_476_U77, P3_ADD_476_U78, P3_ADD_476_U79, P3_ADD_476_U80, P3_ADD_476_U81, P3_ADD_476_U82, P3_ADD_476_U83, P3_ADD_476_U84, P3_ADD_476_U85, P3_ADD_476_U86, P3_ADD_476_U87, P3_ADD_476_U88, P3_ADD_476_U89, P3_ADD_476_U90, P3_ADD_476_U91, P3_ADD_476_U92, P3_ADD_476_U93, P3_ADD_476_U94, P3_ADD_476_U95, P3_ADD_476_U96, P3_ADD_476_U97, P3_ADD_476_U98, P3_ADD_476_U99, P3_ADD_476_U100, P3_ADD_476_U101, P3_ADD_476_U102, P3_ADD_476_U103, P3_ADD_476_U104, P3_ADD_476_U105, P3_ADD_476_U106, P3_ADD_476_U107, P3_ADD_476_U108, P3_ADD_476_U109, P3_ADD_476_U110, P3_ADD_476_U111, P3_ADD_476_U112, P3_ADD_476_U113, P3_ADD_476_U114, P3_ADD_476_U115, P3_ADD_476_U116, P3_ADD_476_U117, P3_ADD_476_U118, P3_ADD_476_U119, P3_ADD_476_U120, P3_ADD_476_U121, P3_ADD_476_U122, P3_ADD_476_U123, P3_ADD_476_U124, P3_ADD_476_U125, P3_ADD_476_U126, P3_ADD_476_U127, P3_ADD_476_U128, P3_ADD_476_U129, P3_ADD_476_U130, P3_ADD_476_U131, P3_ADD_476_U132, P3_ADD_476_U133, P3_ADD_476_U134, P3_ADD_476_U135, P3_ADD_476_U136, P3_ADD_476_U137, P3_ADD_476_U138, P3_ADD_476_U139, P3_ADD_476_U140, P3_ADD_476_U141, P3_ADD_476_U142, P3_ADD_476_U143, P3_ADD_476_U144, P3_ADD_476_U145, P3_ADD_476_U146, P3_ADD_476_U147, P3_ADD_476_U148, P3_ADD_476_U149, P3_ADD_476_U150, P3_ADD_476_U151, P3_ADD_476_U152, P3_ADD_476_U153, P3_ADD_476_U154, P3_ADD_476_U155, P3_ADD_476_U156, P3_ADD_476_U157, P3_ADD_476_U158, P3_ADD_476_U159, P3_ADD_476_U160, P3_ADD_476_U161, P3_ADD_476_U162, P3_ADD_476_U163, P3_ADD_476_U164, P3_ADD_476_U165, P3_ADD_476_U166, P3_ADD_476_U167, P3_ADD_476_U168, P3_ADD_476_U169, P3_ADD_476_U170, P3_ADD_476_U171, P3_ADD_476_U172, P3_ADD_476_U173, P3_ADD_476_U174, P3_ADD_476_U175, P3_ADD_476_U176, P3_ADD_476_U177, P3_ADD_476_U178, P3_ADD_476_U179, P3_ADD_476_U180, P3_ADD_476_U181, P3_ADD_476_U182, P3_GTE_390_U6, P3_GTE_390_U7, P3_GTE_390_U8, P3_GTE_390_U9, P3_ADD_531_U5, P3_ADD_531_U6, P3_ADD_531_U7, P3_ADD_531_U8, P3_ADD_531_U9, P3_ADD_531_U10, P3_ADD_531_U11, P3_ADD_531_U12, P3_ADD_531_U13, P3_ADD_531_U14, P3_ADD_531_U15, P3_ADD_531_U16, P3_ADD_531_U17, P3_ADD_531_U18, P3_ADD_531_U19, P3_ADD_531_U20, P3_ADD_531_U21, P3_ADD_531_U22, P3_ADD_531_U23, P3_ADD_531_U24, P3_ADD_531_U25, P3_ADD_531_U26, P3_ADD_531_U27, P3_ADD_531_U28, P3_ADD_531_U29, P3_ADD_531_U30, P3_ADD_531_U31, P3_ADD_531_U32, P3_ADD_531_U33, P3_ADD_531_U34, P3_ADD_531_U35, P3_ADD_531_U36, P3_ADD_531_U37, P3_ADD_531_U38, P3_ADD_531_U39, P3_ADD_531_U40, P3_ADD_531_U41, P3_ADD_531_U42, P3_ADD_531_U43, P3_ADD_531_U44, P3_ADD_531_U45, P3_ADD_531_U46, P3_ADD_531_U47, P3_ADD_531_U48, P3_ADD_531_U49, P3_ADD_531_U50, P3_ADD_531_U51, P3_ADD_531_U52, P3_ADD_531_U53, P3_ADD_531_U54, P3_ADD_531_U55, P3_ADD_531_U56, P3_ADD_531_U57, P3_ADD_531_U58, P3_ADD_531_U59, P3_ADD_531_U60, P3_ADD_531_U61, P3_ADD_531_U62, P3_ADD_531_U63, P3_ADD_531_U64, P3_ADD_531_U65, P3_ADD_531_U66, P3_ADD_531_U67, P3_ADD_531_U68, P3_ADD_531_U69, P3_ADD_531_U70, P3_ADD_531_U71, P3_ADD_531_U72, P3_ADD_531_U73, P3_ADD_531_U74, P3_ADD_531_U75, P3_ADD_531_U76, P3_ADD_531_U77, P3_ADD_531_U78, P3_ADD_531_U79, P3_ADD_531_U80, P3_ADD_531_U81, P3_ADD_531_U82, P3_ADD_531_U83, P3_ADD_531_U84, P3_ADD_531_U85, P3_ADD_531_U86, P3_ADD_531_U87, P3_ADD_531_U88, P3_ADD_531_U89, P3_ADD_531_U90, P3_ADD_531_U91, P3_ADD_531_U92, P3_ADD_531_U93, P3_ADD_531_U94, P3_ADD_531_U95, P3_ADD_531_U96, P3_ADD_531_U97, P3_ADD_531_U98, P3_ADD_531_U99, P3_ADD_531_U100, P3_ADD_531_U101, P3_ADD_531_U102, P3_ADD_531_U103, P3_ADD_531_U104, P3_ADD_531_U105, P3_ADD_531_U106, P3_ADD_531_U107, P3_ADD_531_U108, P3_ADD_531_U109, P3_ADD_531_U110, P3_ADD_531_U111, P3_ADD_531_U112, P3_ADD_531_U113, P3_ADD_531_U114, P3_ADD_531_U115, P3_ADD_531_U116, P3_ADD_531_U117, P3_ADD_531_U118, P3_ADD_531_U119, P3_ADD_531_U120, P3_ADD_531_U121, P3_ADD_531_U122, P3_ADD_531_U123, P3_ADD_531_U124, P3_ADD_531_U125, P3_ADD_531_U126, P3_ADD_531_U127, P3_ADD_531_U128, P3_ADD_531_U129, P3_ADD_531_U130, P3_ADD_531_U131, P3_ADD_531_U132, P3_ADD_531_U133, P3_ADD_531_U134, P3_ADD_531_U135, P3_ADD_531_U136, P3_ADD_531_U137, P3_ADD_531_U138, P3_ADD_531_U139, P3_ADD_531_U140, P3_ADD_531_U141, P3_ADD_531_U142, P3_ADD_531_U143, P3_ADD_531_U144, P3_ADD_531_U145, P3_ADD_531_U146, P3_ADD_531_U147, P3_ADD_531_U148, P3_ADD_531_U149, P3_ADD_531_U150, P3_ADD_531_U151, P3_ADD_531_U152, P3_ADD_531_U153, P3_ADD_531_U154, P3_ADD_531_U155, P3_ADD_531_U156, P3_ADD_531_U157, P3_ADD_531_U158, P3_ADD_531_U159, P3_ADD_531_U160, P3_ADD_531_U161, P3_ADD_531_U162, P3_ADD_531_U163, P3_ADD_531_U164, P3_ADD_531_U165, P3_ADD_531_U166, P3_ADD_531_U167, P3_ADD_531_U168, P3_ADD_531_U169, P3_ADD_531_U170, P3_ADD_531_U171, P3_ADD_531_U172, P3_ADD_531_U173, P3_ADD_531_U174, P3_ADD_531_U175, P3_ADD_531_U176, P3_ADD_531_U177, P3_ADD_531_U178, P3_ADD_531_U179, P3_ADD_531_U180, P3_ADD_531_U181, P3_ADD_531_U182, P3_ADD_531_U183, P3_ADD_531_U184, P3_ADD_531_U185, P3_ADD_531_U186, P3_ADD_531_U187, P3_ADD_531_U188, P3_ADD_531_U189, P3_SUB_320_U6, P3_SUB_320_U7, P3_SUB_320_U8, P3_SUB_320_U9, P3_SUB_320_U10, P3_SUB_320_U11, P3_SUB_320_U12, P3_SUB_320_U13, P3_SUB_320_U14, P3_SUB_320_U15, P3_SUB_320_U16, P3_SUB_320_U17, P3_SUB_320_U18, P3_SUB_320_U19, P3_SUB_320_U20, P3_SUB_320_U21, P3_SUB_320_U22, P3_SUB_320_U23, P3_SUB_320_U24, P3_SUB_320_U25, P3_SUB_320_U26, P3_SUB_320_U27, P3_SUB_320_U28, P3_SUB_320_U29, P3_SUB_320_U30, P3_SUB_320_U31, P3_SUB_320_U32, P3_SUB_320_U33, P3_SUB_320_U34, P3_SUB_320_U35, P3_SUB_320_U36, P3_SUB_320_U37, P3_SUB_320_U38, P3_SUB_320_U39, P3_SUB_320_U40, P3_SUB_320_U41, P3_SUB_320_U42, P3_SUB_320_U43, P3_SUB_320_U44, P3_SUB_320_U45, P3_SUB_320_U46, P3_SUB_320_U47, P3_SUB_320_U48, P3_SUB_320_U49, P3_SUB_320_U50, P3_SUB_320_U51, P3_SUB_320_U52, P3_SUB_320_U53, P3_SUB_320_U54, P3_SUB_320_U55, P3_SUB_320_U56, P3_SUB_320_U57, P3_SUB_320_U58, P3_SUB_320_U59, P3_SUB_320_U60, P3_SUB_320_U61, P3_SUB_320_U62, P3_SUB_320_U63, P3_SUB_320_U64, P3_SUB_320_U65, P3_SUB_320_U66, P3_SUB_320_U67, P3_SUB_320_U68, P3_SUB_320_U69, P3_SUB_320_U70, P3_SUB_320_U71, P3_SUB_320_U72, P3_SUB_320_U73, P3_SUB_320_U74, P3_SUB_320_U75, P3_SUB_320_U76, P3_SUB_320_U77, P3_SUB_320_U78, P3_SUB_320_U79, P3_SUB_320_U80, P3_SUB_320_U81, P3_SUB_320_U82, P3_SUB_320_U83, P3_SUB_320_U84, P3_SUB_320_U85, P3_SUB_320_U86, P3_SUB_320_U87, P3_SUB_320_U88, P3_SUB_320_U89, P3_SUB_320_U90, P3_SUB_320_U91, P3_SUB_320_U92, P3_SUB_320_U93, P3_SUB_320_U94, P3_SUB_320_U95, P3_SUB_320_U96, P3_SUB_320_U97, P3_SUB_320_U98, P3_SUB_320_U99, P3_SUB_320_U100, P3_SUB_320_U101, P3_SUB_320_U102, P3_SUB_320_U103, P3_SUB_320_U104, P3_SUB_320_U105, P3_SUB_320_U106, P3_SUB_320_U107, P3_SUB_320_U108, P3_SUB_320_U109, P3_SUB_320_U110, P3_SUB_320_U111, P3_SUB_320_U112, P3_SUB_320_U113, P3_SUB_320_U114, P3_SUB_320_U115, P3_SUB_320_U116, P3_SUB_320_U117, P3_SUB_320_U118, P3_SUB_320_U119, P3_SUB_320_U120, P3_SUB_320_U121, P3_SUB_320_U122, P3_SUB_320_U123, P3_SUB_320_U124, P3_SUB_320_U125, P3_SUB_320_U126, P3_SUB_320_U127, P3_SUB_320_U128, P3_SUB_320_U129, P3_SUB_320_U130, P3_SUB_320_U131, P3_SUB_320_U132, P3_SUB_320_U133, P3_SUB_320_U134, P3_SUB_320_U135, P3_SUB_320_U136, P3_SUB_320_U137, P3_SUB_320_U138, P3_SUB_320_U139, P3_SUB_320_U140, P3_SUB_320_U141, P3_SUB_320_U142, P3_SUB_320_U143, P3_SUB_320_U144, P3_SUB_320_U145, P3_SUB_320_U146, P3_SUB_320_U147, P3_SUB_320_U148, P3_SUB_320_U149, P3_SUB_320_U150, P3_SUB_320_U151, P3_SUB_320_U152, P3_SUB_320_U153, P3_SUB_320_U154, P3_SUB_320_U155, P3_SUB_320_U156, P3_SUB_320_U157, P3_SUB_320_U158, P3_SUB_320_U159, P3_ADD_505_U5, P3_ADD_505_U6, P3_ADD_505_U7, P3_ADD_505_U8, P3_ADD_505_U9, P3_ADD_505_U10, P3_ADD_505_U11, P3_ADD_505_U12, P3_ADD_505_U13, P3_ADD_505_U14, P3_ADD_505_U15, P3_ADD_505_U16, P3_ADD_505_U17, P3_ADD_505_U18, P3_ADD_505_U19, P3_ADD_505_U20, P3_ADD_505_U21, P3_ADD_505_U22, P3_ADD_505_U23, P3_ADD_505_U24, P3_ADD_505_U25, P3_ADD_505_U26, P3_ADD_505_U27, P3_ADD_505_U28, P3_GTE_485_U6, P3_GTE_485_U7, P3_ADD_318_U4, P3_ADD_318_U5, P3_ADD_318_U6, P3_ADD_318_U7, P3_ADD_318_U8, P3_ADD_318_U9, P3_ADD_318_U10, P3_ADD_318_U11, P3_ADD_318_U12, P3_ADD_318_U13, P3_ADD_318_U14, P3_ADD_318_U15, P3_ADD_318_U16, P3_ADD_318_U17, P3_ADD_318_U18, P3_ADD_318_U19, P3_ADD_318_U20, P3_ADD_318_U21, P3_ADD_318_U22, P3_ADD_318_U23, P3_ADD_318_U24, P3_ADD_318_U25, P3_ADD_318_U26, P3_ADD_318_U27, P3_ADD_318_U28, P3_ADD_318_U29, P3_ADD_318_U30, P3_ADD_318_U31, P3_ADD_318_U32, P3_ADD_318_U33, P3_ADD_318_U34, P3_ADD_318_U35, P3_ADD_318_U36, P3_ADD_318_U37, P3_ADD_318_U38, P3_ADD_318_U39, P3_ADD_318_U40, P3_ADD_318_U41, P3_ADD_318_U42, P3_ADD_318_U43, P3_ADD_318_U44, P3_ADD_318_U45, P3_ADD_318_U46, P3_ADD_318_U47, P3_ADD_318_U48, P3_ADD_318_U49, P3_ADD_318_U50, P3_ADD_318_U51, P3_ADD_318_U52, P3_ADD_318_U53, P3_ADD_318_U54, P3_ADD_318_U55, P3_ADD_318_U56, P3_ADD_318_U57, P3_ADD_318_U58, P3_ADD_318_U59, P3_ADD_318_U60, P3_ADD_318_U61, P3_ADD_318_U62, P3_ADD_318_U63, P3_ADD_318_U64, P3_ADD_318_U65, P3_ADD_318_U66, P3_ADD_318_U67, P3_ADD_318_U68, P3_ADD_318_U69, P3_ADD_318_U70, P3_ADD_318_U71, P3_ADD_318_U72, P3_ADD_318_U73, P3_ADD_318_U74, P3_ADD_318_U75, P3_ADD_318_U76, P3_ADD_318_U77, P3_ADD_318_U78, P3_ADD_318_U79, P3_ADD_318_U80, P3_ADD_318_U81, P3_ADD_318_U82, P3_ADD_318_U83, P3_ADD_318_U84, P3_ADD_318_U85, P3_ADD_318_U86, P3_ADD_318_U87, P3_ADD_318_U88, P3_ADD_318_U89, P3_ADD_318_U90, P3_ADD_318_U91, P3_ADD_318_U92, P3_ADD_318_U93, P3_ADD_318_U94, P3_ADD_318_U95, P3_ADD_318_U96, P3_ADD_318_U97, P3_ADD_318_U98, P3_ADD_318_U99, P3_ADD_318_U100, P3_ADD_318_U101, P3_ADD_318_U102, P3_ADD_318_U103, P3_ADD_318_U104, P3_ADD_318_U105, P3_ADD_318_U106, P3_ADD_318_U107, P3_ADD_318_U108, P3_ADD_318_U109, P3_ADD_318_U110, P3_ADD_318_U111, P3_ADD_318_U112, P3_ADD_318_U113, P3_ADD_318_U114, P3_ADD_318_U115, P3_ADD_318_U116, P3_ADD_318_U117, P3_ADD_318_U118, P3_ADD_318_U119, P3_ADD_318_U120, P3_ADD_318_U121, P3_ADD_318_U122, P3_ADD_318_U123, P3_ADD_318_U124, P3_ADD_318_U125, P3_ADD_318_U126, P3_ADD_318_U127, P3_ADD_318_U128, P3_ADD_318_U129, P3_ADD_318_U130, P3_ADD_318_U131, P3_ADD_318_U132, P3_ADD_318_U133, P3_ADD_318_U134, P3_ADD_318_U135, P3_ADD_318_U136, P3_ADD_318_U137, P3_ADD_318_U138, P3_ADD_318_U139, P3_ADD_318_U140, P3_ADD_318_U141, P3_ADD_318_U142, P3_ADD_318_U143, P3_ADD_318_U144, P3_ADD_318_U145, P3_ADD_318_U146, P3_ADD_318_U147, P3_ADD_318_U148, P3_ADD_318_U149, P3_ADD_318_U150, P3_ADD_318_U151, P3_ADD_318_U152, P3_ADD_318_U153, P3_ADD_318_U154, P3_ADD_318_U155, P3_ADD_318_U156, P3_ADD_318_U157, P3_ADD_318_U158, P3_ADD_318_U159, P3_ADD_318_U160, P3_ADD_318_U161, P3_ADD_318_U162, P3_ADD_318_U163, P3_ADD_318_U164, P3_ADD_318_U165, P3_ADD_318_U166, P3_ADD_318_U167, P3_ADD_318_U168, P3_ADD_318_U169, P3_ADD_318_U170, P3_ADD_318_U171, P3_ADD_318_U172, P3_ADD_318_U173, P3_ADD_318_U174, P3_ADD_318_U175, P3_ADD_318_U176, P3_ADD_318_U177, P3_ADD_318_U178, P3_ADD_318_U179, P3_ADD_318_U180, P3_ADD_318_U181, P3_ADD_318_U182, P3_SUB_370_U6, P3_SUB_370_U7, P3_SUB_370_U8, P3_SUB_370_U9, P3_SUB_370_U10, P3_SUB_370_U11, P3_SUB_370_U12, P3_SUB_370_U13, P3_SUB_370_U14, P3_SUB_370_U15, P3_SUB_370_U16, P3_SUB_370_U17, P3_SUB_370_U18, P3_SUB_370_U19, P3_SUB_370_U20, P3_SUB_370_U21, P3_SUB_370_U22, P3_SUB_370_U23, P3_SUB_370_U24, P3_SUB_370_U25, P3_SUB_370_U26, P3_SUB_370_U27, P3_SUB_370_U28, P3_SUB_370_U29, P3_SUB_370_U30, P3_SUB_370_U31, P3_SUB_370_U32, P3_SUB_370_U33, P3_SUB_370_U34, P3_SUB_370_U35, P3_SUB_370_U36, P3_SUB_370_U37, P3_SUB_370_U38, P3_SUB_370_U39, P3_SUB_370_U40, P3_SUB_370_U41, P3_SUB_370_U42, P3_SUB_370_U43, P3_SUB_370_U44, P3_SUB_370_U45, P3_SUB_370_U46, P3_SUB_370_U47, P3_SUB_370_U48, P3_SUB_370_U49, P3_SUB_370_U50, P3_SUB_370_U51, P3_SUB_370_U52, P3_SUB_370_U53, P3_SUB_370_U54, P3_SUB_370_U55, P3_SUB_370_U56, P3_SUB_370_U57, P3_SUB_370_U58, P3_SUB_370_U59, P3_SUB_370_U60, P3_SUB_370_U61, P3_SUB_370_U62, P3_SUB_370_U63, P3_SUB_370_U64, P3_SUB_370_U65, P3_SUB_370_U66, P3_ADD_315_U4, P3_ADD_315_U5, P3_ADD_315_U6, P3_ADD_315_U7, P3_ADD_315_U8, P3_ADD_315_U9, P3_ADD_315_U10, P3_ADD_315_U11, P3_ADD_315_U12, P3_ADD_315_U13, P3_ADD_315_U14, P3_ADD_315_U15, P3_ADD_315_U16, P3_ADD_315_U17, P3_ADD_315_U18, P3_ADD_315_U19, P3_ADD_315_U20, P3_ADD_315_U21, P3_ADD_315_U22, P3_ADD_315_U23, P3_ADD_315_U24, P3_ADD_315_U25, P3_ADD_315_U26, P3_ADD_315_U27, P3_ADD_315_U28, P3_ADD_315_U29, P3_ADD_315_U30, P3_ADD_315_U31, P3_ADD_315_U32, P3_ADD_315_U33, P3_ADD_315_U34, P3_ADD_315_U35, P3_ADD_315_U36, P3_ADD_315_U37, P3_ADD_315_U38, P3_ADD_315_U39, P3_ADD_315_U40, P3_ADD_315_U41, P3_ADD_315_U42, P3_ADD_315_U43, P3_ADD_315_U44, P3_ADD_315_U45, P3_ADD_315_U46, P3_ADD_315_U47, P3_ADD_315_U48, P3_ADD_315_U49, P3_ADD_315_U50, P3_ADD_315_U51, P3_ADD_315_U52, P3_ADD_315_U53, P3_ADD_315_U54, P3_ADD_315_U55, P3_ADD_315_U56, P3_ADD_315_U57, P3_ADD_315_U58, P3_ADD_315_U59, P3_ADD_315_U60, P3_ADD_315_U61, P3_ADD_315_U62, P3_ADD_315_U63, P3_ADD_315_U64, P3_ADD_315_U65, P3_ADD_315_U66, P3_ADD_315_U67, P3_ADD_315_U68, P3_ADD_315_U69, P3_ADD_315_U70, P3_ADD_315_U71, P3_ADD_315_U72, P3_ADD_315_U73, P3_ADD_315_U74, P3_ADD_315_U75, P3_ADD_315_U76, P3_ADD_315_U77, P3_ADD_315_U78, P3_ADD_315_U79, P3_ADD_315_U80, P3_ADD_315_U81, P3_ADD_315_U82, P3_ADD_315_U83, P3_ADD_315_U84, P3_ADD_315_U85, P3_ADD_315_U86, P3_ADD_315_U87, P3_ADD_315_U88, P3_ADD_315_U89, P3_ADD_315_U90, P3_ADD_315_U91, P3_ADD_315_U92, P3_ADD_315_U93, P3_ADD_315_U94, P3_ADD_315_U95, P3_ADD_315_U96, P3_ADD_315_U97, P3_ADD_315_U98, P3_ADD_315_U99, P3_ADD_315_U100, P3_ADD_315_U101, P3_ADD_315_U102, P3_ADD_315_U103, P3_ADD_315_U104, P3_ADD_315_U105, P3_ADD_315_U106, P3_ADD_315_U107, P3_ADD_315_U108, P3_ADD_315_U109, P3_ADD_315_U110, P3_ADD_315_U111, P3_ADD_315_U112, P3_ADD_315_U113, P3_ADD_315_U114, P3_ADD_315_U115, P3_ADD_315_U116, P3_ADD_315_U117, P3_ADD_315_U118, P3_ADD_315_U119, P3_ADD_315_U120, P3_ADD_315_U121, P3_ADD_315_U122, P3_ADD_315_U123, P3_ADD_315_U124, P3_ADD_315_U125, P3_ADD_315_U126, P3_ADD_315_U127, P3_ADD_315_U128, P3_ADD_315_U129, P3_ADD_315_U130, P3_ADD_315_U131, P3_ADD_315_U132, P3_ADD_315_U133, P3_ADD_315_U134, P3_ADD_315_U135, P3_ADD_315_U136, P3_ADD_315_U137, P3_ADD_315_U138, P3_ADD_315_U139, P3_ADD_315_U140, P3_ADD_315_U141, P3_ADD_315_U142, P3_ADD_315_U143, P3_ADD_315_U144, P3_ADD_315_U145, P3_ADD_315_U146, P3_ADD_315_U147, P3_ADD_315_U148, P3_ADD_315_U149, P3_ADD_315_U150, P3_ADD_315_U151, P3_ADD_315_U152, P3_ADD_315_U153, P3_ADD_315_U154, P3_ADD_315_U155, P3_ADD_315_U156, P3_ADD_315_U157, P3_ADD_315_U158, P3_ADD_315_U159, P3_ADD_315_U160, P3_ADD_315_U161, P3_ADD_315_U162, P3_ADD_315_U163, P3_ADD_315_U164, P3_ADD_315_U165, P3_ADD_315_U166, P3_ADD_315_U167, P3_ADD_315_U168, P3_ADD_315_U169, P3_ADD_315_U170, P3_ADD_315_U171, P3_ADD_315_U172, P3_ADD_315_U173, P3_ADD_315_U174, P3_ADD_315_U175, P3_ADD_315_U176, P3_GTE_355_U6, P3_GTE_355_U7, P3_GTE_355_U8, P3_ADD_360_1242_U4, P3_ADD_360_1242_U5, P3_ADD_360_1242_U6, P3_ADD_360_1242_U7, P3_ADD_360_1242_U8, P3_ADD_360_1242_U9, P3_ADD_360_1242_U10, P3_ADD_360_1242_U11, P3_ADD_360_1242_U12, P3_ADD_360_1242_U13, P3_ADD_360_1242_U14, P3_ADD_360_1242_U15, P3_ADD_360_1242_U16, P3_ADD_360_1242_U17, P3_ADD_360_1242_U18, P3_ADD_360_1242_U19, P3_ADD_360_1242_U20, P3_ADD_360_1242_U21, P3_ADD_360_1242_U22, P3_ADD_360_1242_U23, P3_ADD_360_1242_U24, P3_ADD_360_1242_U25, P3_ADD_360_1242_U26, P3_ADD_360_1242_U27, P3_ADD_360_1242_U28, P3_ADD_360_1242_U29, P3_ADD_360_1242_U30, P3_ADD_360_1242_U31, P3_ADD_360_1242_U32, P3_ADD_360_1242_U33, P3_ADD_360_1242_U34, P3_ADD_360_1242_U35, P3_ADD_360_1242_U36, P3_ADD_360_1242_U37, P3_ADD_360_1242_U38, P3_ADD_360_1242_U39, P3_ADD_360_1242_U40, P3_ADD_360_1242_U41, P3_ADD_360_1242_U42, P3_ADD_360_1242_U43, P3_ADD_360_1242_U44, P3_ADD_360_1242_U45, P3_ADD_360_1242_U46, P3_ADD_360_1242_U47, P3_ADD_360_1242_U48, P3_ADD_360_1242_U49, P3_ADD_360_1242_U50, P3_ADD_360_1242_U51, P3_ADD_360_1242_U52, P3_ADD_360_1242_U53, P3_ADD_360_1242_U54, P3_ADD_360_1242_U55, P3_ADD_360_1242_U56, P3_ADD_360_1242_U57, P3_ADD_360_1242_U58, P3_ADD_360_1242_U59, P3_ADD_360_1242_U60, P3_ADD_360_1242_U61, P3_ADD_360_1242_U62, P3_ADD_360_1242_U63, P3_ADD_360_1242_U64, P3_ADD_360_1242_U65, P3_ADD_360_1242_U66, P3_ADD_360_1242_U67, P3_ADD_360_1242_U68, P3_ADD_360_1242_U69, P3_ADD_360_1242_U70, P3_ADD_360_1242_U71, P3_ADD_360_1242_U72, P3_ADD_360_1242_U73, P3_ADD_360_1242_U74, P3_ADD_360_1242_U75, P3_ADD_360_1242_U76, P3_ADD_360_1242_U77, P3_ADD_360_1242_U78, P3_ADD_360_1242_U79, P3_ADD_360_1242_U80, P3_ADD_360_1242_U81, P3_ADD_360_1242_U82, P3_ADD_360_1242_U83, P3_ADD_360_1242_U84, P3_ADD_360_1242_U85, P3_ADD_360_1242_U86, P3_ADD_360_1242_U87, P3_ADD_360_1242_U88, P3_ADD_360_1242_U89, P3_ADD_360_1242_U90, P3_ADD_360_1242_U91, P3_ADD_360_1242_U92, P3_ADD_360_1242_U93, P3_ADD_360_1242_U94, P3_ADD_360_1242_U95, P3_ADD_360_1242_U96, P3_ADD_360_1242_U97, P3_ADD_360_1242_U98, P3_ADD_360_1242_U99, P3_ADD_360_1242_U100, P3_ADD_360_1242_U101, P3_ADD_360_1242_U102, P3_ADD_360_1242_U103, P3_ADD_360_1242_U104, P3_ADD_360_1242_U105, P3_ADD_360_1242_U106, P3_ADD_360_1242_U107, P3_ADD_360_1242_U108, P3_ADD_360_1242_U109, P3_ADD_360_1242_U110, P3_ADD_360_1242_U111, P3_ADD_360_1242_U112, P3_ADD_360_1242_U113, P3_ADD_360_1242_U114, P3_ADD_360_1242_U115, P3_ADD_360_1242_U116, P3_ADD_360_1242_U117, P3_ADD_360_1242_U118, P3_ADD_360_1242_U119, P3_ADD_360_1242_U120, P3_ADD_360_1242_U121, P3_ADD_360_1242_U122, P3_ADD_360_1242_U123, P3_ADD_360_1242_U124, P3_ADD_360_1242_U125, P3_ADD_360_1242_U126, P3_ADD_360_1242_U127, P3_ADD_360_1242_U128, P3_ADD_360_1242_U129, P3_ADD_360_1242_U130, P3_ADD_360_1242_U131, P3_ADD_360_1242_U132, P3_ADD_360_1242_U133, P3_ADD_360_1242_U134, P3_ADD_360_1242_U135, P3_ADD_360_1242_U136, P3_ADD_360_1242_U137, P3_ADD_360_1242_U138, P3_ADD_360_1242_U139, P3_ADD_360_1242_U140, P3_ADD_360_1242_U141, P3_ADD_360_1242_U142, P3_ADD_360_1242_U143, P3_ADD_360_1242_U144, P3_ADD_360_1242_U145, P3_ADD_360_1242_U146, P3_ADD_360_1242_U147, P3_ADD_360_1242_U148, P3_ADD_360_1242_U149, P3_ADD_360_1242_U150, P3_ADD_360_1242_U151, P3_ADD_360_1242_U152, P3_ADD_360_1242_U153, P3_ADD_360_1242_U154, P3_ADD_360_1242_U155, P3_ADD_360_1242_U156, P3_ADD_360_1242_U157, P3_ADD_360_1242_U158, P3_ADD_360_1242_U159, P3_ADD_360_1242_U160, P3_ADD_360_1242_U161, P3_ADD_360_1242_U162, P3_ADD_360_1242_U163, P3_ADD_360_1242_U164, P3_ADD_360_1242_U165, P3_ADD_360_1242_U166, P3_ADD_360_1242_U167, P3_ADD_360_1242_U168, P3_ADD_360_1242_U169, P3_ADD_360_1242_U170, P3_ADD_360_1242_U171, P3_ADD_360_1242_U172, P3_ADD_360_1242_U173, P3_ADD_360_1242_U174, P3_ADD_360_1242_U175, P3_ADD_360_1242_U176, P3_ADD_360_1242_U177, P3_ADD_360_1242_U178, P3_ADD_360_1242_U179, P3_ADD_360_1242_U180, P3_ADD_360_1242_U181, P3_ADD_360_1242_U182, P3_ADD_360_1242_U183, P3_ADD_360_1242_U184, P3_ADD_360_1242_U185, P3_ADD_360_1242_U186, P3_ADD_360_1242_U187, P3_ADD_360_1242_U188, P3_ADD_360_1242_U189, P3_ADD_360_1242_U190, P3_ADD_360_1242_U191, P3_ADD_360_1242_U192, P3_ADD_360_1242_U193, P3_ADD_360_1242_U194, P3_ADD_360_1242_U195, P3_ADD_360_1242_U196, P3_ADD_360_1242_U197, P3_ADD_360_1242_U198, P3_ADD_360_1242_U199, P3_ADD_360_1242_U200, P3_ADD_360_1242_U201, P3_ADD_360_1242_U202, P3_ADD_360_1242_U203, P3_ADD_360_1242_U204, P3_ADD_360_1242_U205, P3_ADD_360_1242_U206, P3_ADD_360_1242_U207, P3_ADD_360_1242_U208, P3_ADD_360_1242_U209, P3_ADD_360_1242_U210, P3_ADD_360_1242_U211, P3_ADD_360_1242_U212, P3_ADD_360_1242_U213, P3_ADD_360_1242_U214, P3_ADD_360_1242_U215, P3_ADD_360_1242_U216, P3_ADD_360_1242_U217, P3_ADD_360_1242_U218, P3_ADD_360_1242_U219, P3_ADD_360_1242_U220, P3_ADD_360_1242_U221, P3_ADD_360_1242_U222, P3_ADD_360_1242_U223, P3_ADD_360_1242_U224, P3_ADD_360_1242_U225, P3_ADD_360_1242_U226, P3_ADD_360_1242_U227, P3_ADD_360_1242_U228, P3_ADD_360_1242_U229, P3_ADD_360_1242_U230, P3_ADD_360_1242_U231, P3_ADD_360_1242_U232, P3_ADD_360_1242_U233, P3_ADD_360_1242_U234, P3_ADD_360_1242_U235, P3_ADD_360_1242_U236, P3_ADD_360_1242_U237, P3_ADD_360_1242_U238, P3_ADD_360_1242_U239, P3_ADD_360_1242_U240, P3_ADD_360_1242_U241, P3_ADD_360_1242_U242, P3_ADD_360_1242_U243, P3_ADD_360_1242_U244, P3_ADD_360_1242_U245, P3_ADD_360_1242_U246, P3_ADD_360_1242_U247, P3_ADD_360_1242_U248, P3_ADD_360_1242_U249, P3_ADD_360_1242_U250, P3_ADD_360_1242_U251, P3_ADD_360_1242_U252, P3_ADD_360_1242_U253, P3_ADD_360_1242_U254, P3_ADD_360_1242_U255, P3_ADD_360_1242_U256, P3_ADD_360_1242_U257, P3_ADD_360_1242_U258, P3_LT_563_1260_U6, P3_LT_563_1260_U7, P3_SUB_589_U6, P3_SUB_589_U7, P3_SUB_589_U8, P3_SUB_589_U9, P3_ADD_467_U4, P3_ADD_467_U5, P3_ADD_467_U6, P3_ADD_467_U7, P3_ADD_467_U8, P3_ADD_467_U9, P3_ADD_467_U10, P3_ADD_467_U11, P3_ADD_467_U12, P3_ADD_467_U13, P3_ADD_467_U14, P3_ADD_467_U15, P3_ADD_467_U16, P3_ADD_467_U17, P3_ADD_467_U18, P3_ADD_467_U19, P3_ADD_467_U20, P3_ADD_467_U21, P3_ADD_467_U22, P3_ADD_467_U23, P3_ADD_467_U24, P3_ADD_467_U25, P3_ADD_467_U26, P3_ADD_467_U27, P3_ADD_467_U28, P3_ADD_467_U29, P3_ADD_467_U30, P3_ADD_467_U31, P3_ADD_467_U32, P3_ADD_467_U33, P3_ADD_467_U34, P3_ADD_467_U35, P3_ADD_467_U36, P3_ADD_467_U37, P3_ADD_467_U38, P3_ADD_467_U39, P3_ADD_467_U40, P3_ADD_467_U41, P3_ADD_467_U42, P3_ADD_467_U43, P3_ADD_467_U44, P3_ADD_467_U45, P3_ADD_467_U46, P3_ADD_467_U47, P3_ADD_467_U48, P3_ADD_467_U49, P3_ADD_467_U50, P3_ADD_467_U51, P3_ADD_467_U52, P3_ADD_467_U53, P3_ADD_467_U54, P3_ADD_467_U55, P3_ADD_467_U56, P3_ADD_467_U57, P3_ADD_467_U58, P3_ADD_467_U59, P3_ADD_467_U60, P3_ADD_467_U61, P3_ADD_467_U62, P3_ADD_467_U63, P3_ADD_467_U64, P3_ADD_467_U65, P3_ADD_467_U66, P3_ADD_467_U67, P3_ADD_467_U68, P3_ADD_467_U69, P3_ADD_467_U70, P3_ADD_467_U71, P3_ADD_467_U72, P3_ADD_467_U73, P3_ADD_467_U74, P3_ADD_467_U75, P3_ADD_467_U76, P3_ADD_467_U77, P3_ADD_467_U78, P3_ADD_467_U79, P3_ADD_467_U80, P3_ADD_467_U81, P3_ADD_467_U82, P3_ADD_467_U83, P3_ADD_467_U84, P3_ADD_467_U85, P3_ADD_467_U86, P3_ADD_467_U87, P3_ADD_467_U88, P3_ADD_467_U89, P3_ADD_467_U90, P3_ADD_467_U91, P3_ADD_467_U92, P3_ADD_467_U93, P3_ADD_467_U94, P3_ADD_467_U95, P3_ADD_467_U96, P3_ADD_467_U97, P3_ADD_467_U98, P3_ADD_467_U99, P3_ADD_467_U100, P3_ADD_467_U101, P3_ADD_467_U102, P3_ADD_467_U103, P3_ADD_467_U104, P3_ADD_467_U105, P3_ADD_467_U106, P3_ADD_467_U107, P3_ADD_467_U108, P3_ADD_467_U109, P3_ADD_467_U110, P3_ADD_467_U111, P3_ADD_467_U112, P3_ADD_467_U113, P3_ADD_467_U114, P3_ADD_467_U115, P3_ADD_467_U116, P3_ADD_467_U117, P3_ADD_467_U118, P3_ADD_467_U119, P3_ADD_467_U120, P3_ADD_467_U121, P3_ADD_467_U122, P3_ADD_467_U123, P3_ADD_467_U124, P3_ADD_467_U125, P3_ADD_467_U126, P3_ADD_467_U127, P3_ADD_467_U128, P3_ADD_467_U129, P3_ADD_467_U130, P3_ADD_467_U131, P3_ADD_467_U132, P3_ADD_467_U133, P3_ADD_467_U134, P3_ADD_467_U135, P3_ADD_467_U136, P3_ADD_467_U137, P3_ADD_467_U138, P3_ADD_467_U139, P3_ADD_467_U140, P3_ADD_467_U141, P3_ADD_467_U142, P3_ADD_467_U143, P3_ADD_467_U144, P3_ADD_467_U145, P3_ADD_467_U146, P3_ADD_467_U147, P3_ADD_467_U148, P3_ADD_467_U149, P3_ADD_467_U150, P3_ADD_467_U151, P3_ADD_467_U152, P3_ADD_467_U153, P3_ADD_467_U154, P3_ADD_467_U155, P3_ADD_467_U156, P3_ADD_467_U157, P3_ADD_467_U158, P3_ADD_467_U159, P3_ADD_467_U160, P3_ADD_467_U161, P3_ADD_467_U162, P3_ADD_467_U163, P3_ADD_467_U164, P3_ADD_467_U165, P3_ADD_467_U166, P3_ADD_467_U167, P3_ADD_467_U168, P3_ADD_467_U169, P3_ADD_467_U170, P3_ADD_467_U171, P3_ADD_467_U172, P3_ADD_467_U173, P3_ADD_467_U174, P3_ADD_467_U175, P3_ADD_467_U176, P3_ADD_467_U177, P3_ADD_467_U178, P3_ADD_467_U179, P3_ADD_467_U180, P3_ADD_467_U181, P3_ADD_467_U182, P3_ADD_430_U4, P3_ADD_430_U5, P3_ADD_430_U6, P3_ADD_430_U7, P3_ADD_430_U8, P3_ADD_430_U9, P3_ADD_430_U10, P3_ADD_430_U11, P3_ADD_430_U12, P3_ADD_430_U13, P3_ADD_430_U14, P3_ADD_430_U15, P3_ADD_430_U16, P3_ADD_430_U17, P3_ADD_430_U18, P3_ADD_430_U19, P3_ADD_430_U20, P3_ADD_430_U21, P3_ADD_430_U22, P3_ADD_430_U23, P3_ADD_430_U24, P3_ADD_430_U25, P3_ADD_430_U26, P3_ADD_430_U27, P3_ADD_430_U28, P3_ADD_430_U29, P3_ADD_430_U30, P3_ADD_430_U31, P3_ADD_430_U32, P3_ADD_430_U33, P3_ADD_430_U34, P3_ADD_430_U35, P3_ADD_430_U36, P3_ADD_430_U37, P3_ADD_430_U38, P3_ADD_430_U39, P3_ADD_430_U40, P3_ADD_430_U41, P3_ADD_430_U42, P3_ADD_430_U43, P3_ADD_430_U44, P3_ADD_430_U45, P3_ADD_430_U46, P3_ADD_430_U47, P3_ADD_430_U48, P3_ADD_430_U49, P3_ADD_430_U50, P3_ADD_430_U51, P3_ADD_430_U52, P3_ADD_430_U53, P3_ADD_430_U54, P3_ADD_430_U55, P3_ADD_430_U56, P3_ADD_430_U57, P3_ADD_430_U58, P3_ADD_430_U59, P3_ADD_430_U60, P3_ADD_430_U61, P3_ADD_430_U62, P3_ADD_430_U63, P3_ADD_430_U64, P3_ADD_430_U65, P3_ADD_430_U66, P3_ADD_430_U67, P3_ADD_430_U68, P3_ADD_430_U69, P3_ADD_430_U70, P3_ADD_430_U71, P3_ADD_430_U72, P3_ADD_430_U73, P3_ADD_430_U74, P3_ADD_430_U75, P3_ADD_430_U76, P3_ADD_430_U77, P3_ADD_430_U78, P3_ADD_430_U79, P3_ADD_430_U80, P3_ADD_430_U81, P3_ADD_430_U82, P3_ADD_430_U83, P3_ADD_430_U84, P3_ADD_430_U85, P3_ADD_430_U86, P3_ADD_430_U87, P3_ADD_430_U88, P3_ADD_430_U89, P3_ADD_430_U90, P3_ADD_430_U91, P3_ADD_430_U92, P3_ADD_430_U93, P3_ADD_430_U94, P3_ADD_430_U95, P3_ADD_430_U96, P3_ADD_430_U97, P3_ADD_430_U98, P3_ADD_430_U99, P3_ADD_430_U100, P3_ADD_430_U101, P3_ADD_430_U102, P3_ADD_430_U103, P3_ADD_430_U104, P3_ADD_430_U105, P3_ADD_430_U106, P3_ADD_430_U107, P3_ADD_430_U108, P3_ADD_430_U109, P3_ADD_430_U110, P3_ADD_430_U111, P3_ADD_430_U112, P3_ADD_430_U113, P3_ADD_430_U114, P3_ADD_430_U115, P3_ADD_430_U116, P3_ADD_430_U117, P3_ADD_430_U118, P3_ADD_430_U119, P3_ADD_430_U120, P3_ADD_430_U121, P3_ADD_430_U122, P3_ADD_430_U123, P3_ADD_430_U124, P3_ADD_430_U125, P3_ADD_430_U126, P3_ADD_430_U127, P3_ADD_430_U128, P3_ADD_430_U129, P3_ADD_430_U130, P3_ADD_430_U131, P3_ADD_430_U132, P3_ADD_430_U133, P3_ADD_430_U134, P3_ADD_430_U135, P3_ADD_430_U136, P3_ADD_430_U137, P3_ADD_430_U138, P3_ADD_430_U139, P3_ADD_430_U140, P3_ADD_430_U141, P3_ADD_430_U142, P3_ADD_430_U143, P3_ADD_430_U144, P3_ADD_430_U145, P3_ADD_430_U146, P3_ADD_430_U147, P3_ADD_430_U148, P3_ADD_430_U149, P3_ADD_430_U150, P3_ADD_430_U151, P3_ADD_430_U152, P3_ADD_430_U153, P3_ADD_430_U154, P3_ADD_430_U155, P3_ADD_430_U156, P3_ADD_430_U157, P3_ADD_430_U158, P3_ADD_430_U159, P3_ADD_430_U160, P3_ADD_430_U161, P3_ADD_430_U162, P3_ADD_430_U163, P3_ADD_430_U164, P3_ADD_430_U165, P3_ADD_430_U166, P3_ADD_430_U167, P3_ADD_430_U168, P3_ADD_430_U169, P3_ADD_430_U170, P3_ADD_430_U171, P3_ADD_430_U172, P3_ADD_430_U173, P3_ADD_430_U174, P3_ADD_430_U175, P3_ADD_430_U176, P3_ADD_430_U177, P3_ADD_430_U178, P3_ADD_430_U179, P3_ADD_430_U180, P3_ADD_430_U181, P3_ADD_430_U182, P3_ADD_380_U5, P3_ADD_380_U6, P3_ADD_380_U7, P3_ADD_380_U8, P3_ADD_380_U9, P3_ADD_380_U10, P3_ADD_380_U11, P3_ADD_380_U12, P3_ADD_380_U13, P3_ADD_380_U14, P3_ADD_380_U15, P3_ADD_380_U16, P3_ADD_380_U17, P3_ADD_380_U18, P3_ADD_380_U19, P3_ADD_380_U20, P3_ADD_380_U21, P3_ADD_380_U22, P3_ADD_380_U23, P3_ADD_380_U24, P3_ADD_380_U25, P3_ADD_380_U26, P3_ADD_380_U27, P3_ADD_380_U28, P3_ADD_380_U29, P3_ADD_380_U30, P3_ADD_380_U31, P3_ADD_380_U32, P3_ADD_380_U33, P3_ADD_380_U34, P3_ADD_380_U35, P3_ADD_380_U36, P3_ADD_380_U37, P3_ADD_380_U38, P3_ADD_380_U39, P3_ADD_380_U40, P3_ADD_380_U41, P3_ADD_380_U42, P3_ADD_380_U43, P3_ADD_380_U44, P3_ADD_380_U45, P3_ADD_380_U46, P3_ADD_380_U47, P3_ADD_380_U48, P3_ADD_380_U49, P3_ADD_380_U50, P3_ADD_380_U51, P3_ADD_380_U52, P3_ADD_380_U53, P3_ADD_380_U54, P3_ADD_380_U55, P3_ADD_380_U56, P3_ADD_380_U57, P3_ADD_380_U58, P3_ADD_380_U59, P3_ADD_380_U60, P3_ADD_380_U61, P3_ADD_380_U62, P3_ADD_380_U63, P3_ADD_380_U64, P3_ADD_380_U65, P3_ADD_380_U66, P3_ADD_380_U67, P3_ADD_380_U68, P3_ADD_380_U69, P3_ADD_380_U70, P3_ADD_380_U71, P3_ADD_380_U72, P3_ADD_380_U73, P3_ADD_380_U74, P3_ADD_380_U75, P3_ADD_380_U76, P3_ADD_380_U77, P3_ADD_380_U78, P3_ADD_380_U79, P3_ADD_380_U80, P3_ADD_380_U81, P3_ADD_380_U82, P3_ADD_380_U83, P3_ADD_380_U84, P3_ADD_380_U85, P3_ADD_380_U86, P3_ADD_380_U87, P3_ADD_380_U88, P3_ADD_380_U89, P3_ADD_380_U90, P3_ADD_380_U91, P3_ADD_380_U92, P3_ADD_380_U93, P3_ADD_380_U94, P3_ADD_380_U95, P3_ADD_380_U96, P3_ADD_380_U97, P3_ADD_380_U98, P3_ADD_380_U99, P3_ADD_380_U100, P3_ADD_380_U101, P3_ADD_380_U102, P3_ADD_380_U103, P3_ADD_380_U104, P3_ADD_380_U105, P3_ADD_380_U106, P3_ADD_380_U107, P3_ADD_380_U108, P3_ADD_380_U109, P3_ADD_380_U110, P3_ADD_380_U111, P3_ADD_380_U112, P3_ADD_380_U113, P3_ADD_380_U114, P3_ADD_380_U115, P3_ADD_380_U116, P3_ADD_380_U117, P3_ADD_380_U118, P3_ADD_380_U119, P3_ADD_380_U120, P3_ADD_380_U121, P3_ADD_380_U122, P3_ADD_380_U123, P3_ADD_380_U124, P3_ADD_380_U125, P3_ADD_380_U126, P3_ADD_380_U127, P3_ADD_380_U128, P3_ADD_380_U129, P3_ADD_380_U130, P3_ADD_380_U131, P3_ADD_380_U132, P3_ADD_380_U133, P3_ADD_380_U134, P3_ADD_380_U135, P3_ADD_380_U136, P3_ADD_380_U137, P3_ADD_380_U138, P3_ADD_380_U139, P3_ADD_380_U140, P3_ADD_380_U141, P3_ADD_380_U142, P3_ADD_380_U143, P3_ADD_380_U144, P3_ADD_380_U145, P3_ADD_380_U146, P3_ADD_380_U147, P3_ADD_380_U148, P3_ADD_380_U149, P3_ADD_380_U150, P3_ADD_380_U151, P3_ADD_380_U152, P3_ADD_380_U153, P3_ADD_380_U154, P3_ADD_380_U155, P3_ADD_380_U156, P3_ADD_380_U157, P3_ADD_380_U158, P3_ADD_380_U159, P3_ADD_380_U160, P3_ADD_380_U161, P3_ADD_380_U162, P3_ADD_380_U163, P3_ADD_380_U164, P3_ADD_380_U165, P3_ADD_380_U166, P3_ADD_380_U167, P3_ADD_380_U168, P3_ADD_380_U169, P3_ADD_380_U170, P3_ADD_380_U171, P3_ADD_380_U172, P3_ADD_380_U173, P3_ADD_380_U174, P3_ADD_380_U175, P3_ADD_380_U176, P3_ADD_380_U177, P3_ADD_380_U178, P3_ADD_380_U179, P3_ADD_380_U180, P3_ADD_380_U181, P3_ADD_380_U182, P3_ADD_380_U183, P3_ADD_380_U184, P3_ADD_380_U185, P3_ADD_380_U186, P3_ADD_380_U187, P3_ADD_380_U188, P3_ADD_380_U189, P3_GTE_370_U6, P3_GTE_370_U7, P3_GTE_370_U8, P3_GTE_370_U9, P3_ADD_344_U5, P3_ADD_344_U6, P3_ADD_344_U7, P3_ADD_344_U8, P3_ADD_344_U9, P3_ADD_344_U10, P3_ADD_344_U11, P3_ADD_344_U12, P3_ADD_344_U13, P3_ADD_344_U14, P3_ADD_344_U15, P3_ADD_344_U16, P3_ADD_344_U17, P3_ADD_344_U18, P3_ADD_344_U19, P3_ADD_344_U20, P3_ADD_344_U21, P3_ADD_344_U22, P3_ADD_344_U23, P3_ADD_344_U24, P3_ADD_344_U25, P3_ADD_344_U26, P3_ADD_344_U27, P3_ADD_344_U28, P3_ADD_344_U29, P3_ADD_344_U30, P3_ADD_344_U31, P3_ADD_344_U32, P3_ADD_344_U33, P3_ADD_344_U34, P3_ADD_344_U35, P3_ADD_344_U36, P3_ADD_344_U37, P3_ADD_344_U38, P3_ADD_344_U39, P3_ADD_344_U40, P3_ADD_344_U41, P3_ADD_344_U42, P3_ADD_344_U43, P3_ADD_344_U44, P3_ADD_344_U45, P3_ADD_344_U46, P3_ADD_344_U47, P3_ADD_344_U48, P3_ADD_344_U49, P3_ADD_344_U50, P3_ADD_344_U51, P3_ADD_344_U52, P3_ADD_344_U53, P3_ADD_344_U54, P3_ADD_344_U55, P3_ADD_344_U56, P3_ADD_344_U57, P3_ADD_344_U58, P3_ADD_344_U59, P3_ADD_344_U60, P3_ADD_344_U61, P3_ADD_344_U62, P3_ADD_344_U63, P3_ADD_344_U64, P3_ADD_344_U65, P3_ADD_344_U66, P3_ADD_344_U67, P3_ADD_344_U68, P3_ADD_344_U69, P3_ADD_344_U70, P3_ADD_344_U71, P3_ADD_344_U72, P3_ADD_344_U73, P3_ADD_344_U74, P3_ADD_344_U75, P3_ADD_344_U76, P3_ADD_344_U77, P3_ADD_344_U78, P3_ADD_344_U79, P3_ADD_344_U80, P3_ADD_344_U81, P3_ADD_344_U82, P3_ADD_344_U83, P3_ADD_344_U84, P3_ADD_344_U85, P3_ADD_344_U86, P3_ADD_344_U87, P3_ADD_344_U88, P3_ADD_344_U89, P3_ADD_344_U90, P3_ADD_344_U91, P3_ADD_344_U92, P3_ADD_344_U93, P3_ADD_344_U94, P3_ADD_344_U95, P3_ADD_344_U96, P3_ADD_344_U97, P3_ADD_344_U98, P3_ADD_344_U99, P3_ADD_344_U100, P3_ADD_344_U101, P3_ADD_344_U102, P3_ADD_344_U103, P3_ADD_344_U104, P3_ADD_344_U105, P3_ADD_344_U106, P3_ADD_344_U107, P3_ADD_344_U108, P3_ADD_344_U109, P3_ADD_344_U110, P3_ADD_344_U111, P3_ADD_344_U112, P3_ADD_344_U113, P3_ADD_344_U114, P3_ADD_344_U115, P3_ADD_344_U116, P3_ADD_344_U117, P3_ADD_344_U118, P3_ADD_344_U119, P3_ADD_344_U120, P3_ADD_344_U121, P3_ADD_344_U122, P3_ADD_344_U123, P3_ADD_344_U124, P3_ADD_344_U125, P3_ADD_344_U126, P3_ADD_344_U127, P3_ADD_344_U128, P3_ADD_344_U129, P3_ADD_344_U130, P3_ADD_344_U131, P3_ADD_344_U132, P3_ADD_344_U133, P3_ADD_344_U134, P3_ADD_344_U135, P3_ADD_344_U136, P3_ADD_344_U137, P3_ADD_344_U138, P3_ADD_344_U139, P3_ADD_344_U140, P3_ADD_344_U141, P3_ADD_344_U142, P3_ADD_344_U143, P3_ADD_344_U144, P3_ADD_344_U145, P3_ADD_344_U146, P3_ADD_344_U147, P3_ADD_344_U148, P3_ADD_344_U149, P3_ADD_344_U150, P3_ADD_344_U151, P3_ADD_344_U152, P3_ADD_344_U153, P3_ADD_344_U154, P3_ADD_344_U155, P3_ADD_344_U156, P3_ADD_344_U157, P3_ADD_344_U158, P3_ADD_344_U159, P3_ADD_344_U160, P3_ADD_344_U161, P3_ADD_344_U162, P3_ADD_344_U163, P3_ADD_344_U164, P3_ADD_344_U165, P3_ADD_344_U166, P3_ADD_344_U167, P3_ADD_344_U168, P3_ADD_344_U169, P3_ADD_344_U170, P3_ADD_344_U171, P3_ADD_344_U172, P3_ADD_344_U173, P3_ADD_344_U174, P3_ADD_344_U175, P3_ADD_344_U176, P3_ADD_344_U177, P3_ADD_344_U178, P3_ADD_344_U179, P3_ADD_344_U180, P3_ADD_344_U181, P3_ADD_344_U182, P3_ADD_344_U183, P3_ADD_344_U184, P3_ADD_344_U185, P3_ADD_344_U186, P3_ADD_344_U187, P3_ADD_344_U188, P3_ADD_344_U189, P3_LT_563_U6, P3_LT_563_U7, P3_LT_563_U8, P3_LT_563_U9, P3_LT_563_U10, P3_LT_563_U11, P3_LT_563_U12, P3_LT_563_U13, P3_LT_563_U14, P3_LT_563_U15, P3_LT_563_U16, P3_LT_563_U17, P3_LT_563_U18, P3_LT_563_U19, P3_LT_563_U20, P3_LT_563_U21, P3_LT_563_U22, P3_LT_563_U23, P3_LT_563_U24, P3_LT_563_U25, P3_LT_563_U26, P3_LT_563_U27, P3_LT_563_U28, P3_ADD_339_U4, P3_ADD_339_U5, P3_ADD_339_U6, P3_ADD_339_U7, P3_ADD_339_U8, P3_ADD_339_U9, P3_ADD_339_U10, P3_ADD_339_U11, P3_ADD_339_U12, P3_ADD_339_U13, P3_ADD_339_U14, P3_ADD_339_U15, P3_ADD_339_U16, P3_ADD_339_U17, P3_ADD_339_U18, P3_ADD_339_U19, P3_ADD_339_U20, P3_ADD_339_U21, P3_ADD_339_U22, P3_ADD_339_U23, P3_ADD_339_U24, P3_ADD_339_U25, P3_ADD_339_U26, P3_ADD_339_U27, P3_ADD_339_U28, P3_ADD_339_U29, P3_ADD_339_U30, P3_ADD_339_U31, P3_ADD_339_U32, P3_ADD_339_U33, P3_ADD_339_U34, P3_ADD_339_U35, P3_ADD_339_U36, P3_ADD_339_U37, P3_ADD_339_U38, P3_ADD_339_U39, P3_ADD_339_U40, P3_ADD_339_U41, P3_ADD_339_U42, P3_ADD_339_U43, P3_ADD_339_U44, P3_ADD_339_U45, P3_ADD_339_U46, P3_ADD_339_U47, P3_ADD_339_U48, P3_ADD_339_U49, P3_ADD_339_U50, P3_ADD_339_U51, P3_ADD_339_U52, P3_ADD_339_U53, P3_ADD_339_U54, P3_ADD_339_U55, P3_ADD_339_U56, P3_ADD_339_U57, P3_ADD_339_U58, P3_ADD_339_U59, P3_ADD_339_U60, P3_ADD_339_U61, P3_ADD_339_U62, P3_ADD_339_U63, P3_ADD_339_U64, P3_ADD_339_U65, P3_ADD_339_U66, P3_ADD_339_U67, P3_ADD_339_U68, P3_ADD_339_U69, P3_ADD_339_U70, P3_ADD_339_U71, P3_ADD_339_U72, P3_ADD_339_U73, P3_ADD_339_U74, P3_ADD_339_U75, P3_ADD_339_U76, P3_ADD_339_U77, P3_ADD_339_U78, P3_ADD_339_U79, P3_ADD_339_U80, P3_ADD_339_U81, P3_ADD_339_U82, P3_ADD_339_U83, P3_ADD_339_U84, P3_ADD_339_U85, P3_ADD_339_U86, P3_ADD_339_U87, P3_ADD_339_U88, P3_ADD_339_U89, P3_ADD_339_U90, P3_ADD_339_U91, P3_ADD_339_U92, P3_ADD_339_U93, P3_ADD_339_U94, P3_ADD_339_U95, P3_ADD_339_U96, P3_ADD_339_U97, P3_ADD_339_U98, P3_ADD_339_U99, P3_ADD_339_U100, P3_ADD_339_U101, P3_ADD_339_U102, P3_ADD_339_U103, P3_ADD_339_U104, P3_ADD_339_U105, P3_ADD_339_U106, P3_ADD_339_U107, P3_ADD_339_U108, P3_ADD_339_U109, P3_ADD_339_U110, P3_ADD_339_U111, P3_ADD_339_U112, P3_ADD_339_U113, P3_ADD_339_U114, P3_ADD_339_U115, P3_ADD_339_U116, P3_ADD_339_U117, P3_ADD_339_U118, P3_ADD_339_U119, P3_ADD_339_U120, P3_ADD_339_U121, P3_ADD_339_U122, P3_ADD_339_U123, P3_ADD_339_U124, P3_ADD_339_U125, P3_ADD_339_U126, P3_ADD_339_U127, P3_ADD_339_U128, P3_ADD_339_U129, P3_ADD_339_U130, P3_ADD_339_U131, P3_ADD_339_U132, P3_ADD_339_U133, P3_ADD_339_U134, P3_ADD_339_U135, P3_ADD_339_U136, P3_ADD_339_U137, P3_ADD_339_U138, P3_ADD_339_U139, P3_ADD_339_U140, P3_ADD_339_U141, P3_ADD_339_U142, P3_ADD_339_U143, P3_ADD_339_U144, P3_ADD_339_U145, P3_ADD_339_U146, P3_ADD_339_U147, P3_ADD_339_U148, P3_ADD_339_U149, P3_ADD_339_U150, P3_ADD_339_U151, P3_ADD_339_U152, P3_ADD_339_U153, P3_ADD_339_U154, P3_ADD_339_U155, P3_ADD_339_U156, P3_ADD_339_U157, P3_ADD_339_U158, P3_ADD_339_U159, P3_ADD_339_U160, P3_ADD_339_U161, P3_ADD_339_U162, P3_ADD_339_U163, P3_ADD_339_U164, P3_ADD_339_U165, P3_ADD_339_U166, P3_ADD_339_U167, P3_ADD_339_U168, P3_ADD_339_U169, P3_ADD_339_U170, P3_ADD_339_U171, P3_ADD_339_U172, P3_ADD_339_U173, P3_ADD_339_U174, P3_ADD_339_U175, P3_ADD_339_U176, P3_ADD_339_U177, P3_ADD_339_U178, P3_ADD_339_U179, P3_ADD_339_U180, P3_ADD_339_U181, P3_ADD_339_U182, P3_ADD_360_U4, P3_ADD_360_U5, P3_ADD_360_U6, P3_ADD_360_U7, P3_ADD_360_U8, P3_ADD_360_U9, P3_ADD_360_U10, P3_ADD_360_U11, P3_ADD_360_U12, P3_ADD_360_U13, P3_ADD_360_U14, P3_ADD_360_U15, P3_ADD_360_U16, P3_ADD_360_U17, P3_ADD_360_U18, P3_ADD_360_U19, P3_ADD_360_U20, P3_ADD_360_U21, P3_ADD_360_U22, P3_ADD_360_U23, P3_ADD_360_U24, P3_ADD_360_U25, P3_ADD_360_U26, P3_ADD_360_U27, P3_ADD_360_U28, P3_ADD_360_U29, P3_ADD_360_U30, P3_ADD_360_U31, P3_ADD_360_U32, P3_ADD_360_U33, P3_ADD_360_U34, P3_ADD_360_U35, P3_ADD_360_U36, P3_ADD_360_U37, P3_ADD_360_U38, P3_ADD_360_U39, P3_ADD_360_U40, P3_LTE_597_U6, P3_SUB_580_U6, P3_SUB_580_U7, P3_SUB_580_U8, P3_SUB_580_U9, P3_SUB_580_U10, P3_LT_589_U6, P3_LT_589_U7, P3_LT_589_U8, P3_ADD_541_U4, P3_ADD_541_U5, P3_ADD_541_U6, P3_ADD_541_U7, P3_ADD_541_U8, P3_ADD_541_U9, P3_ADD_541_U10, P3_ADD_541_U11, P3_ADD_541_U12, P3_ADD_541_U13, P3_ADD_541_U14, P3_ADD_541_U15, P3_ADD_541_U16, P3_ADD_541_U17, P3_ADD_541_U18, P3_ADD_541_U19, P3_ADD_541_U20, P3_ADD_541_U21, P3_ADD_541_U22, P3_ADD_541_U23, P3_ADD_541_U24, P3_ADD_541_U25, P3_ADD_541_U26, P3_ADD_541_U27, P3_ADD_541_U28, P3_ADD_541_U29, P3_ADD_541_U30, P3_ADD_541_U31, P3_ADD_541_U32, P3_ADD_541_U33, P3_ADD_541_U34, P3_ADD_541_U35, P3_ADD_541_U36, P3_ADD_541_U37, P3_ADD_541_U38, P3_ADD_541_U39, P3_ADD_541_U40, P3_ADD_541_U41, P3_ADD_541_U42, P3_ADD_541_U43, P3_ADD_541_U44, P3_ADD_541_U45, P3_ADD_541_U46, P3_ADD_541_U47, P3_ADD_541_U48, P3_ADD_541_U49, P3_ADD_541_U50, P3_ADD_541_U51, P3_ADD_541_U52, P3_ADD_541_U53, P3_ADD_541_U54, P3_ADD_541_U55, P3_ADD_541_U56, P3_ADD_541_U57, P3_ADD_541_U58, P3_ADD_541_U59, P3_ADD_541_U60, P3_ADD_541_U61, P3_ADD_541_U62, P3_ADD_541_U63, P3_ADD_541_U64, P3_ADD_541_U65, P3_ADD_541_U66, P3_ADD_541_U67, P3_ADD_541_U68, P3_ADD_541_U69, P3_ADD_541_U70, P3_ADD_541_U71, P3_ADD_541_U72, P3_ADD_541_U73, P3_ADD_541_U74, P3_ADD_541_U75, P3_ADD_541_U76, P3_ADD_541_U77, P3_ADD_541_U78, P3_ADD_541_U79, P3_ADD_541_U80, P3_ADD_541_U81, P3_ADD_541_U82, P3_ADD_541_U83, P3_ADD_541_U84, P3_ADD_541_U85, P3_ADD_541_U86, P3_ADD_541_U87, P3_ADD_541_U88, P3_ADD_541_U89, P3_ADD_541_U90, P3_ADD_541_U91, P3_ADD_541_U92, P3_ADD_541_U93, P3_ADD_541_U94, P3_ADD_541_U95, P3_ADD_541_U96, P3_ADD_541_U97, P3_ADD_541_U98, P3_ADD_541_U99, P3_ADD_541_U100, P3_ADD_541_U101, P3_ADD_541_U102, P3_ADD_541_U103, P3_ADD_541_U104, P3_ADD_541_U105, P3_ADD_541_U106, P3_ADD_541_U107, P3_ADD_541_U108, P3_ADD_541_U109, P3_ADD_541_U110, P3_ADD_541_U111, P3_ADD_541_U112, P3_ADD_541_U113, P3_ADD_541_U114, P3_ADD_541_U115, P3_ADD_541_U116, P3_ADD_541_U117, P3_ADD_541_U118, P3_ADD_541_U119, P3_ADD_541_U120, P3_ADD_541_U121, P3_ADD_541_U122, P3_ADD_541_U123, P3_ADD_541_U124, P3_ADD_541_U125, P3_ADD_541_U126, P3_ADD_541_U127, P3_ADD_541_U128, P3_ADD_541_U129, P3_ADD_541_U130, P3_ADD_541_U131, P3_ADD_541_U132, P3_ADD_541_U133, P3_ADD_541_U134, P3_ADD_541_U135, P3_ADD_541_U136, P3_ADD_541_U137, P3_ADD_541_U138, P3_ADD_541_U139, P3_ADD_541_U140, P3_ADD_541_U141, P3_ADD_541_U142, P3_ADD_541_U143, P3_ADD_541_U144, P3_ADD_541_U145, P3_ADD_541_U146, P3_ADD_541_U147, P3_ADD_541_U148, P3_ADD_541_U149, P3_ADD_541_U150, P3_ADD_541_U151, P3_ADD_541_U152, P3_ADD_541_U153, P3_ADD_541_U154, P3_ADD_541_U155, P3_ADD_541_U156, P3_ADD_541_U157, P3_ADD_541_U158, P3_ADD_541_U159, P3_ADD_541_U160, P3_ADD_541_U161, P3_ADD_541_U162, P3_ADD_541_U163, P3_ADD_541_U164, P3_ADD_541_U165, P3_ADD_541_U166, P3_ADD_541_U167, P3_ADD_541_U168, P3_ADD_541_U169, P3_ADD_541_U170, P3_ADD_541_U171, P3_ADD_541_U172, P3_ADD_541_U173, P3_ADD_541_U174, P3_ADD_541_U175, P3_ADD_541_U176, P3_ADD_541_U177, P3_ADD_541_U178, P3_ADD_541_U179, P3_ADD_541_U180, P3_ADD_541_U181, P3_ADD_541_U182, P3_SUB_355_U6, P3_SUB_355_U7, P3_SUB_355_U8, P3_SUB_355_U9, P3_SUB_355_U10, P3_SUB_355_U11, P3_SUB_355_U12, P3_SUB_355_U13, P3_SUB_355_U14, P3_SUB_355_U15, P3_SUB_355_U16, P3_SUB_355_U17, P3_SUB_355_U18, P3_SUB_355_U19, P3_SUB_355_U20, P3_SUB_355_U21, P3_SUB_355_U22, P3_SUB_355_U23, P3_SUB_355_U24, P3_SUB_355_U25, P3_SUB_355_U26, P3_SUB_355_U27, P3_SUB_355_U28, P3_SUB_355_U29, P3_SUB_355_U30, P3_SUB_355_U31, P3_SUB_355_U32, P3_SUB_355_U33, P3_SUB_355_U34, P3_SUB_355_U35, P3_SUB_355_U36, P3_SUB_355_U37, P3_SUB_355_U38, P3_SUB_355_U39, P3_SUB_355_U40, P3_SUB_355_U41, P3_SUB_355_U42, P3_SUB_355_U43, P3_SUB_355_U44, P3_SUB_355_U45, P3_SUB_355_U46, P3_SUB_355_U47, P3_SUB_355_U48, P3_SUB_355_U49, P3_SUB_355_U50, P3_SUB_355_U51, P3_SUB_355_U52, P3_SUB_355_U53, P3_SUB_355_U54, P3_SUB_355_U55, P3_SUB_355_U56, P3_SUB_355_U57, P3_SUB_355_U58, P3_SUB_355_U59, P3_SUB_355_U60, P3_SUB_355_U61, P3_SUB_355_U62, P3_SUB_355_U63, P3_SUB_355_U64, P3_SUB_355_U65, P3_SUB_355_U66, P3_SUB_450_U6, P3_SUB_450_U7, P3_SUB_450_U8, P3_SUB_450_U9, P3_SUB_450_U10, P3_SUB_450_U11, P3_SUB_450_U12, P3_SUB_450_U13, P3_SUB_450_U14, P3_SUB_450_U15, P3_SUB_450_U16, P3_SUB_450_U17, P3_SUB_450_U18, P3_SUB_450_U19, P3_SUB_450_U20, P3_SUB_450_U21, P3_SUB_450_U22, P3_SUB_450_U23, P3_SUB_450_U24, P3_SUB_450_U25, P3_SUB_450_U26, P3_SUB_450_U27, P3_SUB_450_U28, P3_SUB_450_U29, P3_SUB_450_U30, P3_SUB_450_U31, P3_SUB_450_U32, P3_SUB_450_U33, P3_SUB_450_U34, P3_SUB_450_U35, P3_SUB_450_U36, P3_SUB_450_U37, P3_SUB_450_U38, P3_SUB_450_U39, P3_SUB_450_U40, P3_SUB_450_U41, P3_SUB_450_U42, P3_SUB_450_U43, P3_SUB_450_U44, P3_SUB_450_U45, P3_SUB_450_U46, P3_SUB_450_U47, P3_SUB_450_U48, P3_SUB_450_U49, P3_SUB_450_U50, P3_SUB_450_U51, P3_SUB_450_U52, P3_SUB_450_U53, P3_SUB_450_U54, P3_SUB_450_U55, P3_SUB_450_U56, P3_SUB_450_U57, P3_SUB_450_U58, P3_SUB_450_U59, P3_SUB_450_U60, P3_SUB_450_U61, P3_SUB_450_U62, P3_SUB_450_U63, P3_SUB_357_1258_U4, P3_SUB_357_1258_U5, P3_SUB_357_1258_U6, P3_SUB_357_1258_U7, P3_SUB_357_1258_U8, P3_SUB_357_1258_U9, P3_SUB_357_1258_U10, P3_SUB_357_1258_U11, P3_SUB_357_1258_U12, P3_SUB_357_1258_U13, P3_SUB_357_1258_U14, P3_SUB_357_1258_U15, P3_SUB_357_1258_U16, P3_SUB_357_1258_U17, P3_SUB_357_1258_U18, P3_SUB_357_1258_U19, P3_SUB_357_1258_U20, P3_SUB_357_1258_U21, P3_SUB_357_1258_U22, P3_SUB_357_1258_U23, P3_SUB_357_1258_U24, P3_SUB_357_1258_U25, P3_SUB_357_1258_U26, P3_SUB_357_1258_U27, P3_SUB_357_1258_U28, P3_SUB_357_1258_U29, P3_SUB_357_1258_U30, P3_SUB_357_1258_U31, P3_SUB_357_1258_U32, P3_SUB_357_1258_U33, P3_SUB_357_1258_U34, P3_SUB_357_1258_U35, P3_SUB_357_1258_U36, P3_SUB_357_1258_U37, P3_SUB_357_1258_U38, P3_SUB_357_1258_U39, P3_SUB_357_1258_U40, P3_SUB_357_1258_U41, P3_SUB_357_1258_U42, P3_SUB_357_1258_U43, P3_SUB_357_1258_U44, P3_SUB_357_1258_U45, P3_SUB_357_1258_U46, P3_SUB_357_1258_U47, P3_SUB_357_1258_U48, P3_SUB_357_1258_U49, P3_SUB_357_1258_U50, P3_SUB_357_1258_U51, P3_SUB_357_1258_U52, P3_SUB_357_1258_U53, P3_SUB_357_1258_U54, P3_SUB_357_1258_U55, P3_SUB_357_1258_U56, P3_SUB_357_1258_U57, P3_SUB_357_1258_U58, P3_SUB_357_1258_U59, P3_SUB_357_1258_U60, P3_SUB_357_1258_U61, P3_SUB_357_1258_U62, P3_SUB_357_1258_U63, P3_SUB_357_1258_U64, P3_SUB_357_1258_U65, P3_SUB_357_1258_U66, P3_SUB_357_1258_U67, P3_SUB_357_1258_U68, P3_SUB_357_1258_U69, P3_SUB_357_1258_U70, P3_SUB_357_1258_U71, P3_SUB_357_1258_U72, P3_SUB_357_1258_U73, P3_SUB_357_1258_U74, P3_SUB_357_1258_U75, P3_SUB_357_1258_U76, P3_SUB_357_1258_U77, P3_SUB_357_1258_U78, P3_SUB_357_1258_U79, P3_SUB_357_1258_U80, P3_SUB_357_1258_U81, P3_SUB_357_1258_U82, P3_SUB_357_1258_U83, P3_SUB_357_1258_U84, P3_SUB_357_1258_U85, P3_SUB_357_1258_U86, P3_SUB_357_1258_U87, P3_SUB_357_1258_U88, P3_SUB_357_1258_U89, P3_SUB_357_1258_U90, P3_SUB_357_1258_U91, P3_SUB_357_1258_U92, P3_SUB_357_1258_U93, P3_SUB_357_1258_U94, P3_SUB_357_1258_U95, P3_SUB_357_1258_U96, P3_SUB_357_1258_U97, P3_SUB_357_1258_U98, P3_SUB_357_1258_U99, P3_SUB_357_1258_U100, P3_SUB_357_1258_U101, P3_SUB_357_1258_U102, P3_SUB_357_1258_U103, P3_SUB_357_1258_U104, P3_SUB_357_1258_U105, P3_SUB_357_1258_U106, P3_SUB_357_1258_U107, P3_SUB_357_1258_U108, P3_SUB_357_1258_U109, P3_SUB_357_1258_U110, P3_SUB_357_1258_U111, P3_SUB_357_1258_U112, P3_SUB_357_1258_U113, P3_SUB_357_1258_U114, P3_SUB_357_1258_U115, P3_SUB_357_1258_U116, P3_SUB_357_1258_U117, P3_SUB_357_1258_U118, P3_SUB_357_1258_U119, P3_SUB_357_1258_U120, P3_SUB_357_1258_U121, P3_SUB_357_1258_U122, P3_SUB_357_1258_U123, P3_SUB_357_1258_U124, P3_SUB_357_1258_U125, P3_SUB_357_1258_U126, P3_SUB_357_1258_U127, P3_SUB_357_1258_U128, P3_SUB_357_1258_U129, P3_SUB_357_1258_U130, P3_SUB_357_1258_U131, P3_SUB_357_1258_U132, P3_SUB_357_1258_U133, P3_SUB_357_1258_U134, P3_SUB_357_1258_U135, P3_SUB_357_1258_U136, P3_SUB_357_1258_U137, P3_SUB_357_1258_U138, P3_SUB_357_1258_U139, P3_SUB_357_1258_U140, P3_SUB_357_1258_U141, P3_SUB_357_1258_U142, P3_SUB_357_1258_U143, P3_SUB_357_1258_U144, P3_SUB_357_1258_U145, P3_SUB_357_1258_U146, P3_SUB_357_1258_U147, P3_SUB_357_1258_U148, P3_SUB_357_1258_U149, P3_SUB_357_1258_U150, P3_SUB_357_1258_U151, P3_SUB_357_1258_U152, P3_SUB_357_1258_U153, P3_SUB_357_1258_U154, P3_SUB_357_1258_U155, P3_SUB_357_1258_U156, P3_SUB_357_1258_U157, P3_SUB_357_1258_U158, P3_SUB_357_1258_U159, P3_SUB_357_1258_U160, P3_SUB_357_1258_U161, P3_SUB_357_1258_U162, P3_SUB_357_1258_U163, P3_SUB_357_1258_U164, P3_SUB_357_1258_U165, P3_SUB_357_1258_U166, P3_SUB_357_1258_U167, P3_SUB_357_1258_U168, P3_SUB_357_1258_U169, P3_SUB_357_1258_U170, P3_SUB_357_1258_U171, P3_SUB_357_1258_U172, P3_SUB_357_1258_U173, P3_SUB_357_1258_U174, P3_SUB_357_1258_U175, P3_SUB_357_1258_U176, P3_SUB_357_1258_U177, P3_SUB_357_1258_U178, P3_SUB_357_1258_U179, P3_SUB_357_1258_U180, P3_SUB_357_1258_U181, P3_SUB_357_1258_U182, P3_SUB_357_1258_U183, P3_SUB_357_1258_U184, P3_SUB_357_1258_U185, P3_SUB_357_1258_U186, P3_SUB_357_1258_U187, P3_SUB_357_1258_U188, P3_SUB_357_1258_U189, P3_SUB_357_1258_U190, P3_SUB_357_1258_U191, P3_SUB_357_1258_U192, P3_SUB_357_1258_U193, P3_SUB_357_1258_U194, P3_SUB_357_1258_U195, P3_SUB_357_1258_U196, P3_SUB_357_1258_U197, P3_SUB_357_1258_U198, P3_SUB_357_1258_U199, P3_SUB_357_1258_U200, P3_SUB_357_1258_U201, P3_SUB_357_1258_U202, P3_SUB_357_1258_U203, P3_SUB_357_1258_U204, P3_SUB_357_1258_U205, P3_SUB_357_1258_U206, P3_SUB_357_1258_U207, P3_SUB_357_1258_U208, P3_SUB_357_1258_U209, P3_SUB_357_1258_U210, P3_SUB_357_1258_U211, P3_SUB_357_1258_U212, P3_SUB_357_1258_U213, P3_SUB_357_1258_U214, P3_SUB_357_1258_U215, P3_SUB_357_1258_U216, P3_SUB_357_1258_U217, P3_SUB_357_1258_U218, P3_SUB_357_1258_U219, P3_SUB_357_1258_U220, P3_SUB_357_1258_U221, P3_SUB_357_1258_U222, P3_SUB_357_1258_U223, P3_SUB_357_1258_U224, P3_SUB_357_1258_U225, P3_SUB_357_1258_U226, P3_SUB_357_1258_U227, P3_SUB_357_1258_U228, P3_SUB_357_1258_U229, P3_SUB_357_1258_U230, P3_SUB_357_1258_U231, P3_SUB_357_1258_U232, P3_SUB_357_1258_U233, P3_SUB_357_1258_U234, P3_SUB_357_1258_U235, P3_SUB_357_1258_U236, P3_SUB_357_1258_U237, P3_SUB_357_1258_U238, P3_SUB_357_1258_U239, P3_SUB_357_1258_U240, P3_SUB_357_1258_U241, P3_SUB_357_1258_U242, P3_SUB_357_1258_U243, P3_SUB_357_1258_U244, P3_SUB_357_1258_U245, P3_SUB_357_1258_U246, P3_SUB_357_1258_U247, P3_SUB_357_1258_U248, P3_SUB_357_1258_U249, P3_SUB_357_1258_U250, P3_SUB_357_1258_U251, P3_SUB_357_1258_U252, P3_SUB_357_1258_U253, P3_SUB_357_1258_U254, P3_SUB_357_1258_U255, P3_SUB_357_1258_U256, P3_SUB_357_1258_U257, P3_SUB_357_1258_U258, P3_SUB_357_1258_U259, P3_SUB_357_1258_U260, P3_SUB_357_1258_U261, P3_SUB_357_1258_U262, P3_SUB_357_1258_U263, P3_SUB_357_1258_U264, P3_SUB_357_1258_U265, P3_SUB_357_1258_U266, P3_SUB_357_1258_U267, P3_SUB_357_1258_U268, P3_SUB_357_1258_U269, P3_SUB_357_1258_U270, P3_SUB_357_1258_U271, P3_SUB_357_1258_U272, P3_SUB_357_1258_U273, P3_SUB_357_1258_U274, P3_SUB_357_1258_U275, P3_SUB_357_1258_U276, P3_SUB_357_1258_U277, P3_SUB_357_1258_U278, P3_SUB_357_1258_U279, P3_SUB_357_1258_U280, P3_SUB_357_1258_U281, P3_SUB_357_1258_U282, P3_SUB_357_1258_U283, P3_SUB_357_1258_U284, P3_SUB_357_1258_U285, P3_SUB_357_1258_U286, P3_SUB_357_1258_U287, P3_SUB_357_1258_U288, P3_SUB_357_1258_U289, P3_SUB_357_1258_U290, P3_SUB_357_1258_U291, P3_SUB_357_1258_U292, P3_SUB_357_1258_U293, P3_SUB_357_1258_U294, P3_SUB_357_1258_U295, P3_SUB_357_1258_U296, P3_SUB_357_1258_U297, P3_SUB_357_1258_U298, P3_SUB_357_1258_U299, P3_SUB_357_1258_U300, P3_SUB_357_1258_U301, P3_SUB_357_1258_U302, P3_SUB_357_1258_U303, P3_SUB_357_1258_U304, P3_SUB_357_1258_U305, P3_SUB_357_1258_U306, P3_SUB_357_1258_U307, P3_SUB_357_1258_U308, P3_SUB_357_1258_U309, P3_SUB_357_1258_U310, P3_SUB_357_1258_U311, P3_SUB_357_1258_U312, P3_SUB_357_1258_U313, P3_SUB_357_1258_U314, P3_SUB_357_1258_U315, P3_SUB_357_1258_U316, P3_SUB_357_1258_U317, P3_SUB_357_1258_U318, P3_SUB_357_1258_U319, P3_SUB_357_1258_U320, P3_SUB_357_1258_U321, P3_SUB_357_1258_U322, P3_SUB_357_1258_U323, P3_SUB_357_1258_U324, P3_SUB_357_1258_U325, P3_SUB_357_1258_U326, P3_SUB_357_1258_U327, P3_SUB_357_1258_U328, P3_SUB_357_1258_U329, P3_SUB_357_1258_U330, P3_SUB_357_1258_U331, P3_SUB_357_1258_U332, P3_SUB_357_1258_U333, P3_SUB_357_1258_U334, P3_SUB_357_1258_U335, P3_SUB_357_1258_U336, P3_SUB_357_1258_U337, P3_SUB_357_1258_U338, P3_SUB_357_1258_U339, P3_SUB_357_1258_U340, P3_SUB_357_1258_U341, P3_SUB_357_1258_U342, P3_SUB_357_1258_U343, P3_SUB_357_1258_U344, P3_SUB_357_1258_U345, P3_SUB_357_1258_U346, P3_SUB_357_1258_U347, P3_SUB_357_1258_U348, P3_SUB_357_1258_U349, P3_SUB_357_1258_U350, P3_SUB_357_1258_U351, P3_SUB_357_1258_U352, P3_SUB_357_1258_U353, P3_SUB_357_1258_U354, P3_SUB_357_1258_U355, P3_SUB_357_1258_U356, P3_SUB_357_1258_U357, P3_SUB_357_1258_U358, P3_SUB_357_1258_U359, P3_SUB_357_1258_U360, P3_SUB_357_1258_U361, P3_SUB_357_1258_U362, P3_SUB_357_1258_U363, P3_SUB_357_1258_U364, P3_SUB_357_1258_U365, P3_SUB_357_1258_U366, P3_SUB_357_1258_U367, P3_SUB_357_1258_U368, P3_SUB_357_1258_U369, P3_SUB_357_1258_U370, P3_SUB_357_1258_U371, P3_SUB_357_1258_U372, P3_SUB_357_1258_U373, P3_SUB_357_1258_U374, P3_SUB_357_1258_U375, P3_SUB_357_1258_U376, P3_SUB_357_1258_U377, P3_SUB_357_1258_U378, P3_SUB_357_1258_U379, P3_SUB_357_1258_U380, P3_SUB_357_1258_U381, P3_SUB_357_1258_U382, P3_SUB_357_1258_U383, P3_SUB_357_1258_U384, P3_SUB_357_1258_U385, P3_SUB_357_1258_U386, P3_SUB_357_1258_U387, P3_SUB_357_1258_U388, P3_SUB_357_1258_U389, P3_SUB_357_1258_U390, P3_SUB_357_1258_U391, P3_SUB_357_1258_U392, P3_SUB_357_1258_U393, P3_SUB_357_1258_U394, P3_SUB_357_1258_U395, P3_SUB_357_1258_U396, P3_SUB_357_1258_U397, P3_SUB_357_1258_U398, P3_SUB_357_1258_U399, P3_SUB_357_1258_U400, P3_SUB_357_1258_U401, P3_SUB_357_1258_U402, P3_SUB_357_1258_U403, P3_SUB_357_1258_U404, P3_SUB_357_1258_U405, P3_SUB_357_1258_U406, P3_SUB_357_1258_U407, P3_SUB_357_1258_U408, P3_SUB_357_1258_U409, P3_SUB_357_1258_U410, P3_SUB_357_1258_U411, P3_SUB_357_1258_U412, P3_SUB_357_1258_U413, P3_SUB_357_1258_U414, P3_SUB_357_1258_U415, P3_SUB_357_1258_U416, P3_SUB_357_1258_U417, P3_SUB_357_1258_U418, P3_SUB_357_1258_U419, P3_SUB_357_1258_U420, P3_SUB_357_1258_U421, P3_SUB_357_1258_U422, P3_SUB_357_1258_U423, P3_SUB_357_1258_U424, P3_SUB_357_1258_U425, P3_SUB_357_1258_U426, P3_SUB_357_1258_U427, P3_SUB_357_1258_U428, P3_SUB_357_1258_U429, P3_SUB_357_1258_U430, P3_SUB_357_1258_U431, P3_SUB_357_1258_U432, P3_SUB_357_1258_U433, P3_SUB_357_1258_U434, P3_SUB_357_1258_U435, P3_SUB_357_1258_U436, P3_SUB_357_1258_U437, P3_SUB_357_1258_U438, P3_SUB_357_1258_U439, P3_SUB_357_1258_U440, P3_SUB_357_1258_U441, P3_SUB_357_1258_U442, P3_SUB_357_1258_U443, P3_SUB_357_1258_U444, P3_SUB_357_1258_U445, P3_SUB_357_1258_U446, P3_SUB_357_1258_U447, P3_SUB_357_1258_U448, P3_SUB_357_1258_U449, P3_SUB_357_1258_U450, P3_SUB_357_1258_U451, P3_SUB_357_1258_U452, P3_SUB_357_1258_U453, P3_SUB_357_1258_U454, P3_SUB_357_1258_U455, P3_SUB_357_1258_U456, P3_SUB_357_1258_U457, P3_SUB_357_1258_U458, P3_SUB_357_1258_U459, P3_SUB_357_1258_U460, P3_SUB_357_1258_U461, P3_SUB_357_1258_U462, P3_SUB_357_1258_U463, P3_SUB_357_1258_U464, P3_SUB_357_1258_U465, P3_SUB_357_1258_U466, P3_SUB_357_1258_U467, P3_SUB_357_1258_U468, P3_SUB_357_1258_U469, P3_SUB_357_1258_U470, P3_SUB_357_1258_U471, P3_SUB_357_1258_U472, P3_SUB_357_1258_U473, P3_SUB_357_1258_U474, P3_SUB_357_1258_U475, P3_SUB_357_1258_U476, P3_SUB_357_1258_U477, P3_SUB_357_1258_U478, P3_SUB_357_1258_U479, P3_SUB_357_1258_U480, P3_SUB_357_1258_U481, P3_SUB_357_1258_U482, P3_SUB_357_1258_U483, P3_SUB_357_1258_U484, P3_ADD_486_U5, P3_ADD_486_U6, P3_ADD_486_U7, P3_ADD_486_U8, P3_ADD_486_U9, P3_ADD_486_U10, P3_ADD_486_U11, P3_ADD_486_U12, P3_ADD_486_U13, P3_ADD_486_U14, P3_ADD_486_U15, P3_ADD_486_U16, P3_ADD_486_U17, P3_ADD_486_U18, P3_ADD_486_U19, P3_ADD_486_U20, P3_ADD_486_U21, P3_ADD_486_U22, P3_ADD_486_U23, P3_ADD_486_U24, P3_ADD_486_U25, P3_ADD_486_U26, P3_ADD_486_U27, P3_ADD_486_U28, P3_SUB_485_U6, P3_SUB_485_U7, P3_SUB_485_U8, P3_SUB_485_U9, P3_SUB_485_U10, P3_SUB_485_U11, P3_SUB_485_U12, P3_SUB_485_U13, P3_SUB_485_U14, P3_SUB_485_U15, P3_SUB_485_U16, P3_SUB_485_U17, P3_SUB_485_U18, P3_SUB_485_U19, P3_SUB_485_U20, P3_SUB_485_U21, P3_SUB_485_U22, P3_SUB_485_U23, P3_SUB_485_U24, P3_SUB_485_U25, P3_SUB_485_U26, P3_SUB_485_U27, P3_SUB_485_U28, P3_SUB_485_U29, P3_SUB_485_U30, P3_SUB_485_U31, P3_SUB_485_U32, P3_SUB_485_U33, P3_SUB_485_U34, P3_SUB_485_U35, P3_SUB_485_U36, P3_SUB_485_U37, P3_SUB_485_U38, P3_SUB_485_U39, P3_SUB_485_U40, P3_SUB_485_U41, P3_SUB_485_U42, P3_SUB_485_U43, P3_SUB_485_U44, P3_SUB_485_U45, P3_SUB_485_U46, P3_SUB_485_U47, P3_SUB_485_U48, P3_SUB_485_U49, P3_SUB_485_U50, P3_SUB_485_U51, P3_SUB_485_U52, P3_SUB_485_U53, P3_SUB_485_U54, P3_SUB_485_U55, P3_SUB_485_U56, P3_SUB_485_U57, P3_SUB_485_U58, P3_SUB_485_U59, P3_SUB_485_U60, P3_SUB_485_U61, P3_SUB_485_U62, P3_SUB_485_U63, P3_SUB_563_U6, P3_SUB_563_U7, P3_ADD_515_U4, P3_ADD_515_U5, P3_ADD_515_U6, P3_ADD_515_U7, P3_ADD_515_U8, P3_ADD_515_U9, P3_ADD_515_U10, P3_ADD_515_U11, P3_ADD_515_U12, P3_ADD_515_U13, P3_ADD_515_U14, P3_ADD_515_U15, P3_ADD_515_U16, P3_ADD_515_U17, P3_ADD_515_U18, P3_ADD_515_U19, P3_ADD_515_U20, P3_ADD_515_U21, P3_ADD_515_U22, P3_ADD_515_U23, P3_ADD_515_U24, P3_ADD_515_U25, P3_ADD_515_U26, P3_ADD_515_U27, P3_ADD_515_U28, P3_ADD_515_U29, P3_ADD_515_U30, P3_ADD_515_U31, P3_ADD_515_U32, P3_ADD_515_U33, P3_ADD_515_U34, P3_ADD_515_U35, P3_ADD_515_U36, P3_ADD_515_U37, P3_ADD_515_U38, P3_ADD_515_U39, P3_ADD_515_U40, P3_ADD_515_U41, P3_ADD_515_U42, P3_ADD_515_U43, P3_ADD_515_U44, P3_ADD_515_U45, P3_ADD_515_U46, P3_ADD_515_U47, P3_ADD_515_U48, P3_ADD_515_U49, P3_ADD_515_U50, P3_ADD_515_U51, P3_ADD_515_U52, P3_ADD_515_U53, P3_ADD_515_U54, P3_ADD_515_U55, P3_ADD_515_U56, P3_ADD_515_U57, P3_ADD_515_U58, P3_ADD_515_U59, P3_ADD_515_U60, P3_ADD_515_U61, P3_ADD_515_U62, P3_ADD_515_U63, P3_ADD_515_U64, P3_ADD_515_U65, P3_ADD_515_U66, P3_ADD_515_U67, P3_ADD_515_U68, P3_ADD_515_U69, P3_ADD_515_U70, P3_ADD_515_U71, P3_ADD_515_U72, P3_ADD_515_U73, P3_ADD_515_U74, P3_ADD_515_U75, P3_ADD_515_U76, P3_ADD_515_U77, P3_ADD_515_U78, P3_ADD_515_U79, P3_ADD_515_U80, P3_ADD_515_U81, P3_ADD_515_U82, P3_ADD_515_U83, P3_ADD_515_U84, P3_ADD_515_U85, P3_ADD_515_U86, P3_ADD_515_U87, P3_ADD_515_U88, P3_ADD_515_U89, P3_ADD_515_U90, P3_ADD_515_U91, P3_ADD_515_U92, P3_ADD_515_U93, P3_ADD_515_U94, P3_ADD_515_U95, P3_ADD_515_U96, P3_ADD_515_U97, P3_ADD_515_U98, P3_ADD_515_U99, P3_ADD_515_U100, P3_ADD_515_U101, P3_ADD_515_U102, P3_ADD_515_U103, P3_ADD_515_U104, P3_ADD_515_U105, P3_ADD_515_U106, P3_ADD_515_U107, P3_ADD_515_U108, P3_ADD_515_U109, P3_ADD_515_U110, P3_ADD_515_U111, P3_ADD_515_U112, P3_ADD_515_U113, P3_ADD_515_U114, P3_ADD_515_U115, P3_ADD_515_U116, P3_ADD_515_U117, P3_ADD_515_U118, P3_ADD_515_U119, P3_ADD_515_U120, P3_ADD_515_U121, P3_ADD_515_U122, P3_ADD_515_U123, P3_ADD_515_U124, P3_ADD_515_U125, P3_ADD_515_U126, P3_ADD_515_U127, P3_ADD_515_U128, P3_ADD_515_U129, P3_ADD_515_U130, P3_ADD_515_U131, P3_ADD_515_U132, P3_ADD_515_U133, P3_ADD_515_U134, P3_ADD_515_U135, P3_ADD_515_U136, P3_ADD_515_U137, P3_ADD_515_U138, P3_ADD_515_U139, P3_ADD_515_U140, P3_ADD_515_U141, P3_ADD_515_U142, P3_ADD_515_U143, P3_ADD_515_U144, P3_ADD_515_U145, P3_ADD_515_U146, P3_ADD_515_U147, P3_ADD_515_U148, P3_ADD_515_U149, P3_ADD_515_U150, P3_ADD_515_U151, P3_ADD_515_U152, P3_ADD_515_U153, P3_ADD_515_U154, P3_ADD_515_U155, P3_ADD_515_U156, P3_ADD_515_U157, P3_ADD_515_U158, P3_ADD_515_U159, P3_ADD_515_U160, P3_ADD_515_U161, P3_ADD_515_U162, P3_ADD_515_U163, P3_ADD_515_U164, P3_ADD_515_U165, P3_ADD_515_U166, P3_ADD_515_U167, P3_ADD_515_U168, P3_ADD_515_U169, P3_ADD_515_U170, P3_ADD_515_U171, P3_ADD_515_U172, P3_ADD_515_U173, P3_ADD_515_U174, P3_ADD_515_U175, P3_ADD_515_U176, P3_ADD_515_U177, P3_ADD_515_U178, P3_ADD_515_U179, P3_ADD_515_U180, P3_ADD_515_U181, P3_ADD_515_U182, P3_ADD_394_U4, P3_ADD_394_U5, P3_ADD_394_U6, P3_ADD_394_U7, P3_ADD_394_U8, P3_ADD_394_U9, P3_ADD_394_U10, P3_ADD_394_U11, P3_ADD_394_U12, P3_ADD_394_U13, P3_ADD_394_U14, P3_ADD_394_U15, P3_ADD_394_U16, P3_ADD_394_U17, P3_ADD_394_U18, P3_ADD_394_U19, P3_ADD_394_U20, P3_ADD_394_U21, P3_ADD_394_U22, P3_ADD_394_U23, P3_ADD_394_U24, P3_ADD_394_U25, P3_ADD_394_U26, P3_ADD_394_U27, P3_ADD_394_U28, P3_ADD_394_U29, P3_ADD_394_U30, P3_ADD_394_U31, P3_ADD_394_U32, P3_ADD_394_U33, P3_ADD_394_U34, P3_ADD_394_U35, P3_ADD_394_U36, P3_ADD_394_U37, P3_ADD_394_U38, P3_ADD_394_U39, P3_ADD_394_U40, P3_ADD_394_U41, P3_ADD_394_U42, P3_ADD_394_U43, P3_ADD_394_U44, P3_ADD_394_U45, P3_ADD_394_U46, P3_ADD_394_U47, P3_ADD_394_U48, P3_ADD_394_U49, P3_ADD_394_U50, P3_ADD_394_U51, P3_ADD_394_U52, P3_ADD_394_U53, P3_ADD_394_U54, P3_ADD_394_U55, P3_ADD_394_U56, P3_ADD_394_U57, P3_ADD_394_U58, P3_ADD_394_U59, P3_ADD_394_U60, P3_ADD_394_U61, P3_ADD_394_U62, P3_ADD_394_U63, P3_ADD_394_U64, P3_ADD_394_U65, P3_ADD_394_U66, P3_ADD_394_U67, P3_ADD_394_U68, P3_ADD_394_U69, P3_ADD_394_U70, P3_ADD_394_U71, P3_ADD_394_U72, P3_ADD_394_U73, P3_ADD_394_U74, P3_ADD_394_U75, P3_ADD_394_U76, P3_ADD_394_U77, P3_ADD_394_U78, P3_ADD_394_U79, P3_ADD_394_U80, P3_ADD_394_U81, P3_ADD_394_U82, P3_ADD_394_U83, P3_ADD_394_U84, P3_ADD_394_U85, P3_ADD_394_U86, P3_ADD_394_U87, P3_ADD_394_U88, P3_ADD_394_U89, P3_ADD_394_U90, P3_ADD_394_U91, P3_ADD_394_U92, P3_ADD_394_U93, P3_ADD_394_U94, P3_ADD_394_U95, P3_ADD_394_U96, P3_ADD_394_U97, P3_ADD_394_U98, P3_ADD_394_U99, P3_ADD_394_U100, P3_ADD_394_U101, P3_ADD_394_U102, P3_ADD_394_U103, P3_ADD_394_U104, P3_ADD_394_U105, P3_ADD_394_U106, P3_ADD_394_U107, P3_ADD_394_U108, P3_ADD_394_U109, P3_ADD_394_U110, P3_ADD_394_U111, P3_ADD_394_U112, P3_ADD_394_U113, P3_ADD_394_U114, P3_ADD_394_U115, P3_ADD_394_U116, P3_ADD_394_U117, P3_ADD_394_U118, P3_ADD_394_U119, P3_ADD_394_U120, P3_ADD_394_U121, P3_ADD_394_U122, P3_ADD_394_U123, P3_ADD_394_U124, P3_ADD_394_U125, P3_ADD_394_U126, P3_ADD_394_U127, P3_ADD_394_U128, P3_ADD_394_U129, P3_ADD_394_U130, P3_ADD_394_U131, P3_ADD_394_U132, P3_ADD_394_U133, P3_ADD_394_U134, P3_ADD_394_U135, P3_ADD_394_U136, P3_ADD_394_U137, P3_ADD_394_U138, P3_ADD_394_U139, P3_ADD_394_U140, P3_ADD_394_U141, P3_ADD_394_U142, P3_ADD_394_U143, P3_ADD_394_U144, P3_ADD_394_U145, P3_ADD_394_U146, P3_ADD_394_U147, P3_ADD_394_U148, P3_ADD_394_U149, P3_ADD_394_U150, P3_ADD_394_U151, P3_ADD_394_U152, P3_ADD_394_U153, P3_ADD_394_U154, P3_ADD_394_U155, P3_ADD_394_U156, P3_ADD_394_U157, P3_ADD_394_U158, P3_ADD_394_U159, P3_ADD_394_U160, P3_ADD_394_U161, P3_ADD_394_U162, P3_ADD_394_U163, P3_ADD_394_U164, P3_ADD_394_U165, P3_ADD_394_U166, P3_ADD_394_U167, P3_ADD_394_U168, P3_ADD_394_U169, P3_ADD_394_U170, P3_ADD_394_U171, P3_ADD_394_U172, P3_ADD_394_U173, P3_ADD_394_U174, P3_ADD_394_U175, P3_ADD_394_U176, P3_ADD_394_U177, P3_ADD_394_U178, P3_ADD_394_U179, P3_ADD_394_U180, P3_ADD_394_U181, P3_ADD_394_U182, P3_ADD_394_U183, P3_ADD_394_U184, P3_ADD_394_U185, P3_ADD_394_U186, P3_GTE_450_U6, P3_GTE_450_U7, P3_SUB_414_U6, P3_SUB_414_U7, P3_SUB_414_U8, P3_SUB_414_U9, P3_SUB_414_U10, P3_SUB_414_U11, P3_SUB_414_U12, P3_SUB_414_U13, P3_SUB_414_U14, P3_SUB_414_U15, P3_SUB_414_U16, P3_SUB_414_U17, P3_SUB_414_U18, P3_SUB_414_U19, P3_SUB_414_U20, P3_SUB_414_U21, P3_SUB_414_U22, P3_SUB_414_U23, P3_SUB_414_U24, P3_SUB_414_U25, P3_SUB_414_U26, P3_SUB_414_U27, P3_SUB_414_U28, P3_SUB_414_U29, P3_SUB_414_U30, P3_SUB_414_U31, P3_SUB_414_U32, P3_SUB_414_U33, P3_SUB_414_U34, P3_SUB_414_U35, P3_SUB_414_U36, P3_SUB_414_U37, P3_SUB_414_U38, P3_SUB_414_U39, P3_SUB_414_U40, P3_SUB_414_U41, P3_SUB_414_U42, P3_SUB_414_U43, P3_SUB_414_U44, P3_SUB_414_U45, P3_SUB_414_U46, P3_SUB_414_U47, P3_SUB_414_U48, P3_SUB_414_U49, P3_SUB_414_U50, P3_SUB_414_U51, P3_SUB_414_U52, P3_SUB_414_U53, P3_SUB_414_U54, P3_SUB_414_U55, P3_SUB_414_U56, P3_SUB_414_U57, P3_SUB_414_U58, P3_SUB_414_U59, P3_SUB_414_U60, P3_SUB_414_U61, P3_SUB_414_U62, P3_SUB_414_U63, P3_SUB_414_U64, P3_SUB_414_U65, P3_SUB_414_U66, P3_SUB_414_U67, P3_SUB_414_U68, P3_SUB_414_U69, P3_SUB_414_U70, P3_SUB_414_U71, P3_SUB_414_U72, P3_SUB_414_U73, P3_SUB_414_U74, P3_SUB_414_U75, P3_SUB_414_U76, P3_SUB_414_U77, P3_SUB_414_U78, P3_SUB_414_U79, P3_SUB_414_U80, P3_SUB_414_U81, P3_SUB_414_U82, P3_SUB_414_U83, P3_SUB_414_U84, P3_SUB_414_U85, P3_SUB_414_U86, P3_SUB_414_U87, P3_SUB_414_U88, P3_SUB_414_U89, P3_SUB_414_U90, P3_SUB_414_U91, P3_SUB_414_U92, P3_SUB_414_U93, P3_SUB_414_U94, P3_SUB_414_U95, P3_SUB_414_U96, P3_SUB_414_U97, P3_SUB_414_U98, P3_SUB_414_U99, P3_SUB_414_U100, P3_SUB_414_U101, P3_SUB_414_U102, P3_SUB_414_U103, P3_SUB_414_U104, P3_SUB_414_U105, P3_SUB_414_U106, P3_SUB_414_U107, P3_SUB_414_U108, P3_SUB_414_U109, P3_SUB_414_U110, P3_SUB_414_U111, P3_SUB_414_U112, P3_SUB_414_U113, P3_SUB_414_U114, P3_SUB_414_U115, P3_SUB_414_U116, P3_SUB_414_U117, P3_SUB_414_U118, P3_SUB_414_U119, P3_SUB_414_U120, P3_SUB_414_U121, P3_SUB_414_U122, P3_SUB_414_U123, P3_SUB_414_U124, P3_SUB_414_U125, P3_SUB_414_U126, P3_SUB_414_U127, P3_SUB_414_U128, P3_SUB_414_U129, P3_SUB_414_U130, P3_SUB_414_U131, P3_SUB_414_U132, P3_SUB_414_U133, P3_SUB_414_U134, P3_SUB_414_U135, P3_SUB_414_U136, P3_SUB_414_U137, P3_SUB_414_U138, P3_SUB_414_U139, P3_SUB_414_U140, P3_SUB_414_U141, P3_SUB_414_U142, P3_SUB_414_U143, P3_SUB_414_U144, P3_SUB_414_U145, P3_SUB_414_U146, P3_SUB_414_U147, P3_SUB_414_U148, P3_SUB_414_U149, P3_SUB_414_U150, P3_SUB_414_U151, P3_SUB_414_U152, P3_SUB_414_U153, P3_SUB_414_U154, P3_SUB_414_U155, P3_SUB_414_U156, P3_SUB_414_U157, P3_SUB_414_U158, P3_SUB_414_U159, P3_ADD_441_U4, P3_ADD_441_U5, P3_ADD_441_U6, P3_ADD_441_U7, P3_ADD_441_U8, P3_ADD_441_U9, P3_ADD_441_U10, P3_ADD_441_U11, P3_ADD_441_U12, P3_ADD_441_U13, P3_ADD_441_U14, P3_ADD_441_U15, P3_ADD_441_U16, P3_ADD_441_U17, P3_ADD_441_U18, P3_ADD_441_U19, P3_ADD_441_U20, P3_ADD_441_U21, P3_ADD_441_U22, P3_ADD_441_U23, P3_ADD_441_U24, P3_ADD_441_U25, P3_ADD_441_U26, P3_ADD_441_U27, P3_ADD_441_U28, P3_ADD_441_U29, P3_ADD_441_U30, P3_ADD_441_U31, P3_ADD_441_U32, P3_ADD_441_U33, P3_ADD_441_U34, P3_ADD_441_U35, P3_ADD_441_U36, P3_ADD_441_U37, P3_ADD_441_U38, P3_ADD_441_U39, P3_ADD_441_U40, P3_ADD_441_U41, P3_ADD_441_U42, P3_ADD_441_U43, P3_ADD_441_U44, P3_ADD_441_U45, P3_ADD_441_U46, P3_ADD_441_U47, P3_ADD_441_U48, P3_ADD_441_U49, P3_ADD_441_U50, P3_ADD_441_U51, P3_ADD_441_U52, P3_ADD_441_U53, P3_ADD_441_U54, P3_ADD_441_U55, P3_ADD_441_U56, P3_ADD_441_U57, P3_ADD_441_U58, P3_ADD_441_U59, P3_ADD_441_U60, P3_ADD_441_U61, P3_ADD_441_U62, P3_ADD_441_U63, P3_ADD_441_U64, P3_ADD_441_U65, P3_ADD_441_U66, P3_ADD_441_U67, P3_ADD_441_U68, P3_ADD_441_U69, P3_ADD_441_U70, P3_ADD_441_U71, P3_ADD_441_U72, P3_ADD_441_U73, P3_ADD_441_U74, P3_ADD_441_U75, P3_ADD_441_U76, P3_ADD_441_U77, P3_ADD_441_U78, P3_ADD_441_U79, P3_ADD_441_U80, P3_ADD_441_U81, P3_ADD_441_U82, P3_ADD_441_U83, P3_ADD_441_U84, P3_ADD_441_U85, P3_ADD_441_U86, P3_ADD_441_U87, P3_ADD_441_U88, P3_ADD_441_U89, P3_ADD_441_U90, P3_ADD_441_U91, P3_ADD_441_U92, P3_ADD_441_U93, P3_ADD_441_U94, P3_ADD_441_U95, P3_ADD_441_U96, P3_ADD_441_U97, P3_ADD_441_U98, P3_ADD_441_U99, P3_ADD_441_U100, P3_ADD_441_U101, P3_ADD_441_U102, P3_ADD_441_U103, P3_ADD_441_U104, P3_ADD_441_U105, P3_ADD_441_U106, P3_ADD_441_U107, P3_ADD_441_U108, P3_ADD_441_U109, P3_ADD_441_U110, P3_ADD_441_U111, P3_ADD_441_U112, P3_ADD_441_U113, P3_ADD_441_U114, P3_ADD_441_U115, P3_ADD_441_U116, P3_ADD_441_U117, P3_ADD_441_U118, P3_ADD_441_U119, P3_ADD_441_U120, P3_ADD_441_U121, P3_ADD_441_U122, P3_ADD_441_U123, P3_ADD_441_U124, P3_ADD_441_U125, P3_ADD_441_U126, P3_ADD_441_U127, P3_ADD_441_U128, P3_ADD_441_U129, P3_ADD_441_U130, P3_ADD_441_U131, P3_ADD_441_U132, P3_ADD_441_U133, P3_ADD_441_U134, P3_ADD_441_U135, P3_ADD_441_U136, P3_ADD_441_U137, P3_ADD_441_U138, P3_ADD_441_U139, P3_ADD_441_U140, P3_ADD_441_U141, P3_ADD_441_U142, P3_ADD_441_U143, P3_ADD_441_U144, P3_ADD_441_U145, P3_ADD_441_U146, P3_ADD_441_U147, P3_ADD_441_U148, P3_ADD_441_U149, P3_ADD_441_U150, P3_ADD_441_U151, P3_ADD_441_U152, P3_ADD_441_U153, P3_ADD_441_U154, P3_ADD_441_U155, P3_ADD_441_U156, P3_ADD_441_U157, P3_ADD_441_U158, P3_ADD_441_U159, P3_ADD_441_U160, P3_ADD_441_U161, P3_ADD_441_U162, P3_ADD_441_U163, P3_ADD_441_U164, P3_ADD_441_U165, P3_ADD_441_U166, P3_ADD_441_U167, P3_ADD_441_U168, P3_ADD_441_U169, P3_ADD_441_U170, P3_ADD_441_U171, P3_ADD_441_U172, P3_ADD_441_U173, P3_ADD_441_U174, P3_ADD_441_U175, P3_ADD_441_U176, P3_ADD_441_U177, P3_ADD_441_U178, P3_ADD_441_U179, P3_ADD_441_U180, P3_ADD_441_U181, P3_ADD_441_U182, P3_ADD_349_U5, P3_ADD_349_U6, P3_ADD_349_U7, P3_ADD_349_U8, P3_ADD_349_U9, P3_ADD_349_U10, P3_ADD_349_U11, P3_ADD_349_U12, P3_ADD_349_U13, P3_ADD_349_U14, P3_ADD_349_U15, P3_ADD_349_U16, P3_ADD_349_U17, P3_ADD_349_U18, P3_ADD_349_U19, P3_ADD_349_U20, P3_ADD_349_U21, P3_ADD_349_U22, P3_ADD_349_U23, P3_ADD_349_U24, P3_ADD_349_U25, P3_ADD_349_U26, P3_ADD_349_U27, P3_ADD_349_U28, P3_ADD_349_U29, P3_ADD_349_U30, P3_ADD_349_U31, P3_ADD_349_U32, P3_ADD_349_U33, P3_ADD_349_U34, P3_ADD_349_U35, P3_ADD_349_U36, P3_ADD_349_U37, P3_ADD_349_U38, P3_ADD_349_U39, P3_ADD_349_U40, P3_ADD_349_U41, P3_ADD_349_U42, P3_ADD_349_U43, P3_ADD_349_U44, P3_ADD_349_U45, P3_ADD_349_U46, P3_ADD_349_U47, P3_ADD_349_U48, P3_ADD_349_U49, P3_ADD_349_U50, P3_ADD_349_U51, P3_ADD_349_U52, P3_ADD_349_U53, P3_ADD_349_U54, P3_ADD_349_U55, P3_ADD_349_U56, P3_ADD_349_U57, P3_ADD_349_U58, P3_ADD_349_U59, P3_ADD_349_U60, P3_ADD_349_U61, P3_ADD_349_U62, P3_ADD_349_U63, P3_ADD_349_U64, P3_ADD_349_U65, P3_ADD_349_U66, P3_ADD_349_U67, P3_ADD_349_U68, P3_ADD_349_U69, P3_ADD_349_U70, P3_ADD_349_U71, P3_ADD_349_U72, P3_ADD_349_U73, P3_ADD_349_U74, P3_ADD_349_U75, P3_ADD_349_U76, P3_ADD_349_U77, P3_ADD_349_U78, P3_ADD_349_U79, P3_ADD_349_U80, P3_ADD_349_U81, P3_ADD_349_U82, P3_ADD_349_U83, P3_ADD_349_U84, P3_ADD_349_U85, P3_ADD_349_U86, P3_ADD_349_U87, P3_ADD_349_U88, P3_ADD_349_U89, P3_ADD_349_U90, P3_ADD_349_U91, P3_ADD_349_U92, P3_ADD_349_U93, P3_ADD_349_U94, P3_ADD_349_U95, P3_ADD_349_U96, P3_ADD_349_U97, P3_ADD_349_U98, P3_ADD_349_U99, P3_ADD_349_U100, P3_ADD_349_U101, P3_ADD_349_U102, P3_ADD_349_U103, P3_ADD_349_U104, P3_ADD_349_U105, P3_ADD_349_U106, P3_ADD_349_U107, P3_ADD_349_U108, P3_ADD_349_U109, P3_ADD_349_U110, P3_ADD_349_U111, P3_ADD_349_U112, P3_ADD_349_U113, P3_ADD_349_U114, P3_ADD_349_U115, P3_ADD_349_U116, P3_ADD_349_U117, P3_ADD_349_U118, P3_ADD_349_U119, P3_ADD_349_U120, P3_ADD_349_U121, P3_ADD_349_U122, P3_ADD_349_U123, P3_ADD_349_U124, P3_ADD_349_U125, P3_ADD_349_U126, P3_ADD_349_U127, P3_ADD_349_U128, P3_ADD_349_U129, P3_ADD_349_U130, P3_ADD_349_U131, P3_ADD_349_U132, P3_ADD_349_U133, P3_ADD_349_U134, P3_ADD_349_U135, P3_ADD_349_U136, P3_ADD_349_U137, P3_ADD_349_U138, P3_ADD_349_U139, P3_ADD_349_U140, P3_ADD_349_U141, P3_ADD_349_U142, P3_ADD_349_U143, P3_ADD_349_U144, P3_ADD_349_U145, P3_ADD_349_U146, P3_ADD_349_U147, P3_ADD_349_U148, P3_ADD_349_U149, P3_ADD_349_U150, P3_ADD_349_U151, P3_ADD_349_U152, P3_ADD_349_U153, P3_ADD_349_U154, P3_ADD_349_U155, P3_ADD_349_U156, P3_ADD_349_U157, P3_ADD_349_U158, P3_ADD_349_U159, P3_ADD_349_U160, P3_ADD_349_U161, P3_ADD_349_U162, P3_ADD_349_U163, P3_ADD_349_U164, P3_ADD_349_U165, P3_ADD_349_U166, P3_ADD_349_U167, P3_ADD_349_U168, P3_ADD_349_U169, P3_ADD_349_U170, P3_ADD_349_U171, P3_ADD_349_U172, P3_ADD_349_U173, P3_ADD_349_U174, P3_ADD_349_U175, P3_ADD_349_U176, P3_ADD_349_U177, P3_ADD_349_U178, P3_ADD_349_U179, P3_ADD_349_U180, P3_ADD_349_U181, P3_ADD_349_U182, P3_ADD_349_U183, P3_ADD_349_U184, P3_ADD_349_U185, P3_ADD_349_U186, P3_ADD_349_U187, P3_ADD_349_U188, P3_ADD_349_U189, P3_ADD_405_U4, P3_ADD_405_U5, P3_ADD_405_U6, P3_ADD_405_U7, P3_ADD_405_U8, P3_ADD_405_U9, P3_ADD_405_U10, P3_ADD_405_U11, P3_ADD_405_U12, P3_ADD_405_U13, P3_ADD_405_U14, P3_ADD_405_U15, P3_ADD_405_U16, P3_ADD_405_U17, P3_ADD_405_U18, P3_ADD_405_U19, P3_ADD_405_U20, P3_ADD_405_U21, P3_ADD_405_U22, P3_ADD_405_U23, P3_ADD_405_U24, P3_ADD_405_U25, P3_ADD_405_U26, P3_ADD_405_U27, P3_ADD_405_U28, P3_ADD_405_U29, P3_ADD_405_U30, P3_ADD_405_U31, P3_ADD_405_U32, P3_ADD_405_U33, P3_ADD_405_U34, P3_ADD_405_U35, P3_ADD_405_U36, P3_ADD_405_U37, P3_ADD_405_U38, P3_ADD_405_U39, P3_ADD_405_U40, P3_ADD_405_U41, P3_ADD_405_U42, P3_ADD_405_U43, P3_ADD_405_U44, P3_ADD_405_U45, P3_ADD_405_U46, P3_ADD_405_U47, P3_ADD_405_U48, P3_ADD_405_U49, P3_ADD_405_U50, P3_ADD_405_U51, P3_ADD_405_U52, P3_ADD_405_U53, P3_ADD_405_U54, P3_ADD_405_U55, P3_ADD_405_U56, P3_ADD_405_U57, P3_ADD_405_U58, P3_ADD_405_U59, P3_ADD_405_U60, P3_ADD_405_U61, P3_ADD_405_U62, P3_ADD_405_U63, P3_ADD_405_U64, P3_ADD_405_U65, P3_ADD_405_U66, P3_ADD_405_U67, P3_ADD_405_U68, P3_ADD_405_U69, P3_ADD_405_U70, P3_ADD_405_U71, P3_ADD_405_U72, P3_ADD_405_U73, P3_ADD_405_U74, P3_ADD_405_U75, P3_ADD_405_U76, P3_ADD_405_U77, P3_ADD_405_U78, P3_ADD_405_U79, P3_ADD_405_U80, P3_ADD_405_U81, P3_ADD_405_U82, P3_ADD_405_U83, P3_ADD_405_U84, P3_ADD_405_U85, P3_ADD_405_U86, P3_ADD_405_U87, P3_ADD_405_U88, P3_ADD_405_U89, P3_ADD_405_U90, P3_ADD_405_U91, P3_ADD_405_U92, P3_ADD_405_U93, P3_ADD_405_U94, P3_ADD_405_U95, P3_ADD_405_U96, P3_ADD_405_U97, P3_ADD_405_U98, P3_ADD_405_U99, P3_ADD_405_U100, P3_ADD_405_U101, P3_ADD_405_U102, P3_ADD_405_U103, P3_ADD_405_U104, P3_ADD_405_U105, P3_ADD_405_U106, P3_ADD_405_U107, P3_ADD_405_U108, P3_ADD_405_U109, P3_ADD_405_U110, P3_ADD_405_U111, P3_ADD_405_U112, P3_ADD_405_U113, P3_ADD_405_U114, P3_ADD_405_U115, P3_ADD_405_U116, P3_ADD_405_U117, P3_ADD_405_U118, P3_ADD_405_U119, P3_ADD_405_U120, P3_ADD_405_U121, P3_ADD_405_U122, P3_ADD_405_U123, P3_ADD_405_U124, P3_ADD_405_U125, P3_ADD_405_U126, P3_ADD_405_U127, P3_ADD_405_U128, P3_ADD_405_U129, P3_ADD_405_U130, P3_ADD_405_U131, P3_ADD_405_U132, P3_ADD_405_U133, P3_ADD_405_U134, P3_ADD_405_U135, P3_ADD_405_U136, P3_ADD_405_U137, P3_ADD_405_U138, P3_ADD_405_U139, P3_ADD_405_U140, P3_ADD_405_U141, P3_ADD_405_U142, P3_ADD_405_U143, P3_ADD_405_U144, P3_ADD_405_U145, P3_ADD_405_U146, P3_ADD_405_U147, P3_ADD_405_U148, P3_ADD_405_U149, P3_ADD_405_U150, P3_ADD_405_U151, P3_ADD_405_U152, P3_ADD_405_U153, P3_ADD_405_U154, P3_ADD_405_U155, P3_ADD_405_U156, P3_ADD_405_U157, P3_ADD_405_U158, P3_ADD_405_U159, P3_ADD_405_U160, P3_ADD_405_U161, P3_ADD_405_U162, P3_ADD_405_U163, P3_ADD_405_U164, P3_ADD_405_U165, P3_ADD_405_U166, P3_ADD_405_U167, P3_ADD_405_U168, P3_ADD_405_U169, P3_ADD_405_U170, P3_ADD_405_U171, P3_ADD_405_U172, P3_ADD_405_U173, P3_ADD_405_U174, P3_ADD_405_U175, P3_ADD_405_U176, P3_ADD_405_U177, P3_ADD_405_U178, P3_ADD_405_U179, P3_ADD_405_U180, P3_ADD_405_U181, P3_ADD_405_U182, P3_ADD_405_U183, P3_ADD_405_U184, P3_ADD_405_U185, P3_ADD_405_U186, P3_ADD_553_U5, P3_ADD_553_U6, P3_ADD_553_U7, P3_ADD_553_U8, P3_ADD_553_U9, P3_ADD_553_U10, P3_ADD_553_U11, P3_ADD_553_U12, P3_ADD_553_U13, P3_ADD_553_U14, P3_ADD_553_U15, P3_ADD_553_U16, P3_ADD_553_U17, P3_ADD_553_U18, P3_ADD_553_U19, P3_ADD_553_U20, P3_ADD_553_U21, P3_ADD_553_U22, P3_ADD_553_U23, P3_ADD_553_U24, P3_ADD_553_U25, P3_ADD_553_U26, P3_ADD_553_U27, P3_ADD_553_U28, P3_ADD_553_U29, P3_ADD_553_U30, P3_ADD_553_U31, P3_ADD_553_U32, P3_ADD_553_U33, P3_ADD_553_U34, P3_ADD_553_U35, P3_ADD_553_U36, P3_ADD_553_U37, P3_ADD_553_U38, P3_ADD_553_U39, P3_ADD_553_U40, P3_ADD_553_U41, P3_ADD_553_U42, P3_ADD_553_U43, P3_ADD_553_U44, P3_ADD_553_U45, P3_ADD_553_U46, P3_ADD_553_U47, P3_ADD_553_U48, P3_ADD_553_U49, P3_ADD_553_U50, P3_ADD_553_U51, P3_ADD_553_U52, P3_ADD_553_U53, P3_ADD_553_U54, P3_ADD_553_U55, P3_ADD_553_U56, P3_ADD_553_U57, P3_ADD_553_U58, P3_ADD_553_U59, P3_ADD_553_U60, P3_ADD_553_U61, P3_ADD_553_U62, P3_ADD_553_U63, P3_ADD_553_U64, P3_ADD_553_U65, P3_ADD_553_U66, P3_ADD_553_U67, P3_ADD_553_U68, P3_ADD_553_U69, P3_ADD_553_U70, P3_ADD_553_U71, P3_ADD_553_U72, P3_ADD_553_U73, P3_ADD_553_U74, P3_ADD_553_U75, P3_ADD_553_U76, P3_ADD_553_U77, P3_ADD_553_U78, P3_ADD_553_U79, P3_ADD_553_U80, P3_ADD_553_U81, P3_ADD_553_U82, P3_ADD_553_U83, P3_ADD_553_U84, P3_ADD_553_U85, P3_ADD_553_U86, P3_ADD_553_U87, P3_ADD_553_U88, P3_ADD_553_U89, P3_ADD_553_U90, P3_ADD_553_U91, P3_ADD_553_U92, P3_ADD_553_U93, P3_ADD_553_U94, P3_ADD_553_U95, P3_ADD_553_U96, P3_ADD_553_U97, P3_ADD_553_U98, P3_ADD_553_U99, P3_ADD_553_U100, P3_ADD_553_U101, P3_ADD_553_U102, P3_ADD_553_U103, P3_ADD_553_U104, P3_ADD_553_U105, P3_ADD_553_U106, P3_ADD_553_U107, P3_ADD_553_U108, P3_ADD_553_U109, P3_ADD_553_U110, P3_ADD_553_U111, P3_ADD_553_U112, P3_ADD_553_U113, P3_ADD_553_U114, P3_ADD_553_U115, P3_ADD_553_U116, P3_ADD_553_U117, P3_ADD_553_U118, P3_ADD_553_U119, P3_ADD_553_U120, P3_ADD_553_U121, P3_ADD_553_U122, P3_ADD_553_U123, P3_ADD_553_U124, P3_ADD_553_U125, P3_ADD_553_U126, P3_ADD_553_U127, P3_ADD_553_U128, P3_ADD_553_U129, P3_ADD_553_U130, P3_ADD_553_U131, P3_ADD_553_U132, P3_ADD_553_U133, P3_ADD_553_U134, P3_ADD_553_U135, P3_ADD_553_U136, P3_ADD_553_U137, P3_ADD_553_U138, P3_ADD_553_U139, P3_ADD_553_U140, P3_ADD_553_U141, P3_ADD_553_U142, P3_ADD_553_U143, P3_ADD_553_U144, P3_ADD_553_U145, P3_ADD_553_U146, P3_ADD_553_U147, P3_ADD_553_U148, P3_ADD_553_U149, P3_ADD_553_U150, P3_ADD_553_U151, P3_ADD_553_U152, P3_ADD_553_U153, P3_ADD_553_U154, P3_ADD_553_U155, P3_ADD_553_U156, P3_ADD_553_U157, P3_ADD_553_U158, P3_ADD_553_U159, P3_ADD_553_U160, P3_ADD_553_U161, P3_ADD_553_U162, P3_ADD_553_U163, P3_ADD_553_U164, P3_ADD_553_U165, P3_ADD_553_U166, P3_ADD_553_U167, P3_ADD_553_U168, P3_ADD_553_U169, P3_ADD_553_U170, P3_ADD_553_U171, P3_ADD_553_U172, P3_ADD_553_U173, P3_ADD_553_U174, P3_ADD_553_U175, P3_ADD_553_U176, P3_ADD_553_U177, P3_ADD_553_U178, P3_ADD_553_U179, P3_ADD_553_U180, P3_ADD_553_U181, P3_ADD_553_U182, P3_ADD_553_U183, P3_ADD_553_U184, P3_ADD_553_U185, P3_ADD_553_U186, P3_ADD_553_U187, P3_ADD_553_U188, P3_ADD_553_U189, P3_ADD_558_U5, P3_ADD_558_U6, P3_ADD_558_U7, P3_ADD_558_U8, P3_ADD_558_U9, P3_ADD_558_U10, P3_ADD_558_U11, P3_ADD_558_U12, P3_ADD_558_U13, P3_ADD_558_U14, P3_ADD_558_U15, P3_ADD_558_U16, P3_ADD_558_U17, P3_ADD_558_U18, P3_ADD_558_U19, P3_ADD_558_U20, P3_ADD_558_U21, P3_ADD_558_U22, P3_ADD_558_U23, P3_ADD_558_U24, P3_ADD_558_U25, P3_ADD_558_U26, P3_ADD_558_U27, P3_ADD_558_U28, P3_ADD_558_U29, P3_ADD_558_U30, P3_ADD_558_U31, P3_ADD_558_U32, P3_ADD_558_U33, P3_ADD_558_U34, P3_ADD_558_U35, P3_ADD_558_U36, P3_ADD_558_U37, P3_ADD_558_U38, P3_ADD_558_U39, P3_ADD_558_U40, P3_ADD_558_U41, P3_ADD_558_U42, P3_ADD_558_U43, P3_ADD_558_U44, P3_ADD_558_U45, P3_ADD_558_U46, P3_ADD_558_U47, P3_ADD_558_U48, P3_ADD_558_U49, P3_ADD_558_U50, P3_ADD_558_U51, P3_ADD_558_U52, P3_ADD_558_U53, P3_ADD_558_U54, P3_ADD_558_U55, P3_ADD_558_U56, P3_ADD_558_U57, P3_ADD_558_U58, P3_ADD_558_U59, P3_ADD_558_U60, P3_ADD_558_U61, P3_ADD_558_U62, P3_ADD_558_U63, P3_ADD_558_U64, P3_ADD_558_U65, P3_ADD_558_U66, P3_ADD_558_U67, P3_ADD_558_U68, P3_ADD_558_U69, P3_ADD_558_U70, P3_ADD_558_U71, P3_ADD_558_U72, P3_ADD_558_U73, P3_ADD_558_U74, P3_ADD_558_U75, P3_ADD_558_U76, P3_ADD_558_U77, P3_ADD_558_U78, P3_ADD_558_U79, P3_ADD_558_U80, P3_ADD_558_U81, P3_ADD_558_U82, P3_ADD_558_U83, P3_ADD_558_U84, P3_ADD_558_U85, P3_ADD_558_U86, P3_ADD_558_U87, P3_ADD_558_U88, P3_ADD_558_U89, P3_ADD_558_U90, P3_ADD_558_U91, P3_ADD_558_U92, P3_ADD_558_U93, P3_ADD_558_U94, P3_ADD_558_U95, P3_ADD_558_U96, P3_ADD_558_U97, P3_ADD_558_U98, P3_ADD_558_U99, P3_ADD_558_U100, P3_ADD_558_U101, P3_ADD_558_U102, P3_ADD_558_U103, P3_ADD_558_U104, P3_ADD_558_U105, P3_ADD_558_U106, P3_ADD_558_U107, P3_ADD_558_U108, P3_ADD_558_U109, P3_ADD_558_U110, P3_ADD_558_U111, P3_ADD_558_U112, P3_ADD_558_U113, P3_ADD_558_U114, P3_ADD_558_U115, P3_ADD_558_U116, P3_ADD_558_U117, P3_ADD_558_U118, P3_ADD_558_U119, P3_ADD_558_U120, P3_ADD_558_U121, P3_ADD_558_U122, P3_ADD_558_U123, P3_ADD_558_U124, P3_ADD_558_U125, P3_ADD_558_U126, P3_ADD_558_U127, P3_ADD_558_U128, P3_ADD_558_U129, P3_ADD_558_U130, P3_ADD_558_U131, P3_ADD_558_U132, P3_ADD_558_U133, P3_ADD_558_U134, P3_ADD_558_U135, P3_ADD_558_U136, P3_ADD_558_U137, P3_ADD_558_U138, P3_ADD_558_U139, P3_ADD_558_U140, P3_ADD_558_U141, P3_ADD_558_U142, P3_ADD_558_U143, P3_ADD_558_U144, P3_ADD_558_U145, P3_ADD_558_U146, P3_ADD_558_U147, P3_ADD_558_U148, P3_ADD_558_U149, P3_ADD_558_U150, P3_ADD_558_U151, P3_ADD_558_U152, P3_ADD_558_U153, P3_ADD_558_U154, P3_ADD_558_U155, P3_ADD_558_U156, P3_ADD_558_U157, P3_ADD_558_U158, P3_ADD_558_U159, P3_ADD_558_U160, P3_ADD_558_U161, P3_ADD_558_U162, P3_ADD_558_U163, P3_ADD_558_U164, P3_ADD_558_U165, P3_ADD_558_U166, P3_ADD_558_U167, P3_ADD_558_U168, P3_ADD_558_U169, P3_ADD_558_U170, P3_ADD_558_U171, P3_ADD_558_U172, P3_ADD_558_U173, P3_ADD_558_U174, P3_ADD_558_U175, P3_ADD_558_U176, P3_ADD_558_U177, P3_ADD_558_U178, P3_ADD_558_U179, P3_ADD_558_U180, P3_ADD_558_U181, P3_ADD_558_U182, P3_ADD_558_U183, P3_ADD_558_U184, P3_ADD_558_U185, P3_ADD_558_U186, P3_ADD_558_U187, P3_ADD_558_U188, P3_ADD_558_U189, P3_ADD_385_U5, P3_ADD_385_U6, P3_ADD_385_U7, P3_ADD_385_U8, P3_ADD_385_U9, P3_ADD_385_U10, P3_ADD_385_U11, P3_ADD_385_U12, P3_ADD_385_U13, P3_ADD_385_U14, P3_ADD_385_U15, P3_ADD_385_U16, P3_ADD_385_U17, P3_ADD_385_U18, P3_ADD_385_U19, P3_ADD_385_U20, P3_ADD_385_U21, P3_ADD_385_U22, P3_ADD_385_U23, P3_ADD_385_U24, P3_ADD_385_U25, P3_ADD_385_U26, P3_ADD_385_U27, P3_ADD_385_U28, P3_ADD_385_U29, P3_ADD_385_U30, P3_ADD_385_U31, P3_ADD_385_U32, P3_ADD_385_U33, P3_ADD_385_U34, P3_ADD_385_U35, P3_ADD_385_U36, P3_ADD_385_U37, P3_ADD_385_U38, P3_ADD_385_U39, P3_ADD_385_U40, P3_ADD_385_U41, P3_ADD_385_U42, P3_ADD_385_U43, P3_ADD_385_U44, P3_ADD_385_U45, P3_ADD_385_U46, P3_ADD_385_U47, P3_ADD_385_U48, P3_ADD_385_U49, P3_ADD_385_U50, P3_ADD_385_U51, P3_ADD_385_U52, P3_ADD_385_U53, P3_ADD_385_U54, P3_ADD_385_U55, P3_ADD_385_U56, P3_ADD_385_U57, P3_ADD_385_U58, P3_ADD_385_U59, P3_ADD_385_U60, P3_ADD_385_U61, P3_ADD_385_U62, P3_ADD_385_U63, P3_ADD_385_U64, P3_ADD_385_U65, P3_ADD_385_U66, P3_ADD_385_U67, P3_ADD_385_U68, P3_ADD_385_U69, P3_ADD_385_U70, P3_ADD_385_U71, P3_ADD_385_U72, P3_ADD_385_U73, P3_ADD_385_U74, P3_ADD_385_U75, P3_ADD_385_U76, P3_ADD_385_U77, P3_ADD_385_U78, P3_ADD_385_U79, P3_ADD_385_U80, P3_ADD_385_U81, P3_ADD_385_U82, P3_ADD_385_U83, P3_ADD_385_U84, P3_ADD_385_U85, P3_ADD_385_U86, P3_ADD_385_U87, P3_ADD_385_U88, P3_ADD_385_U89, P3_ADD_385_U90, P3_ADD_385_U91, P3_ADD_385_U92, P3_ADD_385_U93, P3_ADD_385_U94, P3_ADD_385_U95, P3_ADD_385_U96, P3_ADD_385_U97, P3_ADD_385_U98, P3_ADD_385_U99, P3_ADD_385_U100, P3_ADD_385_U101, P3_ADD_385_U102, P3_ADD_385_U103, P3_ADD_385_U104, P3_ADD_385_U105, P3_ADD_385_U106, P3_ADD_385_U107, P3_ADD_385_U108, P3_ADD_385_U109, P3_ADD_385_U110, P3_ADD_385_U111, P3_ADD_385_U112, P3_ADD_385_U113, P3_ADD_385_U114, P3_ADD_385_U115, P3_ADD_385_U116, P3_ADD_385_U117, P3_ADD_385_U118, P3_ADD_385_U119, P3_ADD_385_U120, P3_ADD_385_U121, P3_ADD_385_U122, P3_ADD_385_U123, P3_ADD_385_U124, P3_ADD_385_U125, P3_ADD_385_U126, P3_ADD_385_U127, P3_ADD_385_U128, P3_ADD_385_U129, P3_ADD_385_U130, P3_ADD_385_U131, P3_ADD_385_U132, P3_ADD_385_U133, P3_ADD_385_U134, P3_ADD_385_U135, P3_ADD_385_U136, P3_ADD_385_U137, P3_ADD_385_U138, P3_ADD_385_U139, P3_ADD_385_U140, P3_ADD_385_U141, P3_ADD_385_U142, P3_ADD_385_U143, P3_ADD_385_U144, P3_ADD_385_U145, P3_ADD_385_U146, P3_ADD_385_U147, P3_ADD_385_U148, P3_ADD_385_U149, P3_ADD_385_U150, P3_ADD_385_U151, P3_ADD_385_U152, P3_ADD_385_U153, P3_ADD_385_U154, P3_ADD_385_U155, P3_ADD_385_U156, P3_ADD_385_U157, P3_ADD_385_U158, P3_ADD_385_U159, P3_ADD_385_U160, P3_ADD_385_U161, P3_ADD_385_U162, P3_ADD_385_U163, P3_ADD_385_U164, P3_ADD_385_U165, P3_ADD_385_U166, P3_ADD_385_U167, P3_ADD_385_U168, P3_ADD_385_U169, P3_ADD_385_U170, P3_ADD_385_U171, P3_ADD_385_U172, P3_ADD_385_U173, P3_ADD_385_U174, P3_ADD_385_U175, P3_ADD_385_U176, P3_ADD_385_U177, P3_ADD_385_U178, P3_ADD_385_U179, P3_ADD_385_U180, P3_ADD_385_U181, P3_ADD_385_U182, P3_ADD_385_U183, P3_ADD_385_U184, P3_ADD_385_U185, P3_ADD_385_U186, P3_ADD_385_U187, P3_ADD_385_U188, P3_ADD_385_U189, P3_ADD_357_U6, P3_ADD_357_U7, P3_ADD_357_U8, P3_ADD_357_U9, P3_ADD_357_U10, P3_ADD_357_U11, P3_ADD_357_U12, P3_ADD_357_U13, P3_ADD_357_U14, P3_ADD_357_U15, P3_ADD_357_U16, P3_ADD_357_U17, P3_ADD_357_U18, P3_ADD_357_U19, P3_ADD_357_U20, P3_ADD_357_U21, P3_ADD_357_U22, P3_ADD_357_U23, P3_ADD_357_U24, P3_ADD_357_U25, P3_ADD_357_U26, P3_ADD_357_U27, P3_ADD_357_U28, P3_ADD_357_U29, P3_ADD_357_U30, P3_ADD_357_U31, P3_ADD_357_U32, P3_ADD_357_U33, P3_ADD_357_U34, P3_ADD_357_U35, P3_ADD_547_U5, P3_ADD_547_U6, P3_ADD_547_U7, P3_ADD_547_U8, P3_ADD_547_U9, P3_ADD_547_U10, P3_ADD_547_U11, P3_ADD_547_U12, P3_ADD_547_U13, P3_ADD_547_U14, P3_ADD_547_U15, P3_ADD_547_U16, P3_ADD_547_U17, P3_ADD_547_U18, P3_ADD_547_U19, P3_ADD_547_U20, P3_ADD_547_U21, P3_ADD_547_U22, P3_ADD_547_U23, P3_ADD_547_U24, P3_ADD_547_U25, P3_ADD_547_U26, P3_ADD_547_U27, P3_ADD_547_U28, P3_ADD_547_U29, P3_ADD_547_U30, P3_ADD_547_U31, P3_ADD_547_U32, P3_ADD_547_U33, P3_ADD_547_U34, P3_ADD_547_U35, P3_ADD_547_U36, P3_ADD_547_U37, P3_ADD_547_U38, P3_ADD_547_U39, P3_ADD_547_U40, P3_ADD_547_U41, P3_ADD_547_U42, P3_ADD_547_U43, P3_ADD_547_U44, P3_ADD_547_U45, P3_ADD_547_U46, P3_ADD_547_U47, P3_ADD_547_U48, P3_ADD_547_U49, P3_ADD_547_U50, P3_ADD_547_U51, P3_ADD_547_U52, P3_ADD_547_U53, P3_ADD_547_U54, P3_ADD_547_U55, P3_ADD_547_U56, P3_ADD_547_U57, P3_ADD_547_U58, P3_ADD_547_U59, P3_ADD_547_U60, P3_ADD_547_U61, P3_ADD_547_U62, P3_ADD_547_U63, P3_ADD_547_U64, P3_ADD_547_U65, P3_ADD_547_U66, P3_ADD_547_U67, P3_ADD_547_U68, P3_ADD_547_U69, P3_ADD_547_U70, P3_ADD_547_U71, P3_ADD_547_U72, P3_ADD_547_U73, P3_ADD_547_U74, P3_ADD_547_U75, P3_ADD_547_U76, P3_ADD_547_U77, P3_ADD_547_U78, P3_ADD_547_U79, P3_ADD_547_U80, P3_ADD_547_U81, P3_ADD_547_U82, P3_ADD_547_U83, P3_ADD_547_U84, P3_ADD_547_U85, P3_ADD_547_U86, P3_ADD_547_U87, P3_ADD_547_U88, P3_ADD_547_U89, P3_ADD_547_U90, P3_ADD_547_U91, P3_ADD_547_U92, P3_ADD_547_U93, P3_ADD_547_U94, P3_ADD_547_U95, P3_ADD_547_U96, P3_ADD_547_U97, P3_ADD_547_U98, P3_ADD_547_U99, P3_ADD_547_U100, P3_ADD_547_U101, P3_ADD_547_U102, P3_ADD_547_U103, P3_ADD_547_U104, P3_ADD_547_U105, P3_ADD_547_U106, P3_ADD_547_U107, P3_ADD_547_U108, P3_ADD_547_U109, P3_ADD_547_U110, P3_ADD_547_U111, P3_ADD_547_U112, P3_ADD_547_U113, P3_ADD_547_U114, P3_ADD_547_U115, P3_ADD_547_U116, P3_ADD_547_U117, P3_ADD_547_U118, P3_ADD_547_U119, P3_ADD_547_U120, P3_ADD_547_U121, P3_ADD_547_U122, P3_ADD_547_U123, P3_ADD_547_U124, P3_ADD_547_U125, P3_ADD_547_U126, P3_ADD_547_U127, P3_ADD_547_U128, P3_ADD_547_U129, P3_ADD_547_U130, P3_ADD_547_U131, P3_ADD_547_U132, P3_ADD_547_U133, P3_ADD_547_U134, P3_ADD_547_U135, P3_ADD_547_U136, P3_ADD_547_U137, P3_ADD_547_U138, P3_ADD_547_U139, P3_ADD_547_U140, P3_ADD_547_U141, P3_ADD_547_U142, P3_ADD_547_U143, P3_ADD_547_U144, P3_ADD_547_U145, P3_ADD_547_U146, P3_ADD_547_U147, P3_ADD_547_U148, P3_ADD_547_U149, P3_ADD_547_U150, P3_ADD_547_U151, P3_ADD_547_U152, P3_ADD_547_U153, P3_ADD_547_U154, P3_ADD_547_U155, P3_ADD_547_U156, P3_ADD_547_U157, P3_ADD_547_U158, P3_ADD_547_U159, P3_ADD_547_U160, P3_ADD_547_U161, P3_ADD_547_U162, P3_ADD_547_U163, P3_ADD_547_U164, P3_ADD_547_U165, P3_ADD_547_U166, P3_ADD_547_U167, P3_ADD_547_U168, P3_ADD_547_U169, P3_ADD_547_U170, P3_ADD_547_U171, P3_ADD_547_U172, P3_ADD_547_U173, P3_ADD_547_U174, P3_ADD_547_U175, P3_ADD_547_U176, P3_ADD_547_U177, P3_ADD_547_U178, P3_ADD_547_U179, P3_ADD_547_U180, P3_ADD_547_U181, P3_ADD_547_U182, P3_ADD_547_U183, P3_ADD_547_U184, P3_ADD_547_U185, P3_ADD_547_U186, P3_ADD_547_U187, P3_ADD_547_U188, P3_ADD_547_U189, P3_SUB_412_U6, P3_SUB_412_U7, P3_SUB_412_U8, P3_SUB_412_U9, P3_SUB_412_U10, P3_SUB_412_U11, P3_SUB_412_U12, P3_SUB_412_U13, P3_SUB_412_U14, P3_SUB_412_U15, P3_SUB_412_U16, P3_SUB_412_U17, P3_SUB_412_U18, P3_SUB_412_U19, P3_SUB_412_U20, P3_SUB_412_U21, P3_SUB_412_U22, P3_SUB_412_U23, P3_SUB_412_U24, P3_SUB_412_U25, P3_SUB_412_U26, P3_SUB_412_U27, P3_SUB_412_U28, P3_SUB_412_U29, P3_SUB_412_U30, P3_SUB_412_U31, P3_SUB_412_U32, P3_SUB_412_U33, P3_SUB_412_U34, P3_SUB_412_U35, P3_SUB_412_U36, P3_SUB_412_U37, P3_SUB_412_U38, P3_SUB_412_U39, P3_SUB_412_U40, P3_SUB_412_U41, P3_SUB_412_U42, P3_SUB_412_U43, P3_SUB_412_U44, P3_SUB_412_U45, P3_SUB_412_U46, P3_SUB_412_U47, P3_SUB_412_U48, P3_SUB_412_U49, P3_SUB_412_U50, P3_SUB_412_U51, P3_SUB_412_U52, P3_SUB_412_U53, P3_SUB_412_U54, P3_SUB_412_U55, P3_SUB_412_U56, P3_SUB_412_U57, P3_SUB_412_U58, P3_SUB_412_U59, P3_SUB_412_U60, P3_SUB_412_U61, P3_SUB_412_U62, P3_SUB_412_U63, P3_ADD_371_1212_U4, P3_ADD_371_1212_U5, P3_ADD_371_1212_U6, P3_ADD_371_1212_U7, P3_ADD_371_1212_U8, P3_ADD_371_1212_U9, P3_ADD_371_1212_U10, P3_ADD_371_1212_U11, P3_ADD_371_1212_U12, P3_ADD_371_1212_U13, P3_ADD_371_1212_U14, P3_ADD_371_1212_U15, P3_ADD_371_1212_U16, P3_ADD_371_1212_U17, P3_ADD_371_1212_U18, P3_ADD_371_1212_U19, P3_ADD_371_1212_U20, P3_ADD_371_1212_U21, P3_ADD_371_1212_U22, P3_ADD_371_1212_U23, P3_ADD_371_1212_U24, P3_ADD_371_1212_U25, P3_ADD_371_1212_U26, P3_ADD_371_1212_U27, P3_ADD_371_1212_U28, P3_ADD_371_1212_U29, P3_ADD_371_1212_U30, P3_ADD_371_1212_U31, P3_ADD_371_1212_U32, P3_ADD_371_1212_U33, P3_ADD_371_1212_U34, P3_ADD_371_1212_U35, P3_ADD_371_1212_U36, P3_ADD_371_1212_U37, P3_ADD_371_1212_U38, P3_ADD_371_1212_U39, P3_ADD_371_1212_U40, P3_ADD_371_1212_U41, P3_ADD_371_1212_U42, P3_ADD_371_1212_U43, P3_ADD_371_1212_U44, P3_ADD_371_1212_U45, P3_ADD_371_1212_U46, P3_ADD_371_1212_U47, P3_ADD_371_1212_U48, P3_ADD_371_1212_U49, P3_ADD_371_1212_U50, P3_ADD_371_1212_U51, P3_ADD_371_1212_U52, P3_ADD_371_1212_U53, P3_ADD_371_1212_U54, P3_ADD_371_1212_U55, P3_ADD_371_1212_U56, P3_ADD_371_1212_U57, P3_ADD_371_1212_U58, P3_ADD_371_1212_U59, P3_ADD_371_1212_U60, P3_ADD_371_1212_U61, P3_ADD_371_1212_U62, P3_ADD_371_1212_U63, P3_ADD_371_1212_U64, P3_ADD_371_1212_U65, P3_ADD_371_1212_U66, P3_ADD_371_1212_U67, P3_ADD_371_1212_U68, P3_ADD_371_1212_U69, P3_ADD_371_1212_U70, P3_ADD_371_1212_U71, P3_ADD_371_1212_U72, P3_ADD_371_1212_U73, P3_ADD_371_1212_U74, P3_ADD_371_1212_U75, P3_ADD_371_1212_U76, P3_ADD_371_1212_U77, P3_ADD_371_1212_U78, P3_ADD_371_1212_U79, P3_ADD_371_1212_U80, P3_ADD_371_1212_U81, P3_ADD_371_1212_U82, P3_ADD_371_1212_U83, P3_ADD_371_1212_U84, P3_ADD_371_1212_U85, P3_ADD_371_1212_U86, P3_ADD_371_1212_U87, P3_ADD_371_1212_U88, P3_ADD_371_1212_U89, P3_ADD_371_1212_U90, P3_ADD_371_1212_U91, P3_ADD_371_1212_U92, P3_ADD_371_1212_U93, P3_ADD_371_1212_U94, P3_ADD_371_1212_U95, P3_ADD_371_1212_U96, P3_ADD_371_1212_U97, P3_ADD_371_1212_U98, P3_ADD_371_1212_U99, P3_ADD_371_1212_U100, P3_ADD_371_1212_U101, P3_ADD_371_1212_U102, P3_ADD_371_1212_U103, P3_ADD_371_1212_U104, P3_ADD_371_1212_U105, P3_ADD_371_1212_U106, P3_ADD_371_1212_U107, P3_ADD_371_1212_U108, P3_ADD_371_1212_U109, P3_ADD_371_1212_U110, P3_ADD_371_1212_U111, P3_ADD_371_1212_U112, P3_ADD_371_1212_U113, P3_ADD_371_1212_U114, P3_ADD_371_1212_U115, P3_ADD_371_1212_U116, P3_ADD_371_1212_U117, P3_ADD_371_1212_U118, P3_ADD_371_1212_U119, P3_ADD_371_1212_U120, P3_ADD_371_1212_U121, P3_ADD_371_1212_U122, P3_ADD_371_1212_U123, P3_ADD_371_1212_U124, P3_ADD_371_1212_U125, P3_ADD_371_1212_U126, P3_ADD_371_1212_U127, P3_ADD_371_1212_U128, P3_ADD_371_1212_U129, P3_ADD_371_1212_U130, P3_ADD_371_1212_U131, P3_ADD_371_1212_U132, P3_ADD_371_1212_U133, P3_ADD_371_1212_U134, P3_ADD_371_1212_U135, P3_ADD_371_1212_U136, P3_ADD_371_1212_U137, P3_ADD_371_1212_U138, P3_ADD_371_1212_U139, P3_ADD_371_1212_U140, P3_ADD_371_1212_U141, P3_ADD_371_1212_U142, P3_ADD_371_1212_U143, P3_ADD_371_1212_U144, P3_ADD_371_1212_U145, P3_ADD_371_1212_U146, P3_ADD_371_1212_U147, P3_ADD_371_1212_U148, P3_ADD_371_1212_U149, P3_ADD_371_1212_U150, P3_ADD_371_1212_U151, P3_ADD_371_1212_U152, P3_ADD_371_1212_U153, P3_ADD_371_1212_U154, P3_ADD_371_1212_U155, P3_ADD_371_1212_U156, P3_ADD_371_1212_U157, P3_ADD_371_1212_U158, P3_ADD_371_1212_U159, P3_ADD_371_1212_U160, P3_ADD_371_1212_U161, P3_ADD_371_1212_U162, P3_ADD_371_1212_U163, P3_ADD_371_1212_U164, P3_ADD_371_1212_U165, P3_ADD_371_1212_U166, P3_ADD_371_1212_U167, P3_ADD_371_1212_U168, P3_ADD_371_1212_U169, P3_ADD_371_1212_U170, P3_ADD_371_1212_U171, P3_ADD_371_1212_U172, P3_ADD_371_1212_U173, P3_ADD_371_1212_U174, P3_ADD_371_1212_U175, P3_ADD_371_1212_U176, P3_ADD_371_1212_U177, P3_ADD_371_1212_U178, P3_ADD_371_1212_U179, P3_ADD_371_1212_U180, P3_ADD_371_1212_U181, P3_ADD_371_1212_U182, P3_ADD_371_1212_U183, P3_ADD_371_1212_U184, P3_ADD_371_1212_U185, P3_ADD_371_1212_U186, P3_ADD_371_1212_U187, P3_ADD_371_1212_U188, P3_ADD_371_1212_U189, P3_ADD_371_1212_U190, P3_ADD_371_1212_U191, P3_ADD_371_1212_U192, P3_ADD_371_1212_U193, P3_ADD_371_1212_U194, P3_ADD_371_1212_U195, P3_ADD_371_1212_U196, P3_ADD_371_1212_U197, P3_ADD_371_1212_U198, P3_ADD_371_1212_U199, P3_ADD_371_1212_U200, P3_ADD_371_1212_U201, P3_ADD_371_1212_U202, P3_ADD_371_1212_U203, P3_ADD_371_1212_U204, P3_ADD_371_1212_U205, P3_ADD_371_1212_U206, P3_ADD_371_1212_U207, P3_ADD_371_1212_U208, P3_ADD_371_1212_U209, P3_ADD_371_1212_U210, P3_ADD_371_1212_U211, P3_ADD_371_1212_U212, P3_ADD_371_1212_U213, P3_ADD_371_1212_U214, P3_ADD_371_1212_U215, P3_ADD_371_1212_U216, P3_ADD_371_1212_U217, P3_ADD_371_1212_U218, P3_ADD_371_1212_U219, P3_ADD_371_1212_U220, P3_ADD_371_1212_U221, P3_ADD_371_1212_U222, P3_ADD_371_1212_U223, P3_ADD_371_1212_U224, P3_ADD_371_1212_U225, P3_ADD_371_1212_U226, P3_ADD_371_1212_U227, P3_ADD_371_1212_U228, P3_ADD_371_1212_U229, P3_ADD_371_1212_U230, P3_ADD_371_1212_U231, P3_ADD_371_1212_U232, P3_ADD_371_1212_U233, P3_ADD_371_1212_U234, P3_ADD_371_1212_U235, P3_ADD_371_1212_U236, P3_ADD_371_1212_U237, P3_ADD_371_1212_U238, P3_ADD_371_1212_U239, P3_ADD_371_1212_U240, P3_ADD_371_1212_U241, P3_ADD_371_1212_U242, P3_ADD_371_1212_U243, P3_ADD_371_1212_U244, P3_ADD_371_1212_U245, P3_ADD_371_1212_U246, P3_ADD_371_1212_U247, P3_ADD_371_1212_U248, P3_ADD_371_1212_U249, P3_ADD_371_1212_U250, P3_ADD_371_1212_U251, P3_ADD_371_1212_U252, P3_ADD_371_1212_U253, P3_ADD_371_1212_U254, P3_ADD_371_1212_U255, P3_ADD_371_1212_U256, P3_ADD_371_1212_U257, P3_ADD_371_1212_U258, P3_ADD_371_1212_U259, P3_ADD_371_1212_U260, P3_ADD_371_1212_U261, P3_ADD_371_1212_U262, P3_ADD_371_1212_U263, P3_ADD_371_1212_U264, P3_ADD_371_1212_U265, P3_SUB_504_U6, P3_SUB_504_U7, P3_SUB_504_U8, P3_SUB_504_U9, P3_SUB_504_U10, P3_SUB_504_U11, P3_SUB_504_U12, P3_SUB_504_U13, P3_SUB_504_U14, P3_SUB_504_U15, P3_SUB_504_U16, P3_SUB_504_U17, P3_SUB_504_U18, P3_SUB_504_U19, P3_SUB_504_U20, P3_SUB_504_U21, P3_SUB_504_U22, P3_SUB_504_U23, P3_SUB_504_U24, P3_SUB_504_U25, P3_SUB_504_U26, P3_SUB_504_U27, P3_SUB_504_U28, P3_SUB_504_U29, P3_SUB_504_U30, P3_SUB_504_U31, P3_SUB_504_U32, P3_SUB_504_U33, P3_SUB_504_U34, P3_SUB_504_U35, P3_SUB_504_U36, P3_SUB_504_U37, P3_SUB_504_U38, P3_SUB_504_U39, P3_SUB_504_U40, P3_SUB_504_U41, P3_SUB_504_U42, P3_SUB_504_U43, P3_SUB_504_U44, P3_SUB_504_U45, P3_SUB_504_U46, P3_SUB_504_U47, P3_SUB_504_U48, P3_SUB_504_U49, P3_SUB_504_U50, P3_SUB_504_U51, P3_SUB_504_U52, P3_SUB_504_U53, P3_SUB_504_U54, P3_SUB_504_U55, P3_SUB_504_U56, P3_SUB_504_U57, P3_SUB_504_U58, P3_SUB_504_U59, P3_SUB_504_U60, P3_SUB_504_U61, P3_SUB_504_U62, P3_SUB_504_U63, P3_SUB_401_U6, P3_SUB_401_U7, P3_SUB_401_U8, P3_SUB_401_U9, P3_SUB_401_U10, P3_SUB_401_U11, P3_SUB_401_U12, P3_SUB_401_U13, P3_SUB_401_U14, P3_SUB_401_U15, P3_SUB_401_U16, P3_SUB_401_U17, P3_SUB_401_U18, P3_SUB_401_U19, P3_SUB_401_U20, P3_SUB_401_U21, P3_SUB_401_U22, P3_SUB_401_U23, P3_SUB_401_U24, P3_SUB_401_U25, P3_SUB_401_U26, P3_SUB_401_U27, P3_SUB_401_U28, P3_SUB_401_U29, P3_SUB_401_U30, P3_SUB_401_U31, P3_SUB_401_U32, P3_SUB_401_U33, P3_SUB_401_U34, P3_SUB_401_U35, P3_SUB_401_U36, P3_SUB_401_U37, P3_SUB_401_U38, P3_SUB_401_U39, P3_SUB_401_U40, P3_SUB_401_U41, P3_SUB_401_U42, P3_SUB_401_U43, P3_SUB_401_U44, P3_SUB_401_U45, P3_SUB_401_U46, P3_SUB_401_U47, P3_SUB_401_U48, P3_SUB_401_U49, P3_SUB_401_U50, P3_SUB_401_U51, P3_SUB_401_U52, P3_SUB_401_U53, P3_SUB_401_U54, P3_SUB_401_U55, P3_SUB_401_U56, P3_SUB_401_U57, P3_SUB_401_U58, P3_SUB_401_U59, P3_SUB_401_U60, P3_SUB_401_U61, P3_SUB_401_U62, P3_SUB_401_U63, P3_SUB_401_U64, P3_SUB_401_U65, P3_SUB_401_U66, P3_ADD_371_U4, P3_ADD_371_U5, P3_ADD_371_U6, P3_ADD_371_U7, P3_ADD_371_U8, P3_ADD_371_U9, P3_ADD_371_U10, P3_ADD_371_U11, P3_ADD_371_U12, P3_ADD_371_U13, P3_ADD_371_U14, P3_ADD_371_U15, P3_ADD_371_U16, P3_ADD_371_U17, P3_ADD_371_U18, P3_ADD_371_U19, P3_ADD_371_U20, P3_ADD_371_U21, P3_ADD_371_U22, P3_ADD_371_U23, P3_ADD_371_U24, P3_ADD_371_U25, P3_ADD_371_U26, P3_ADD_371_U27, P3_ADD_371_U28, P3_ADD_371_U29, P3_ADD_371_U30, P3_ADD_371_U31, P3_ADD_371_U32, P3_ADD_371_U33, P3_ADD_371_U34, P3_ADD_371_U35, P3_ADD_371_U36, P3_ADD_371_U37, P3_ADD_371_U38, P3_ADD_371_U39, P3_ADD_371_U40, P3_ADD_371_U41, P3_ADD_371_U42, P3_ADD_371_U43, P3_ADD_371_U44, P3_SUB_390_U6, P3_SUB_390_U7, P3_SUB_390_U8, P3_SUB_390_U9, P3_SUB_390_U10, P3_SUB_390_U11, P3_SUB_390_U12, P3_SUB_390_U13, P3_SUB_390_U14, P3_SUB_390_U15, P3_SUB_390_U16, P3_SUB_390_U17, P3_SUB_390_U18, P3_SUB_390_U19, P3_SUB_390_U20, P3_SUB_390_U21, P3_SUB_390_U22, P3_SUB_390_U23, P3_SUB_390_U24, P3_SUB_390_U25, P3_SUB_390_U26, P3_SUB_390_U27, P3_SUB_390_U28, P3_SUB_390_U29, P3_SUB_390_U30, P3_SUB_390_U31, P3_SUB_390_U32, P3_SUB_390_U33, P3_SUB_390_U34, P3_SUB_390_U35, P3_SUB_390_U36, P3_SUB_390_U37, P3_SUB_390_U38, P3_SUB_390_U39, P3_SUB_390_U40, P3_SUB_390_U41, P3_SUB_390_U42, P3_SUB_390_U43, P3_SUB_390_U44, P3_SUB_390_U45, P3_SUB_390_U46, P3_SUB_390_U47, P3_SUB_390_U48, P3_SUB_390_U49, P3_SUB_390_U50, P3_SUB_390_U51, P3_SUB_390_U52, P3_SUB_390_U53, P3_SUB_390_U54, P3_SUB_390_U55, P3_SUB_390_U56, P3_SUB_390_U57, P3_SUB_390_U58, P3_SUB_390_U59, P3_SUB_390_U60, P3_SUB_390_U61, P3_SUB_390_U62, P3_SUB_390_U63, P3_SUB_390_U64, P3_SUB_390_U65, P3_SUB_390_U66, P3_SUB_357_U6, P3_SUB_357_U7, P3_SUB_357_U8, P3_SUB_357_U9, P3_SUB_357_U10, P3_SUB_357_U11, P3_SUB_357_U12, P3_SUB_357_U13, P3_ADD_495_U4, P3_ADD_495_U5, P3_ADD_495_U6, P3_ADD_495_U7, P3_ADD_495_U8, P3_ADD_495_U9, P3_ADD_495_U10, P3_ADD_495_U11, P3_ADD_495_U12, P3_ADD_495_U13, P3_ADD_495_U14, P3_ADD_495_U15, P3_ADD_495_U16, P3_ADD_495_U17, P3_ADD_495_U18, P3_ADD_495_U19, P3_ADD_495_U20, P3_GTE_412_U6, P3_GTE_412_U7, P3_GTE_504_U6, P3_GTE_504_U7, P3_ADD_494_U4, P3_ADD_494_U5, P3_ADD_494_U6, P3_ADD_494_U7, P3_ADD_494_U8, P3_ADD_494_U9, P3_ADD_494_U10, P3_ADD_494_U11, P3_ADD_494_U12, P3_ADD_494_U13, P3_ADD_494_U14, P3_ADD_494_U15, P3_ADD_494_U16, P3_ADD_494_U17, P3_ADD_494_U18, P3_ADD_494_U19, P3_ADD_494_U20, P3_ADD_494_U21, P3_ADD_494_U22, P3_ADD_494_U23, P3_ADD_494_U24, P3_ADD_494_U25, P3_ADD_494_U26, P3_ADD_494_U27, P3_ADD_494_U28, P3_ADD_494_U29, P3_ADD_494_U30, P3_ADD_494_U31, P3_ADD_494_U32, P3_ADD_494_U33, P3_ADD_494_U34, P3_ADD_494_U35, P3_ADD_494_U36, P3_ADD_494_U37, P3_ADD_494_U38, P3_ADD_494_U39, P3_ADD_494_U40, P3_ADD_494_U41, P3_ADD_494_U42, P3_ADD_494_U43, P3_ADD_494_U44, P3_ADD_494_U45, P3_ADD_494_U46, P3_ADD_494_U47, P3_ADD_494_U48, P3_ADD_494_U49, P3_ADD_494_U50, P3_ADD_494_U51, P3_ADD_494_U52, P3_ADD_494_U53, P3_ADD_494_U54, P3_ADD_494_U55, P3_ADD_494_U56, P3_ADD_494_U57, P3_ADD_494_U58, P3_ADD_494_U59, P3_ADD_494_U60, P3_ADD_494_U61, P3_ADD_494_U62, P3_ADD_494_U63, P3_ADD_494_U64, P3_ADD_494_U65, P3_ADD_494_U66, P3_ADD_494_U67, P3_ADD_494_U68, P3_ADD_494_U69, P3_ADD_494_U70, P3_ADD_494_U71, P3_ADD_494_U72, P3_ADD_494_U73, P3_ADD_494_U74, P3_ADD_494_U75, P3_ADD_494_U76, P3_ADD_494_U77, P3_ADD_494_U78, P3_ADD_494_U79, P3_ADD_494_U80, P3_ADD_494_U81, P3_ADD_494_U82, P3_ADD_494_U83, P3_ADD_494_U84, P3_ADD_494_U85, P3_ADD_494_U86, P3_ADD_494_U87, P3_ADD_494_U88, P3_ADD_494_U89, P3_ADD_494_U90, P3_ADD_494_U91, P3_ADD_494_U92, P3_ADD_494_U93, P3_ADD_494_U94, P3_ADD_494_U95, P3_ADD_494_U96, P3_ADD_494_U97, P3_ADD_494_U98, P3_ADD_494_U99, P3_ADD_494_U100, P3_ADD_494_U101, P3_ADD_494_U102, P3_ADD_494_U103, P3_ADD_494_U104, P3_ADD_494_U105, P3_ADD_494_U106, P3_ADD_494_U107, P3_ADD_494_U108, P3_ADD_494_U109, P3_ADD_494_U110, P3_ADD_494_U111, P3_ADD_494_U112, P3_ADD_494_U113, P3_ADD_494_U114, P3_ADD_494_U115, P3_ADD_494_U116, P3_ADD_494_U117, P3_ADD_494_U118, P3_ADD_494_U119, P3_ADD_494_U120, P3_ADD_494_U121, P3_ADD_494_U122, P3_ADD_494_U123, P3_ADD_494_U124, P3_ADD_494_U125, P3_ADD_494_U126, P3_ADD_494_U127, P3_ADD_494_U128, P3_ADD_494_U129, P3_ADD_494_U130, P3_ADD_494_U131, P3_ADD_494_U132, P3_ADD_494_U133, P3_ADD_494_U134, P3_ADD_494_U135, P3_ADD_494_U136, P3_ADD_494_U137, P3_ADD_494_U138, P3_ADD_494_U139, P3_ADD_494_U140, P3_ADD_494_U141, P3_ADD_494_U142, P3_ADD_494_U143, P3_ADD_494_U144, P3_ADD_494_U145, P3_ADD_494_U146, P3_ADD_494_U147, P3_ADD_494_U148, P3_ADD_494_U149, P3_ADD_494_U150, P3_ADD_494_U151, P3_ADD_494_U152, P3_ADD_494_U153, P3_ADD_494_U154, P3_ADD_494_U155, P3_ADD_494_U156, P3_ADD_494_U157, P3_ADD_494_U158, P3_ADD_494_U159, P3_ADD_494_U160, P3_ADD_494_U161, P3_ADD_494_U162, P3_ADD_494_U163, P3_ADD_494_U164, P3_ADD_494_U165, P3_ADD_494_U166, P3_ADD_494_U167, P3_ADD_494_U168, P3_ADD_494_U169, P3_ADD_494_U170, P3_ADD_494_U171, P3_ADD_494_U172, P3_ADD_494_U173, P3_ADD_494_U174, P3_ADD_494_U175, P3_ADD_494_U176, P3_ADD_494_U177, P3_ADD_494_U178, P3_ADD_494_U179, P3_ADD_494_U180, P3_ADD_494_U181, P3_ADD_494_U182, P3_ADD_536_U4, P3_ADD_536_U5, P3_ADD_536_U6, P3_ADD_536_U7, P3_ADD_536_U8, P3_ADD_536_U9, P3_ADD_536_U10, P3_ADD_536_U11, P3_ADD_536_U12, P3_ADD_536_U13, P3_ADD_536_U14, P3_ADD_536_U15, P3_ADD_536_U16, P3_ADD_536_U17, P3_ADD_536_U18, P3_ADD_536_U19, P3_ADD_536_U20, P3_ADD_536_U21, P3_ADD_536_U22, P3_ADD_536_U23, P3_ADD_536_U24, P3_ADD_536_U25, P3_ADD_536_U26, P3_ADD_536_U27, P3_ADD_536_U28, P3_ADD_536_U29, P3_ADD_536_U30, P3_ADD_536_U31, P3_ADD_536_U32, P3_ADD_536_U33, P3_ADD_536_U34, P3_ADD_536_U35, P3_ADD_536_U36, P3_ADD_536_U37, P3_ADD_536_U38, P3_ADD_536_U39, P3_ADD_536_U40, P3_ADD_536_U41, P3_ADD_536_U42, P3_ADD_536_U43, P3_ADD_536_U44, P3_ADD_536_U45, P3_ADD_536_U46, P3_ADD_536_U47, P3_ADD_536_U48, P3_ADD_536_U49, P3_ADD_536_U50, P3_ADD_536_U51, P3_ADD_536_U52, P3_ADD_536_U53, P3_ADD_536_U54, P3_ADD_536_U55, P3_ADD_536_U56, P3_ADD_536_U57, P3_ADD_536_U58, P3_ADD_536_U59, P3_ADD_536_U60, P3_ADD_536_U61, P3_ADD_536_U62, P3_ADD_536_U63, P3_ADD_536_U64, P3_ADD_536_U65, P3_ADD_536_U66, P3_ADD_536_U67, P3_ADD_536_U68, P3_ADD_536_U69, P3_ADD_536_U70, P3_ADD_536_U71, P3_ADD_536_U72, P3_ADD_536_U73, P3_ADD_536_U74, P3_ADD_536_U75, P3_ADD_536_U76, P3_ADD_536_U77, P3_ADD_536_U78, P3_ADD_536_U79, P3_ADD_536_U80, P3_ADD_536_U81, P3_ADD_536_U82, P3_ADD_536_U83, P3_ADD_536_U84, P3_ADD_536_U85, P3_ADD_536_U86, P3_ADD_536_U87, P3_ADD_536_U88, P3_ADD_536_U89, P3_ADD_536_U90, P3_ADD_536_U91, P3_ADD_536_U92, P3_ADD_536_U93, P3_ADD_536_U94, P3_ADD_536_U95, P3_ADD_536_U96, P3_ADD_536_U97, P3_ADD_536_U98, P3_ADD_536_U99, P3_ADD_536_U100, P3_ADD_536_U101, P3_ADD_536_U102, P3_ADD_536_U103, P3_ADD_536_U104, P3_ADD_536_U105, P3_ADD_536_U106, P3_ADD_536_U107, P3_ADD_536_U108, P3_ADD_536_U109, P3_ADD_536_U110, P3_ADD_536_U111, P3_ADD_536_U112, P3_ADD_536_U113, P3_ADD_536_U114, P3_ADD_536_U115, P3_ADD_536_U116, P3_ADD_536_U117, P3_ADD_536_U118, P3_ADD_536_U119, P3_ADD_536_U120, P3_ADD_536_U121, P3_ADD_536_U122, P3_ADD_536_U123, P3_ADD_536_U124, P3_ADD_536_U125, P3_ADD_536_U126, P3_ADD_536_U127, P3_ADD_536_U128, P3_ADD_536_U129, P3_ADD_536_U130, P3_ADD_536_U131, P3_ADD_536_U132, P3_ADD_536_U133, P3_ADD_536_U134, P3_ADD_536_U135, P3_ADD_536_U136, P3_ADD_536_U137, P3_ADD_536_U138, P3_ADD_536_U139, P3_ADD_536_U140, P3_ADD_536_U141, P3_ADD_536_U142, P3_ADD_536_U143, P3_ADD_536_U144, P3_ADD_536_U145, P3_ADD_536_U146, P3_ADD_536_U147, P3_ADD_536_U148, P3_ADD_536_U149, P3_ADD_536_U150, P3_ADD_536_U151, P3_ADD_536_U152, P3_ADD_536_U153, P3_ADD_536_U154, P3_ADD_536_U155, P3_ADD_536_U156, P3_ADD_536_U157, P3_ADD_536_U158, P3_ADD_536_U159, P3_ADD_536_U160, P3_ADD_536_U161, P3_ADD_536_U162, P3_ADD_536_U163, P3_ADD_536_U164, P3_ADD_536_U165, P3_ADD_536_U166, P3_ADD_536_U167, P3_ADD_536_U168, P3_ADD_536_U169, P3_ADD_536_U170, P3_ADD_536_U171, P3_ADD_536_U172, P3_ADD_536_U173, P3_ADD_536_U174, P3_ADD_536_U175, P3_ADD_536_U176, P3_ADD_536_U177, P3_ADD_536_U178, P3_ADD_536_U179, P3_ADD_536_U180, P3_ADD_536_U181, P3_ADD_536_U182, P3_ADD_402_1132_U4, P3_ADD_402_1132_U5, P3_ADD_402_1132_U6, P3_ADD_402_1132_U7, P3_ADD_402_1132_U8, P3_ADD_402_1132_U9, P3_ADD_402_1132_U10, P3_ADD_402_1132_U11, P3_ADD_402_1132_U12, P3_ADD_402_1132_U13, P3_ADD_402_1132_U14, P3_ADD_402_1132_U15, P3_ADD_402_1132_U16, P3_ADD_402_1132_U17, P3_ADD_402_1132_U18, P3_ADD_402_1132_U19, P3_ADD_402_1132_U20, P3_ADD_402_1132_U21, P3_ADD_402_1132_U22, P3_ADD_402_1132_U23, P3_ADD_402_1132_U24, P3_ADD_402_1132_U25, P3_ADD_402_1132_U26, P3_ADD_402_1132_U27, P3_ADD_402_1132_U28, P3_ADD_402_1132_U29, P3_ADD_402_1132_U30, P3_ADD_402_1132_U31, P3_ADD_402_1132_U32, P3_ADD_402_1132_U33, P3_ADD_402_1132_U34, P3_ADD_402_1132_U35, P3_ADD_402_1132_U36, P3_ADD_402_1132_U37, P3_ADD_402_1132_U38, P3_ADD_402_1132_U39, P3_ADD_402_1132_U40, P3_ADD_402_1132_U41, P3_ADD_402_1132_U42, P3_ADD_402_1132_U43, P3_ADD_402_1132_U44, P3_ADD_402_1132_U45, P3_ADD_402_1132_U46, P3_ADD_402_1132_U47, P3_ADD_402_1132_U48, P3_ADD_402_1132_U49, P3_ADD_402_1132_U50, P2_R2099_U5, P2_R2099_U6, P2_R2099_U7, P2_R2099_U8, P2_R2099_U9, P2_R2099_U10, P2_R2099_U11, P2_R2099_U12, P2_R2099_U13, P2_R2099_U14, P2_R2099_U15, P2_R2099_U16, P2_R2099_U17, P2_R2099_U18, P2_R2099_U19, P2_R2099_U20, P2_R2099_U21, P2_R2099_U22, P2_R2099_U23, P2_R2099_U24, P2_R2099_U25, P2_R2099_U26, P2_R2099_U27, P2_R2099_U28, P2_R2099_U29, P2_R2099_U30, P2_R2099_U31, P2_R2099_U32, P2_R2099_U33, P2_R2099_U34, P2_R2099_U35, P2_R2099_U36, P2_R2099_U37, P2_R2099_U38, P2_R2099_U39, P2_R2099_U40, P2_R2099_U41, P2_R2099_U42, P2_R2099_U43, P2_R2099_U44, P2_R2099_U45, P2_R2099_U46, P2_R2099_U47, P2_R2099_U48, P2_R2099_U49, P2_R2099_U50, P2_R2099_U51, P2_R2099_U52, P2_R2099_U53, P2_R2099_U54, P2_R2099_U55, P2_R2099_U56, P2_R2099_U57, P2_R2099_U58, P2_R2099_U59, P2_R2099_U60, P2_R2099_U61, P2_R2099_U62, P2_R2099_U63, P2_R2099_U64, P2_R2099_U65, P2_R2099_U66, P2_R2099_U67, P2_R2099_U68, P2_R2099_U69, P2_R2099_U70, P2_R2099_U71, P2_R2099_U72, P2_R2099_U73, P2_R2099_U74, P2_R2099_U75, P2_R2099_U76, P2_R2099_U77, P2_R2099_U78, P2_R2099_U79, P2_R2099_U80, P2_R2099_U81, P2_R2099_U82, P2_R2099_U83, P2_R2099_U84, P2_R2099_U85, P2_R2099_U86, P2_R2099_U87, P2_R2099_U88, P2_R2099_U89, P2_R2099_U90, P2_R2099_U91, P2_R2099_U92, P2_R2099_U93, P2_R2099_U94, P2_R2099_U95, P2_R2099_U96, P2_R2099_U97, P2_R2099_U98, P2_R2099_U99, P2_R2099_U100, P2_R2099_U101, P2_R2099_U102, P2_R2099_U103, P2_R2099_U104, P2_R2099_U105, P2_R2099_U106, P2_R2099_U107, P2_R2099_U108, P2_R2099_U109, P2_R2099_U110, P2_R2099_U111, P2_R2099_U112, P2_R2099_U113, P2_R2099_U114, P2_R2099_U115, P2_R2099_U116, P2_R2099_U117, P2_R2099_U118, P2_R2099_U119, P2_R2099_U120, P2_R2099_U121, P2_R2099_U122, P2_R2099_U123, P2_R2099_U124, P2_R2099_U125, P2_R2099_U126, P2_R2099_U127, P2_R2099_U128, P2_R2099_U129, P2_R2099_U130, P2_R2099_U131, P2_R2099_U132, P2_R2099_U133, P2_R2099_U134, P2_R2099_U135, P2_R2099_U136, P2_R2099_U137, P2_R2099_U138, P2_R2099_U139, P2_R2099_U140, P2_R2099_U141, P2_R2099_U142, P2_R2099_U143, P2_R2099_U144, P2_R2099_U145, P2_R2099_U146, P2_R2099_U147, P2_R2099_U148, P2_R2099_U149, P2_R2099_U150, P2_R2099_U151, P2_R2099_U152, P2_R2099_U153, P2_R2099_U154, P2_R2099_U155, P2_R2099_U156, P2_R2099_U157, P2_R2099_U158, P2_R2099_U159, P2_R2099_U160, P2_R2099_U161, P2_R2099_U162, P2_R2099_U163, P2_R2099_U164, P2_R2099_U165, P2_R2099_U166, P2_R2099_U167, P2_R2099_U168, P2_R2099_U169, P2_R2099_U170, P2_R2099_U171, P2_R2099_U172, P2_R2099_U173, P2_R2099_U174, P2_R2099_U175, P2_R2099_U176, P2_R2099_U177, P2_R2099_U178, P2_R2099_U179, P2_R2099_U180, P2_R2099_U181, P2_R2099_U182, P2_R2099_U183, P2_R2099_U184, P2_R2099_U185, P2_R2099_U186, P2_R2099_U187, P2_R2099_U188, P2_R2099_U189, P2_R2099_U190, P2_R2099_U191, P2_R2099_U192, P2_R2099_U193, P2_R2099_U194, P2_R2099_U195, P2_R2099_U196, P2_R2099_U197, P2_R2099_U198, P2_R2099_U199, P2_R2099_U200, P2_R2099_U201, P2_R2099_U202, P2_R2099_U203, P2_R2099_U204, P2_R2099_U205, P2_R2099_U206, P2_R2099_U207, P2_R2099_U208, P2_R2099_U209, P2_R2099_U210, P2_R2099_U211, P2_R2099_U212, P2_R2099_U213, P2_R2099_U214, P2_R2099_U215, P2_R2099_U216, P2_R2099_U217, P2_R2099_U218, P2_R2099_U219, P2_R2099_U220, P2_R2099_U221, P2_R2099_U222, P2_R2099_U223, P2_R2099_U224, P2_R2099_U225, P2_ADD_391_1196_U5, P2_ADD_391_1196_U6, P2_ADD_391_1196_U7, P2_ADD_391_1196_U8, P2_ADD_391_1196_U9, P2_ADD_391_1196_U10, P2_ADD_391_1196_U11, P2_ADD_391_1196_U12, P2_ADD_391_1196_U13, P2_ADD_391_1196_U14, P2_ADD_391_1196_U15, P2_ADD_391_1196_U16, P2_ADD_391_1196_U17, P2_ADD_391_1196_U18, P2_ADD_391_1196_U19, P2_ADD_391_1196_U20, P2_ADD_391_1196_U21, P2_ADD_391_1196_U22, P2_ADD_391_1196_U23, P2_ADD_391_1196_U24, P2_ADD_391_1196_U25, P2_ADD_391_1196_U26, P2_ADD_391_1196_U27, P2_ADD_391_1196_U28, P2_ADD_391_1196_U29, P2_ADD_391_1196_U30, P2_ADD_391_1196_U31, P2_ADD_391_1196_U32, P2_ADD_391_1196_U33, P2_ADD_391_1196_U34, P2_ADD_391_1196_U35, P2_ADD_391_1196_U36, P2_ADD_391_1196_U37, P2_ADD_391_1196_U38, P2_ADD_391_1196_U39, P2_ADD_391_1196_U40, P2_ADD_391_1196_U41, P2_ADD_391_1196_U42, P2_ADD_391_1196_U43, P2_ADD_391_1196_U44, P2_ADD_391_1196_U45, P2_ADD_391_1196_U46, P2_ADD_391_1196_U47, P2_ADD_391_1196_U48, P2_ADD_391_1196_U49, P2_ADD_391_1196_U50, P2_ADD_391_1196_U51, P2_ADD_391_1196_U52, P2_ADD_391_1196_U53, P2_ADD_391_1196_U54, P2_ADD_391_1196_U55, P2_ADD_391_1196_U56, P2_ADD_391_1196_U57, P2_ADD_391_1196_U58, P2_ADD_391_1196_U59, P2_ADD_391_1196_U60, P2_ADD_391_1196_U61, P2_ADD_391_1196_U62, P2_ADD_391_1196_U63, P2_ADD_391_1196_U64, P2_ADD_391_1196_U65, P2_ADD_391_1196_U66, P2_ADD_391_1196_U67, P2_ADD_391_1196_U68, P2_ADD_391_1196_U69, P2_ADD_391_1196_U70, P2_ADD_391_1196_U71, P2_ADD_391_1196_U72, P2_ADD_391_1196_U73, P2_ADD_391_1196_U74, P2_ADD_391_1196_U75, P2_ADD_391_1196_U76, P2_ADD_391_1196_U77, P2_ADD_391_1196_U78, P2_ADD_391_1196_U79, P2_ADD_391_1196_U80, P2_ADD_391_1196_U81, P2_ADD_391_1196_U82, P2_ADD_391_1196_U83, P2_ADD_391_1196_U84, P2_ADD_391_1196_U85, P2_ADD_391_1196_U86, P2_ADD_391_1196_U87, P2_ADD_391_1196_U88, P2_ADD_391_1196_U89, P2_ADD_391_1196_U90, P2_ADD_391_1196_U91, P2_ADD_391_1196_U92, P2_ADD_391_1196_U93, P2_ADD_391_1196_U94, P2_ADD_391_1196_U95, P2_ADD_391_1196_U96, P2_ADD_391_1196_U97, P2_ADD_391_1196_U98, P2_ADD_391_1196_U99, P2_ADD_391_1196_U100, P2_ADD_391_1196_U101, P2_ADD_391_1196_U102, P2_ADD_391_1196_U103, P2_ADD_391_1196_U104, P2_ADD_391_1196_U105, P2_ADD_391_1196_U106, P2_ADD_391_1196_U107, P2_ADD_391_1196_U108, P2_ADD_391_1196_U109, P2_ADD_391_1196_U110, P2_ADD_391_1196_U111, P2_ADD_391_1196_U112, P2_ADD_391_1196_U113, P2_ADD_391_1196_U114, P2_ADD_391_1196_U115, P2_ADD_391_1196_U116, P2_ADD_391_1196_U117, P2_ADD_391_1196_U118, P2_ADD_391_1196_U119, P2_ADD_391_1196_U120, P2_ADD_391_1196_U121, P2_ADD_391_1196_U122, P2_ADD_391_1196_U123, P2_ADD_391_1196_U124, P2_ADD_391_1196_U125, P2_ADD_391_1196_U126, P2_ADD_391_1196_U127, P2_ADD_391_1196_U128, P2_ADD_391_1196_U129, P2_ADD_391_1196_U130, P2_ADD_391_1196_U131, P2_ADD_391_1196_U132, P2_ADD_391_1196_U133, P2_ADD_391_1196_U134, P2_ADD_391_1196_U135, P2_ADD_391_1196_U136, P2_ADD_391_1196_U137, P2_ADD_391_1196_U138, P2_ADD_391_1196_U139, P2_ADD_391_1196_U140, P2_ADD_391_1196_U141, P2_ADD_391_1196_U142, P2_ADD_391_1196_U143, P2_ADD_391_1196_U144, P2_ADD_391_1196_U145, P2_ADD_391_1196_U146, P2_ADD_391_1196_U147, P2_ADD_391_1196_U148, P2_ADD_391_1196_U149, P2_ADD_391_1196_U150, P2_ADD_391_1196_U151, P2_ADD_391_1196_U152, P2_ADD_391_1196_U153, P2_ADD_391_1196_U154, P2_ADD_391_1196_U155, P2_ADD_391_1196_U156, P2_ADD_391_1196_U157, P2_ADD_391_1196_U158, P2_ADD_391_1196_U159, P2_ADD_391_1196_U160, P2_ADD_391_1196_U161, P2_ADD_391_1196_U162, P2_ADD_391_1196_U163, P2_ADD_391_1196_U164, P2_ADD_391_1196_U165, P2_ADD_391_1196_U166, P2_ADD_391_1196_U167, P2_ADD_391_1196_U168, P2_ADD_391_1196_U169, P2_ADD_391_1196_U170, P2_ADD_391_1196_U171, P2_ADD_391_1196_U172, P2_ADD_391_1196_U173, P2_ADD_391_1196_U174, P2_ADD_391_1196_U175, P2_ADD_391_1196_U176, P2_ADD_391_1196_U177, P2_ADD_391_1196_U178, P2_ADD_391_1196_U179, P2_ADD_391_1196_U180, P2_ADD_391_1196_U181, P2_ADD_391_1196_U182, P2_ADD_391_1196_U183, P2_ADD_391_1196_U184, P2_ADD_391_1196_U185, P2_ADD_391_1196_U186, P2_ADD_391_1196_U187, P2_ADD_391_1196_U188, P2_ADD_391_1196_U189, P2_ADD_391_1196_U190, P2_ADD_391_1196_U191, P2_ADD_391_1196_U192, P2_ADD_391_1196_U193, P2_ADD_391_1196_U194, P2_ADD_391_1196_U195, P2_ADD_391_1196_U196, P2_ADD_391_1196_U197, P2_ADD_391_1196_U198, P2_ADD_391_1196_U199, P2_ADD_391_1196_U200, P2_ADD_391_1196_U201, P2_ADD_391_1196_U202, P2_ADD_391_1196_U203, P2_ADD_391_1196_U204, P2_ADD_391_1196_U205, P2_ADD_391_1196_U206, P2_ADD_391_1196_U207, P2_ADD_391_1196_U208, P2_ADD_391_1196_U209, P2_ADD_391_1196_U210, P2_ADD_391_1196_U211, P2_ADD_391_1196_U212, P2_ADD_391_1196_U213, P2_ADD_391_1196_U214, P2_ADD_391_1196_U215, P2_ADD_391_1196_U216, P2_ADD_391_1196_U217, P2_ADD_391_1196_U218, P2_ADD_391_1196_U219, P2_ADD_391_1196_U220, P2_ADD_391_1196_U221, P2_ADD_391_1196_U222, P2_ADD_391_1196_U223, P2_ADD_391_1196_U224, P2_ADD_391_1196_U225, P2_ADD_391_1196_U226, P2_ADD_391_1196_U227, P2_ADD_391_1196_U228, P2_ADD_391_1196_U229, P2_ADD_391_1196_U230, P2_ADD_391_1196_U231, P2_ADD_391_1196_U232, P2_ADD_391_1196_U233, P2_ADD_391_1196_U234, P2_ADD_391_1196_U235, P2_ADD_391_1196_U236, P2_ADD_391_1196_U237, P2_ADD_391_1196_U238, P2_ADD_391_1196_U239, P2_ADD_391_1196_U240, P2_ADD_391_1196_U241, P2_ADD_391_1196_U242, P2_ADD_391_1196_U243, P2_ADD_391_1196_U244, P2_ADD_391_1196_U245, P2_ADD_391_1196_U246, P2_ADD_391_1196_U247, P2_ADD_391_1196_U248, P2_ADD_391_1196_U249, P2_ADD_391_1196_U250, P2_ADD_391_1196_U251, P2_ADD_391_1196_U252, P2_ADD_391_1196_U253, P2_ADD_391_1196_U254, P2_ADD_391_1196_U255, P2_ADD_391_1196_U256, P2_ADD_391_1196_U257, P2_ADD_391_1196_U258, P2_ADD_391_1196_U259, P2_ADD_391_1196_U260, P2_ADD_391_1196_U261, P2_ADD_391_1196_U262, P2_ADD_391_1196_U263, P2_ADD_391_1196_U264, P2_ADD_391_1196_U265, P2_ADD_391_1196_U266, P2_ADD_391_1196_U267, P2_ADD_391_1196_U268, P2_ADD_391_1196_U269, P2_ADD_391_1196_U270, P2_ADD_391_1196_U271, P2_ADD_391_1196_U272, P2_ADD_391_1196_U273, P2_ADD_391_1196_U274, P2_ADD_391_1196_U275, P2_ADD_391_1196_U276, P2_ADD_391_1196_U277, P2_ADD_391_1196_U278, P2_ADD_391_1196_U279, P2_ADD_391_1196_U280, P2_ADD_391_1196_U281, P2_ADD_391_1196_U282, P2_ADD_391_1196_U283, P2_ADD_391_1196_U284, P2_ADD_391_1196_U285, P2_ADD_391_1196_U286, P2_ADD_391_1196_U287, P2_ADD_391_1196_U288, P2_ADD_391_1196_U289, P2_ADD_391_1196_U290, P2_ADD_391_1196_U291, P2_ADD_391_1196_U292, P2_ADD_391_1196_U293, P2_ADD_391_1196_U294, P2_ADD_391_1196_U295, P2_ADD_391_1196_U296, P2_ADD_391_1196_U297, P2_ADD_391_1196_U298, P2_ADD_391_1196_U299, P2_ADD_391_1196_U300, P2_ADD_391_1196_U301, P2_ADD_391_1196_U302, P2_ADD_391_1196_U303, P2_ADD_391_1196_U304, P2_ADD_391_1196_U305, P2_ADD_391_1196_U306, P2_ADD_391_1196_U307, P2_ADD_391_1196_U308, P2_ADD_391_1196_U309, P2_ADD_391_1196_U310, P2_ADD_391_1196_U311, P2_ADD_391_1196_U312, P2_ADD_391_1196_U313, P2_ADD_391_1196_U314, P2_ADD_391_1196_U315, P2_ADD_391_1196_U316, P2_ADD_391_1196_U317, P2_ADD_391_1196_U318, P2_ADD_391_1196_U319, P2_ADD_391_1196_U320, P2_ADD_391_1196_U321, P2_ADD_391_1196_U322, P2_ADD_391_1196_U323, P2_ADD_391_1196_U324, P2_ADD_391_1196_U325, P2_ADD_391_1196_U326, P2_ADD_391_1196_U327, P2_ADD_391_1196_U328, P2_ADD_391_1196_U329, P2_ADD_391_1196_U330, P2_ADD_391_1196_U331, P2_ADD_391_1196_U332, P2_ADD_391_1196_U333, P2_ADD_391_1196_U334, P2_ADD_391_1196_U335, P2_ADD_391_1196_U336, P2_ADD_391_1196_U337, P2_ADD_391_1196_U338, P2_ADD_391_1196_U339, P2_ADD_391_1196_U340, P2_ADD_391_1196_U341, P2_ADD_391_1196_U342, P2_ADD_391_1196_U343, P2_ADD_391_1196_U344, P2_ADD_391_1196_U345, P2_ADD_391_1196_U346, P2_ADD_391_1196_U347, P2_ADD_391_1196_U348, P2_ADD_391_1196_U349, P2_ADD_391_1196_U350, P2_ADD_391_1196_U351, P2_ADD_391_1196_U352, P2_ADD_391_1196_U353, P2_ADD_391_1196_U354, P2_ADD_391_1196_U355, P2_ADD_391_1196_U356, P2_ADD_391_1196_U357, P2_ADD_391_1196_U358, P2_ADD_391_1196_U359, P2_ADD_391_1196_U360, P2_ADD_391_1196_U361, P2_ADD_391_1196_U362, P2_ADD_391_1196_U363, P2_ADD_391_1196_U364, P2_ADD_391_1196_U365, P2_ADD_391_1196_U366, P2_ADD_391_1196_U367, P2_ADD_391_1196_U368, P2_ADD_391_1196_U369, P2_ADD_391_1196_U370, P2_ADD_391_1196_U371, P2_ADD_391_1196_U372, P2_ADD_391_1196_U373, P2_ADD_391_1196_U374, P2_ADD_391_1196_U375, P2_ADD_391_1196_U376, P2_ADD_391_1196_U377, P2_ADD_391_1196_U378, P2_ADD_391_1196_U379, P2_ADD_391_1196_U380, P2_ADD_391_1196_U381, P2_ADD_391_1196_U382, P2_ADD_391_1196_U383, P2_ADD_391_1196_U384, P2_ADD_391_1196_U385, P2_ADD_391_1196_U386, P2_ADD_391_1196_U387, P2_ADD_391_1196_U388, P2_ADD_391_1196_U389, P2_ADD_391_1196_U390, P2_ADD_391_1196_U391, P2_ADD_391_1196_U392, P2_ADD_391_1196_U393, P2_ADD_391_1196_U394, P2_ADD_391_1196_U395, P2_ADD_391_1196_U396, P2_ADD_391_1196_U397, P2_ADD_391_1196_U398, P2_ADD_391_1196_U399, P2_ADD_391_1196_U400, P2_ADD_391_1196_U401, P2_ADD_391_1196_U402, P2_ADD_391_1196_U403, P2_ADD_391_1196_U404, P2_ADD_391_1196_U405, P2_ADD_391_1196_U406, P2_ADD_391_1196_U407, P2_ADD_391_1196_U408, P2_ADD_391_1196_U409, P2_ADD_391_1196_U410, P2_ADD_391_1196_U411, P2_ADD_391_1196_U412, P2_ADD_391_1196_U413, P2_ADD_391_1196_U414, P2_ADD_391_1196_U415, P2_ADD_391_1196_U416, P2_ADD_391_1196_U417, P2_ADD_391_1196_U418, P2_ADD_391_1196_U419, P2_ADD_391_1196_U420, P2_ADD_391_1196_U421, P2_ADD_391_1196_U422, P2_ADD_391_1196_U423, P2_ADD_391_1196_U424, P2_ADD_391_1196_U425, P2_ADD_391_1196_U426, P2_ADD_391_1196_U427, P2_ADD_391_1196_U428, P2_ADD_391_1196_U429, P2_ADD_391_1196_U430, P2_ADD_391_1196_U431, P2_ADD_391_1196_U432, P2_ADD_391_1196_U433, P2_ADD_391_1196_U434, P2_ADD_391_1196_U435, P2_ADD_391_1196_U436, P2_ADD_391_1196_U437, P2_ADD_391_1196_U438, P2_ADD_391_1196_U439, P2_ADD_391_1196_U440, P2_ADD_391_1196_U441, P2_ADD_391_1196_U442, P2_ADD_391_1196_U443, P2_ADD_391_1196_U444, P2_ADD_391_1196_U445, P2_ADD_391_1196_U446, P2_ADD_391_1196_U447, P2_ADD_391_1196_U448, P2_ADD_391_1196_U449, P2_ADD_391_1196_U450, P2_ADD_391_1196_U451, P2_ADD_391_1196_U452, P2_ADD_391_1196_U453, P2_ADD_391_1196_U454, P2_ADD_391_1196_U455, P2_ADD_391_1196_U456, P2_ADD_391_1196_U457, P2_ADD_391_1196_U458, P2_ADD_391_1196_U459, P2_ADD_391_1196_U460, P2_ADD_391_1196_U461, P2_ADD_391_1196_U462, P2_ADD_391_1196_U463, P2_ADD_391_1196_U464, P2_ADD_391_1196_U465, P2_ADD_391_1196_U466, P2_ADD_391_1196_U467, P2_ADD_391_1196_U468, P2_ADD_391_1196_U469, P2_ADD_391_1196_U470, P2_ADD_391_1196_U471, P2_ADD_391_1196_U472, P2_ADD_391_1196_U473, P2_ADD_391_1196_U474, P2_ADD_391_1196_U475, P2_ADD_391_1196_U476, P2_ADD_391_1196_U477, P2_ADD_391_1196_U478, P2_ADD_402_1132_U4, P2_ADD_402_1132_U5, P2_ADD_402_1132_U6, P2_ADD_402_1132_U7, P2_ADD_402_1132_U8, P2_ADD_402_1132_U9, P2_ADD_402_1132_U10, P2_ADD_402_1132_U11, P2_ADD_402_1132_U12, P2_ADD_402_1132_U13, P2_ADD_402_1132_U14, P2_ADD_402_1132_U15, P2_ADD_402_1132_U16, P2_ADD_402_1132_U17, P2_ADD_402_1132_U18, P2_ADD_402_1132_U19, P2_ADD_402_1132_U20, P2_ADD_402_1132_U21, P2_ADD_402_1132_U22, P2_ADD_402_1132_U23, P2_ADD_402_1132_U24, P2_ADD_402_1132_U25, P2_ADD_402_1132_U26, P2_ADD_402_1132_U27, P2_ADD_402_1132_U28, P2_ADD_402_1132_U29, P2_ADD_402_1132_U30, P2_ADD_402_1132_U31, P2_ADD_402_1132_U32, P2_ADD_402_1132_U33, P2_ADD_402_1132_U34, P2_ADD_402_1132_U35, P2_ADD_402_1132_U36, P2_ADD_402_1132_U37, P2_ADD_402_1132_U38, P2_ADD_402_1132_U39, P2_ADD_402_1132_U40, P2_ADD_402_1132_U41, P2_ADD_402_1132_U42, P2_ADD_402_1132_U43, P2_ADD_402_1132_U44, P2_ADD_402_1132_U45, P2_ADD_402_1132_U46, P2_ADD_402_1132_U47, P2_ADD_402_1132_U48, P2_ADD_402_1132_U49, P2_ADD_402_1132_U50, P2_SUB_563_U6, P2_SUB_563_U7, P2_R2182_U4, P2_R2182_U5, P2_R2182_U6, P2_R2182_U7, P2_R2182_U8, P2_R2182_U9, P2_R2182_U10, P2_R2182_U11, P2_R2182_U12, P2_R2182_U13, P2_R2182_U14, P2_R2182_U15, P2_R2182_U16, P2_R2182_U17, P2_R2182_U18, P2_R2182_U19, P2_R2182_U20, P2_R2182_U21, P2_R2182_U22, P2_R2182_U23, P2_R2182_U24, P2_R2182_U25, P2_R2182_U26, P2_R2182_U27, P2_R2182_U28, P2_R2182_U29, P2_R2182_U30, P2_R2182_U31, P2_R2182_U32, P2_R2182_U33, P2_R2182_U34, P2_R2182_U35, P2_R2182_U36, P2_R2182_U37, P2_R2182_U38, P2_R2182_U39, P2_R2182_U40, P2_R2182_U41, P2_R2182_U42, P2_R2182_U43, P2_R2182_U44, P2_R2182_U45, P2_R2182_U46, P2_R2182_U47, P2_R2182_U48, P2_R2182_U49, P2_R2182_U50, P2_R2182_U51, P2_R2182_U52, P2_R2182_U53, P2_R2182_U54, P2_R2182_U55, P2_R2182_U56, P2_R2182_U57, P2_R2182_U58, P2_R2182_U59, P2_R2182_U60, P2_R2182_U61, P2_R2182_U62, P2_R2182_U63, P2_R2182_U64, P2_R2182_U65, P2_R2182_U66, P2_R2182_U67, P2_R2182_U68, P2_R2182_U69, P2_R2182_U70, P2_R2182_U71, P2_R2182_U72, P2_R2182_U73, P2_R2182_U74, P2_R2182_U75, P2_R2182_U76, P2_R2182_U77, P2_R2182_U78, P2_R2182_U79, P2_R2182_U80, P2_R2182_U81, P2_R2182_U82, P2_R2182_U83, P2_R2182_U84, P2_R2182_U85, P2_R2182_U86, P2_R2182_U87, P2_R2182_U88, P2_R2182_U89, P2_R2182_U90, P2_R2182_U91, P2_R2182_U92, P2_R2182_U93, P2_R2182_U94, P2_R2182_U95, P2_R2182_U96, P2_R2182_U97, P2_R2182_U98, P2_R2182_U99, P2_R2182_U100, P2_R2182_U101, P2_R2182_U102, P2_R2182_U103, P2_R2182_U104, P2_R2182_U105, P2_R2182_U106, P2_R2182_U107, P2_R2182_U108, P2_R2182_U109, P2_R2182_U110, P2_R2182_U111, P2_R2182_U112, P2_R2182_U113, P2_R2182_U114, P2_R2182_U115, P2_R2182_U116, P2_R2182_U117, P2_R2182_U118, P2_R2182_U119, P2_R2182_U120, P2_R2182_U121, P2_R2182_U122, P2_R2182_U123, P2_R2182_U124, P2_R2182_U125, P2_R2182_U126, P2_R2182_U127, P2_R2182_U128, P2_R2182_U129, P2_R2182_U130, P2_R2182_U131, P2_R2182_U132, P2_R2182_U133, P2_R2182_U134, P2_R2182_U135, P2_R2182_U136, P2_R2182_U137, P2_R2182_U138, P2_R2182_U139, P2_R2182_U140, P2_R2182_U141, P2_R2182_U142, P2_R2182_U143, P2_R2182_U144, P2_R2182_U145, P2_R2182_U146, P2_R2182_U147, P2_R2182_U148, P2_R2182_U149, P2_R2182_U150, P2_R2182_U151, P2_R2182_U152, P2_R2182_U153, P2_R2182_U154, P2_R2182_U155, P2_R2182_U156, P2_R2182_U157, P2_R2182_U158, P2_R2182_U159, P2_R2182_U160, P2_R2182_U161, P2_R2182_U162, P2_R2182_U163, P2_R2182_U164, P2_R2182_U165, P2_R2182_U166, P2_R2182_U167, P2_R2182_U168, P2_R2182_U169, P2_R2182_U170, P2_R2182_U171, P2_R2182_U172, P2_R2182_U173, P2_R2182_U174, P2_R2182_U175, P2_R2182_U176, P2_R2182_U177, P2_R2182_U178, P2_R2182_U179, P2_R2182_U180, P2_R2182_U181, P2_R2182_U182, P2_R2182_U183, P2_R2182_U184, P2_R2182_U185, P2_R2182_U186, P2_R2182_U187, P2_R2182_U188, P2_R2182_U189, P2_R2182_U190, P2_R2182_U191, P2_R2182_U192, P2_R2182_U193, P2_R2182_U194, P2_R2182_U195, P2_R2182_U196, P2_R2182_U197, P2_R2182_U198, P2_R2182_U199, P2_R2182_U200, P2_R2182_U201, P2_R2182_U202, P2_R2182_U203, P2_R2182_U204, P2_R2182_U205, P2_R2182_U206, P2_R2182_U207, P2_R2182_U208, P2_R2182_U209, P2_R2182_U210, P2_R2182_U211, P2_R2182_U212, P2_R2182_U213, P2_R2182_U214, P2_R2182_U215, P2_R2182_U216, P2_R2182_U217, P2_R2182_U218, P2_R2182_U219, P2_R2182_U220, P2_R2182_U221, P2_R2182_U222, P2_R2182_U223, P2_R2182_U224, P2_R2182_U225, P2_R2182_U226, P2_R2182_U227, P2_R2182_U228, P2_R2182_U229, P2_R2182_U230, P2_R2182_U231, P2_R2182_U232, P2_R2182_U233, P2_R2182_U234, P2_R2182_U235, P2_R2182_U236, P2_R2182_U237, P2_R2182_U238, P2_R2182_U239, P2_R2182_U240, P2_R2182_U241, P2_R2182_U242, P2_R2182_U243, P2_R2182_U244, P2_R2182_U245, P2_R2182_U246, P2_R2182_U247, P2_R2182_U248, P2_R2182_U249, P2_R2182_U250, P2_R2182_U251, P2_R2182_U252, P2_R2182_U253, P2_R2182_U254, P2_R2182_U255, P2_R2182_U256, P2_R2182_U257, P2_R2182_U258, P2_R2182_U259, P2_R2182_U260, P2_R2182_U261, P2_R2182_U262, P2_R2182_U263, P2_R2182_U264, P2_R2182_U265, P2_R2182_U266, P2_R2182_U267, P2_R2182_U268, P2_R2182_U269, P2_R2182_U270, P2_R2182_U271, P2_R2182_U272, P2_R2182_U273, P2_R2182_U274, P2_R2182_U275, P2_R2182_U276, P2_R2182_U277, P2_R2182_U278, P2_R2182_U279, P2_R2182_U280, P2_R2182_U281, P2_R2182_U282, P2_R2182_U283, P2_R2182_U284, P2_R2182_U285, P2_R2182_U286, P2_R2182_U287, P2_R2182_U288, P2_R2182_U289, P2_R2182_U290, P2_R2182_U291, P2_R2182_U292, P2_R2182_U293, P2_R2182_U294, P2_R2182_U295, P2_R2182_U296, P2_R2182_U297, P2_R2182_U298, P2_R2182_U299, P2_R2182_U300, P2_R2182_U301, P2_R2182_U302, P2_R2182_U303, P2_R2182_U304, P2_R2182_U305, P2_R2167_U6, P2_R2167_U7, P2_R2167_U8, P2_R2167_U9, P2_R2167_U10, P2_R2167_U11, P2_R2167_U12, P2_R2167_U13, P2_R2167_U14, P2_R2167_U15, P2_R2167_U16, P2_R2167_U17, P2_R2167_U18, P2_R2167_U19, P2_R2167_U20, P2_R2167_U21, P2_R2167_U22, P2_R2167_U23, P2_R2167_U24, P2_R2167_U25, P2_R2167_U26, P2_R2167_U27, P2_R2167_U28, P2_R2167_U29, P2_R2167_U30, P2_R2167_U31, P2_R2167_U32, P2_R2167_U33, P2_R2167_U34, P2_R2167_U35, P2_R2167_U36, P2_R2167_U37, P2_R2167_U38, P2_R2167_U39, P2_R2167_U40, P2_R2167_U41, P2_R2167_U42, P2_R2027_U5, P2_R2027_U6, P2_R2027_U7, P2_R2027_U8, P2_R2027_U9, P2_R2027_U10, P2_R2027_U11, P2_R2027_U12, P2_R2027_U13, P2_R2027_U14, P2_R2027_U15, P2_R2027_U16, P2_R2027_U17, P2_R2027_U18, P2_R2027_U19, P2_R2027_U20, P2_R2027_U21, P2_R2027_U22, P2_R2027_U23, P2_R2027_U24, P2_R2027_U25, P2_R2027_U26, P2_R2027_U27, P2_R2027_U28, P2_R2027_U29, P2_R2027_U30, P2_R2027_U31, P2_R2027_U32, P2_R2027_U33, P2_R2027_U34, P2_R2027_U35, P2_R2027_U36, P2_R2027_U37, P2_R2027_U38, P2_R2027_U39, P2_R2027_U40, P2_R2027_U41, P2_R2027_U42, P2_R2027_U43, P2_R2027_U44, P2_R2027_U45, P2_R2027_U46, P2_R2027_U47, P2_R2027_U48, P2_R2027_U49, P2_R2027_U50, P2_R2027_U51, P2_R2027_U52, P2_R2027_U53, P2_R2027_U54, P2_R2027_U55, P2_R2027_U56, P2_R2027_U57, P2_R2027_U58, P2_R2027_U59, P2_R2027_U60, P2_R2027_U61, P2_R2027_U62, P2_R2027_U63, P2_R2027_U64, P2_R2027_U65, P2_R2027_U66, P2_R2027_U67, P2_R2027_U68, P2_R2027_U69, P2_R2027_U70, P2_R2027_U71, P2_R2027_U72, P2_R2027_U73, P2_R2027_U74, P2_R2027_U75, P2_R2027_U76, P2_R2027_U77, P2_R2027_U78, P2_R2027_U79, P2_R2027_U80, P2_R2027_U81, P2_R2027_U82, P2_R2027_U83, P2_R2027_U84, P2_R2027_U85, P2_R2027_U86, P2_R2027_U87, P2_R2027_U88, P2_R2027_U89, P2_R2027_U90, P2_R2027_U91, P2_R2027_U92, P2_R2027_U93, P2_R2027_U94, P2_R2027_U95, P2_R2027_U96, P2_R2027_U97, P2_R2027_U98, P2_R2027_U99, P2_R2027_U100, P2_R2027_U101, P2_R2027_U102, P2_R2027_U103, P2_R2027_U104, P2_R2027_U105, P2_R2027_U106, P2_R2027_U107, P2_R2027_U108, P2_R2027_U109, P2_R2027_U110, P2_R2027_U111, P2_R2027_U112, P2_R2027_U113, P2_R2027_U114, P2_R2027_U115, P2_R2027_U116, P2_R2027_U117, P2_R2027_U118, P2_R2027_U119, P2_R2027_U120, P2_R2027_U121, P2_R2027_U122, P2_R2027_U123, P2_R2027_U124, P2_R2027_U125, P2_R2027_U126, P2_R2027_U127, P2_R2027_U128, P2_R2027_U129, P2_R2027_U130, P2_R2027_U131, P2_R2027_U132, P2_R2027_U133, P2_R2027_U134, P2_R2027_U135, P2_R2027_U136, P2_R2027_U137, P2_R2027_U138, P2_R2027_U139, P2_R2027_U140, P2_R2027_U141, P2_R2027_U142, P2_R2027_U143, P2_R2027_U144, P2_R2027_U145, P2_R2027_U146, P2_R2027_U147, P2_R2027_U148, P2_R2027_U149, P2_R2027_U150, P2_R2027_U151, P2_R2027_U152, P2_R2027_U153, P2_R2027_U154, P2_R2027_U155, P2_R2027_U156, P2_R2027_U157, P2_R2027_U158, P2_R2027_U159, P2_R2027_U160, P2_R2027_U161, P2_R2027_U162, P2_R2027_U163, P2_R2027_U164, P2_R2027_U165, P2_R2027_U166, P2_R2027_U167, P2_R2027_U168, P2_R2027_U169, P2_R2027_U170, P2_R2027_U171, P2_R2027_U172, P2_R2027_U173, P2_R2027_U174, P2_R2027_U175, P2_R2027_U176, P2_R2027_U177, P2_R2027_U178, P2_R2027_U179, P2_R2027_U180, P2_R2027_U181, P2_R2027_U182, P2_R2027_U183, P2_R2027_U184, P2_R2027_U185, P2_R2027_U186, P2_R2027_U187, P2_R2027_U188, P2_R2027_U189, P2_LT_563_1260_U6, P2_LT_563_1260_U7, P2_R2337_U4, P2_R2337_U5, P2_R2337_U6, P2_R2337_U7, P2_R2337_U8, P2_R2337_U9, P2_R2337_U10, P2_R2337_U11, P2_R2337_U12, P2_R2337_U13, P2_R2337_U14, P2_R2337_U15, P2_R2337_U16, P2_R2337_U17, P2_R2337_U18, P2_R2337_U19, P2_R2337_U20, P2_R2337_U21, P2_R2337_U22, P2_R2337_U23, P2_R2337_U24, P2_R2337_U25, P2_R2337_U26, P2_R2337_U27, P2_R2337_U28, P2_R2337_U29, P2_R2337_U30, P2_R2337_U31, P2_R2337_U32, P2_R2337_U33, P2_R2337_U34, P2_R2337_U35, P2_R2337_U36, P2_R2337_U37, P2_R2337_U38, P2_R2337_U39, P2_R2337_U40, P2_R2337_U41, P2_R2337_U42, P2_R2337_U43, P2_R2337_U44, P2_R2337_U45, P2_R2337_U46, P2_R2337_U47, P2_R2337_U48, P2_R2337_U49, P2_R2337_U50, P2_R2337_U51, P2_R2337_U52, P2_R2337_U53, P2_R2337_U54, P2_R2337_U55, P2_R2337_U56, P2_R2337_U57, P2_R2337_U58, P2_R2337_U59, P2_R2337_U60, P2_R2337_U61, P2_R2337_U62, P2_R2337_U63, P2_R2337_U64, P2_R2337_U65, P2_R2337_U66, P2_R2337_U67, P2_R2337_U68, P2_R2337_U69, P2_R2337_U70, P2_R2337_U71, P2_R2337_U72, P2_R2337_U73, P2_R2337_U74, P2_R2337_U75, P2_R2337_U76, P2_R2337_U77, P2_R2337_U78, P2_R2337_U79, P2_R2337_U80, P2_R2337_U81, P2_R2337_U82, P2_R2337_U83, P2_R2337_U84, P2_R2337_U85, P2_R2337_U86, P2_R2337_U87, P2_R2337_U88, P2_R2337_U89, P2_R2337_U90, P2_R2337_U91, P2_R2337_U92, P2_R2337_U93, P2_R2337_U94, P2_R2337_U95, P2_R2337_U96, P2_R2337_U97, P2_R2337_U98, P2_R2337_U99, P2_R2337_U100, P2_R2337_U101, P2_R2337_U102, P2_R2337_U103, P2_R2337_U104, P2_R2337_U105, P2_R2337_U106, P2_R2337_U107, P2_R2337_U108, P2_R2337_U109, P2_R2337_U110, P2_R2337_U111, P2_R2337_U112, P2_R2337_U113, P2_R2337_U114, P2_R2337_U115, P2_R2337_U116, P2_R2337_U117, P2_R2337_U118, P2_R2337_U119, P2_R2337_U120, P2_R2337_U121, P2_R2337_U122, P2_R2337_U123, P2_R2337_U124, P2_R2337_U125, P2_R2337_U126, P2_R2337_U127, P2_R2337_U128, P2_R2337_U129, P2_R2337_U130, P2_R2337_U131, P2_R2337_U132, P2_R2337_U133, P2_R2337_U134, P2_R2337_U135, P2_R2337_U136, P2_R2337_U137, P2_R2337_U138, P2_R2337_U139, P2_R2337_U140, P2_R2337_U141, P2_R2337_U142, P2_R2337_U143, P2_R2337_U144, P2_R2337_U145, P2_R2337_U146, P2_R2337_U147, P2_R2337_U148, P2_R2337_U149, P2_R2337_U150, P2_R2337_U151, P2_R2337_U152, P2_R2337_U153, P2_R2337_U154, P2_R2337_U155, P2_R2337_U156, P2_R2337_U157, P2_R2337_U158, P2_R2337_U159, P2_R2337_U160, P2_R2337_U161, P2_R2337_U162, P2_R2337_U163, P2_R2337_U164, P2_R2337_U165, P2_R2337_U166, P2_R2337_U167, P2_R2337_U168, P2_R2337_U169, P2_R2337_U170, P2_R2337_U171, P2_R2337_U172, P2_R2337_U173, P2_R2337_U174, P2_R2337_U175, P2_R2337_U176, P2_R2337_U177, P2_R2337_U178, P2_R2337_U179, P2_R2337_U180, P2_R2337_U181, P2_R2337_U182, P2_R2147_U4, P2_R2147_U5, P2_R2147_U6, P2_R2147_U7, P2_R2147_U8, P2_R2147_U9, P2_R2147_U10, P2_R2147_U11, P2_R2147_U12, P2_R2147_U13, P2_R2147_U14, P2_R2147_U15, P2_R2147_U16, P2_R2147_U17, P2_R2147_U18, P2_R2147_U19, P2_R2147_U20, P2_R2219_U6, P2_R2219_U7, P2_R2219_U8, P2_R2219_U9, P2_R2219_U10, P2_R2219_U11, P2_R2219_U12, P2_R2219_U13, P2_R2219_U14, P2_R2219_U15, P2_R2219_U16, P2_R2219_U17, P2_R2219_U18, P2_R2219_U19, P2_R2219_U20, P2_R2219_U21, P2_R2219_U22, P2_R2219_U23, P2_R2219_U24, P2_R2219_U25, P2_R2219_U26, P2_R2219_U27, P2_R2219_U28, P2_R2219_U29, P2_R2219_U30, P2_R2219_U31, P2_R2219_U32, P2_R2219_U33, P2_R2219_U34, P2_R2219_U35, P2_R2219_U36, P2_R2219_U37, P2_R2219_U38, P2_R2219_U39, P2_R2219_U40, P2_R2219_U41, P2_R2219_U42, P2_R2219_U43, P2_R2219_U44, P2_R2219_U45, P2_R2219_U46, P2_R2219_U47, P2_R2219_U48, P2_R2219_U49, P2_R2219_U50, P2_R2219_U51, P2_R2219_U52, P2_R2219_U53, P2_R2219_U54, P2_R2219_U55, P2_R2219_U56, P2_R2219_U57, P2_R2219_U58, P2_R2219_U59, P2_R2219_U60, P2_R2219_U61, P2_R2219_U62, P2_R2219_U63, P2_R2219_U64, P2_R2219_U65, P2_R2219_U66, P2_R2219_U67, P2_R2219_U68, P2_R2219_U69, P2_R2219_U70, P2_R2219_U71, P2_R2219_U72, P2_R2219_U73, P2_R2219_U74, P2_R2219_U75, P2_R2219_U76, P2_R2219_U77, P2_R2219_U78, P2_R2219_U79, P2_R2219_U80, P2_R2219_U81, P2_R2219_U82, P2_R2219_U83, P2_R2219_U84, P2_R2219_U85, P2_R2219_U86, P2_R2219_U87, P2_R2219_U88, P2_R2219_U89, P2_R2219_U90, P2_R2219_U91, P2_R2219_U92, P2_R2219_U93, P2_R2219_U94, P2_R2219_U95, P2_R2219_U96, P2_R2219_U97, P2_R2219_U98, P2_R2219_U99, P2_R2219_U100, P2_R2219_U101, P2_R2219_U102, P2_R2219_U103, P2_R2219_U104, P2_R2219_U105, P2_R2219_U106, P2_R2219_U107, P2_R2219_U108, P2_R2219_U109, P2_R2219_U110, P2_R2219_U111, P2_R2219_U112, P2_R2219_U113, P2_R2219_U114, P2_R2219_U115, P2_R2219_U116, P2_R2243_U6, P2_R2243_U7, P2_R2243_U8, P2_R2243_U9, P2_R2243_U10, P2_R2243_U11, P2_SUB_589_U6, P2_SUB_589_U7, P2_SUB_589_U8, P2_SUB_589_U9, P2_R2096_U4, P2_R2096_U5, P2_R2096_U6, P2_R2096_U7, P2_R2096_U8, P2_R2096_U9, P2_R2096_U10, P2_R2096_U11, P2_R2096_U12, P2_R2096_U13, P2_R2096_U14, P2_R2096_U15, P2_R2096_U16, P2_R2096_U17, P2_R2096_U18, P2_R2096_U19, P2_R2096_U20, P2_R2096_U21, P2_R2096_U22, P2_R2096_U23, P2_R2096_U24, P2_R2096_U25, P2_R2096_U26, P2_R2096_U27, P2_R2096_U28, P2_R2096_U29, P2_R2096_U30, P2_R2096_U31, P2_R2096_U32, P2_R2096_U33, P2_R2096_U34, P2_R2096_U35, P2_R2096_U36, P2_R2096_U37, P2_R2096_U38, P2_R2096_U39, P2_R2096_U40, P2_R2096_U41, P2_R2096_U42, P2_R2096_U43, P2_R2096_U44, P2_R2096_U45, P2_R2096_U46, P2_R2096_U47, P2_R2096_U48, P2_R2096_U49, P2_R2096_U50, P2_R2096_U51, P2_R2096_U52, P2_R2096_U53, P2_R2096_U54, P2_R2096_U55, P2_R2096_U56, P2_R2096_U57, P2_R2096_U58, P2_R2096_U59, P2_R2096_U60, P2_R2096_U61, P2_R2096_U62, P2_R2096_U63, P2_R2096_U64, P2_R2096_U65, P2_R2096_U66, P2_R2096_U67, P2_R2096_U68, P2_R2096_U69, P2_R2096_U70, P2_R2096_U71, P2_R2096_U72, P2_R2096_U73, P2_R2096_U74, P2_R2096_U75, P2_R2096_U76, P2_R2096_U77, P2_R2096_U78, P2_R2096_U79, P2_R2096_U80, P2_R2096_U81, P2_R2096_U82, P2_R2096_U83, P2_R2096_U84, P2_R2096_U85, P2_R2096_U86, P2_R2096_U87, P2_R2096_U88, P2_R2096_U89, P2_R2096_U90, P2_R2096_U91, P2_R2096_U92, P2_R2096_U93, P2_R2096_U94, P2_R2096_U95, P2_R2096_U96, P2_R2096_U97, P2_R2096_U98, P2_R2096_U99, P2_R2096_U100, P2_R2096_U101, P2_R2096_U102, P2_R2096_U103, P2_R2096_U104, P2_R2096_U105, P2_R2096_U106, P2_R2096_U107, P2_R2096_U108, P2_R2096_U109, P2_R2096_U110, P2_R2096_U111, P2_R2096_U112, P2_R2096_U113, P2_R2096_U114, P2_R2096_U115, P2_R2096_U116, P2_R2096_U117, P2_R2096_U118, P2_R2096_U119, P2_R2096_U120, P2_R2096_U121, P2_R2096_U122, P2_R2096_U123, P2_R2096_U124, P2_R2096_U125, P2_R2096_U126, P2_R2096_U127, P2_R2096_U128, P2_R2096_U129, P2_R2096_U130, P2_R2096_U131, P2_R2096_U132, P2_R2096_U133, P2_R2096_U134, P2_R2096_U135, P2_R2096_U136, P2_R2096_U137, P2_R2096_U138, P2_R2096_U139, P2_R2096_U140, P2_R2096_U141, P2_R2096_U142, P2_R2096_U143, P2_R2096_U144, P2_R2096_U145, P2_R2096_U146, P2_R2096_U147, P2_R2096_U148, P2_R2096_U149, P2_R2096_U150, P2_R2096_U151, P2_R2096_U152, P2_R2096_U153, P2_R2096_U154, P2_R2096_U155, P2_R2096_U156, P2_R2096_U157, P2_R2096_U158, P2_R2096_U159, P2_R2096_U160, P2_R2096_U161, P2_R2096_U162, P2_R2096_U163, P2_R2096_U164, P2_R2096_U165, P2_R2096_U166, P2_R2096_U167, P2_R2096_U168, P2_R2096_U169, P2_R2096_U170, P2_R2096_U171, P2_R2096_U172, P2_R2096_U173, P2_R2096_U174, P2_R2096_U175, P2_R2096_U176, P2_R2096_U177, P2_R2096_U178, P2_R2096_U179, P2_R2096_U180, P2_R2096_U181, P2_R2096_U182, P2_R2096_U183, P2_R2096_U184, P2_R2096_U185, P2_R2096_U186, P2_R2096_U187, P2_R2096_U188, P2_R2096_U189, P2_R2096_U190, P2_R2096_U191, P2_R2096_U192, P2_R2096_U193, P2_R2096_U194, P2_R2096_U195, P2_R2096_U196, P2_R2096_U197, P2_R2096_U198, P2_R2096_U199, P2_R2096_U200, P2_R2096_U201, P2_R2096_U202, P2_R2096_U203, P2_R2096_U204, P2_R2096_U205, P2_R2096_U206, P2_R2096_U207, P2_R2096_U208, P2_R2096_U209, P2_R2096_U210, P2_R2096_U211, P2_R2096_U212, P2_R2096_U213, P2_R2096_U214, P2_R2096_U215, P2_R2096_U216, P2_R2096_U217, P2_R2096_U218, P2_R2096_U219, P2_R2096_U220, P2_R2096_U221, P2_R2096_U222, P2_R2096_U223, P2_R2096_U224, P2_R2096_U225, P2_R2096_U226, P2_R2096_U227, P2_R2096_U228, P2_R2096_U229, P2_R2096_U230, P2_R2096_U231, P2_R2096_U232, P2_R2096_U233, P2_R2096_U234, P2_R2096_U235, P2_R2096_U236, P2_R2096_U237, P2_R2096_U238, P2_R2096_U239, P2_R2096_U240, P2_R2096_U241, P2_R2096_U242, P2_R2096_U243, P2_R2096_U244, P2_R2096_U245, P2_R2096_U246, P2_R2096_U247, P2_R2096_U248, P2_R2096_U249, P2_R2096_U250, P2_R2096_U251, P2_R2096_U252, P2_R2096_U253, P2_R2096_U254, P2_R2096_U255, P2_R2096_U256, P2_R2096_U257, P2_R2096_U258, P2_R2096_U259, P2_R2096_U260, P2_R2096_U261, P2_R2096_U262, P2_R2096_U263, P2_R2096_U264, P2_R2096_U265, P2_GTE_370_U6, P2_GTE_370_U7, P2_GTE_370_U8, P2_GTE_370_U9, P2_LT_563_U6, P2_LT_563_U7, P2_LT_563_U8, P2_LT_563_U9, P2_LT_563_U10, P2_LT_563_U11, P2_LT_563_U12, P2_LT_563_U13, P2_LT_563_U14, P2_LT_563_U15, P2_LT_563_U16, P2_LT_563_U17, P2_LT_563_U18, P2_LT_563_U19, P2_LT_563_U20, P2_LT_563_U21, P2_LT_563_U22, P2_LT_563_U23, P2_LT_563_U24, P2_LT_563_U25, P2_LT_563_U26, P2_LT_563_U27, P2_R2256_U4, P2_R2256_U5, P2_R2256_U6, P2_R2256_U7, P2_R2256_U8, P2_R2256_U9, P2_R2256_U10, P2_R2256_U11, P2_R2256_U12, P2_R2256_U13, P2_R2256_U14, P2_R2256_U15, P2_R2256_U16, P2_R2256_U17, P2_R2256_U18, P2_R2256_U19, P2_R2256_U20, P2_R2256_U21, P2_R2256_U22, P2_R2256_U23, P2_R2256_U24, P2_R2256_U25, P2_R2256_U26, P2_R2256_U27, P2_R2256_U28, P2_R2256_U29, P2_R2256_U30, P2_R2256_U31, P2_R2256_U32, P2_R2256_U33, P2_R2256_U34, P2_R2256_U35, P2_R2256_U36, P2_R2256_U37, P2_R2256_U38, P2_R2256_U39, P2_R2256_U40, P2_R2256_U41, P2_R2256_U42, P2_R2256_U43, P2_R2256_U44, P2_R2256_U45, P2_R2256_U46, P2_R2256_U47, P2_R2256_U48, P2_R2256_U49, P2_R2256_U50, P2_R2256_U51, P2_R2256_U52, P2_R2256_U53, P2_R2256_U54, P2_R2256_U55, P2_R2256_U56, P2_R2256_U57, P2_R2256_U58, P2_R2256_U59, P2_R2256_U60, P2_R2256_U61, P2_R2256_U62, P2_R2256_U63, P2_R2256_U64, P2_R2256_U65, P2_R2256_U66, P2_R2256_U67, P2_R2256_U68, P2_R2256_U69, P2_R2256_U70, P2_R2238_U6, P2_R2238_U7, P2_R2238_U8, P2_R2238_U9, P2_R2238_U10, P2_R2238_U11, P2_R2238_U12, P2_R2238_U13, P2_R2238_U14, P2_R2238_U15, P2_R2238_U16, P2_R2238_U17, P2_R2238_U18, P2_R2238_U19, P2_R2238_U20, P2_R2238_U21, P2_R2238_U22, P2_R2238_U23, P2_R2238_U24, P2_R2238_U25, P2_R2238_U26, P2_R2238_U27, P2_R2238_U28, P2_R2238_U29, P2_R2238_U30, P2_R2238_U31, P2_R2238_U32, P2_R2238_U33, P2_R2238_U34, P2_R2238_U35, P2_R2238_U36, P2_R2238_U37, P2_R2238_U38, P2_R2238_U39, P2_R2238_U40, P2_R2238_U41, P2_R2238_U42, P2_R2238_U43, P2_R2238_U44, P2_R2238_U45, P2_R2238_U46, P2_R2238_U47, P2_R2238_U48, P2_R2238_U49, P2_R2238_U50, P2_R2238_U51, P2_R2238_U52, P2_R2238_U53, P2_R2238_U54, P2_R2238_U55, P2_R2238_U56, P2_R2238_U57, P2_R2238_U58, P2_R2238_U59, P2_R2238_U60, P2_R2238_U61, P2_R2238_U62, P2_R2238_U63, P2_R2238_U64, P2_R2238_U65, P2_R2238_U66, P2_R1957_U6, P2_R1957_U7, P2_R1957_U8, P2_R1957_U9, P2_R1957_U10, P2_R1957_U11, P2_R1957_U12, P2_R1957_U13, P2_R1957_U14, P2_R1957_U15, P2_R1957_U16, P2_R1957_U17, P2_R1957_U18, P2_R1957_U19, P2_R1957_U20, P2_R1957_U21, P2_R1957_U22, P2_R1957_U23, P2_R1957_U24, P2_R1957_U25, P2_R1957_U26, P2_R1957_U27, P2_R1957_U28, P2_R1957_U29, P2_R1957_U30, P2_R1957_U31, P2_R1957_U32, P2_R1957_U33, P2_R1957_U34, P2_R1957_U35, P2_R1957_U36, P2_R1957_U37, P2_R1957_U38, P2_R1957_U39, P2_R1957_U40, P2_R1957_U41, P2_R1957_U42, P2_R1957_U43, P2_R1957_U44, P2_R1957_U45, P2_R1957_U46, P2_R1957_U47, P2_R1957_U48, P2_R1957_U49, P2_R1957_U50, P2_R1957_U51, P2_R1957_U52, P2_R1957_U53, P2_R1957_U54, P2_R1957_U55, P2_R1957_U56, P2_R1957_U57, P2_R1957_U58, P2_R1957_U59, P2_R1957_U60, P2_R1957_U61, P2_R1957_U62, P2_R1957_U63, P2_R1957_U64, P2_R1957_U65, P2_R1957_U66, P2_R1957_U67, P2_R1957_U68, P2_R1957_U69, P2_R1957_U70, P2_R1957_U71, P2_R1957_U72, P2_R1957_U73, P2_R1957_U74, P2_R1957_U75, P2_R1957_U76, P2_R1957_U77, P2_R1957_U78, P2_R1957_U79, P2_R1957_U80, P2_R1957_U81, P2_R1957_U82, P2_R1957_U83, P2_R1957_U84, P2_R1957_U85, P2_R1957_U86, P2_R1957_U87, P2_R1957_U88, P2_R1957_U89, P2_R1957_U90, P2_R1957_U91, P2_R1957_U92, P2_R1957_U93, P2_R1957_U94, P2_R1957_U95, P2_R1957_U96, P2_R1957_U97, P2_R1957_U98, P2_R1957_U99, P2_R1957_U100, P2_R1957_U101, P2_R1957_U102, P2_R1957_U103, P2_R1957_U104, P2_R1957_U105, P2_R1957_U106, P2_R1957_U107, P2_R1957_U108, P2_R1957_U109, P2_R1957_U110, P2_R1957_U111, P2_R1957_U112, P2_R1957_U113, P2_R1957_U114, P2_R1957_U115, P2_R1957_U116, P2_R1957_U117, P2_R1957_U118, P2_R1957_U119, P2_R1957_U120, P2_R1957_U121, P2_R1957_U122, P2_R1957_U123, P2_R1957_U124, P2_R1957_U125, P2_R1957_U126, P2_R1957_U127, P2_R1957_U128, P2_R1957_U129, P2_R1957_U130, P2_R1957_U131, P2_R1957_U132, P2_R1957_U133, P2_R1957_U134, P2_R1957_U135, P2_R1957_U136, P2_R1957_U137, P2_R1957_U138, P2_R1957_U139, P2_R1957_U140, P2_R1957_U141, P2_R1957_U142, P2_R1957_U143, P2_R1957_U144, P2_R1957_U145, P2_R1957_U146, P2_R1957_U147, P2_R1957_U148, P2_R1957_U149, P2_R1957_U150, P2_R1957_U151, P2_R1957_U152, P2_R1957_U153, P2_R1957_U154, P2_R1957_U155, P2_R1957_U156, P2_R1957_U157, P2_R1957_U158, P2_R1957_U159, P2_R2278_U4, P2_R2278_U5, P2_R2278_U6, P2_R2278_U7, P2_R2278_U8, P2_R2278_U9, P2_R2278_U10, P2_R2278_U11, P2_R2278_U12, P2_R2278_U13, P2_R2278_U14, P2_R2278_U15, P2_R2278_U16, P2_R2278_U17, P2_R2278_U18, P2_R2278_U19, P2_R2278_U20, P2_R2278_U21, P2_R2278_U22, P2_R2278_U23, P2_R2278_U24, P2_R2278_U25, P2_R2278_U26, P2_R2278_U27, P2_R2278_U28, P2_R2278_U29, P2_R2278_U30, P2_R2278_U31, P2_R2278_U32, P2_R2278_U33, P2_R2278_U34, P2_R2278_U35, P2_R2278_U36, P2_R2278_U37, P2_R2278_U38, P2_R2278_U39, P2_R2278_U40, P2_R2278_U41, P2_R2278_U42, P2_R2278_U43, P2_R2278_U44, P2_R2278_U45, P2_R2278_U46, P2_R2278_U47, P2_R2278_U48, P2_R2278_U49, P2_R2278_U50, P2_R2278_U51, P2_R2278_U52, P2_R2278_U53, P2_R2278_U54, P2_R2278_U55, P2_R2278_U56, P2_R2278_U57, P2_R2278_U58, P2_R2278_U59, P2_R2278_U60, P2_R2278_U61, P2_R2278_U62, P2_R2278_U63, P2_R2278_U64, P2_R2278_U65, P2_R2278_U66, P2_R2278_U67, P2_R2278_U68, P2_R2278_U69, P2_R2278_U70, P2_R2278_U71, P2_R2278_U72, P2_R2278_U73, P2_R2278_U74, P2_R2278_U75, P2_R2278_U76, P2_R2278_U77, P2_R2278_U78, P2_R2278_U79, P2_R2278_U80, P2_R2278_U81, P2_R2278_U82, P2_R2278_U83, P2_R2278_U84, P2_R2278_U85, P2_R2278_U86, P2_R2278_U87, P2_R2278_U88, P2_R2278_U89, P2_R2278_U90, P2_R2278_U91, P2_R2278_U92, P2_R2278_U93, P2_R2278_U94, P2_R2278_U95, P2_R2278_U96, P2_R2278_U97, P2_R2278_U98, P2_R2278_U99, P2_R2278_U100, P2_R2278_U101, P2_R2278_U102, P2_R2278_U103, P2_R2278_U104, P2_R2278_U105, P2_R2278_U106, P2_R2278_U107, P2_R2278_U108, P2_R2278_U109, P2_R2278_U110, P2_R2278_U111, P2_R2278_U112, P2_R2278_U113, P2_R2278_U114, P2_R2278_U115, P2_R2278_U116, P2_R2278_U117, P2_R2278_U118, P2_R2278_U119, P2_R2278_U120, P2_R2278_U121, P2_R2278_U122, P2_R2278_U123, P2_R2278_U124, P2_R2278_U125, P2_R2278_U126, P2_R2278_U127, P2_R2278_U128, P2_R2278_U129, P2_R2278_U130, P2_R2278_U131, P2_R2278_U132, P2_R2278_U133, P2_R2278_U134, P2_R2278_U135, P2_R2278_U136, P2_R2278_U137, P2_R2278_U138, P2_R2278_U139, P2_R2278_U140, P2_R2278_U141, P2_R2278_U142, P2_R2278_U143, P2_R2278_U144, P2_R2278_U145, P2_R2278_U146, P2_R2278_U147, P2_R2278_U148, P2_R2278_U149, P2_R2278_U150, P2_R2278_U151, P2_R2278_U152, P2_R2278_U153, P2_R2278_U154, P2_R2278_U155, P2_R2278_U156, P2_R2278_U157, P2_R2278_U158, P2_R2278_U159, P2_R2278_U160, P2_R2278_U161, P2_R2278_U162, P2_R2278_U163, P2_R2278_U164, P2_R2278_U165, P2_R2278_U166, P2_R2278_U167, P2_R2278_U168, P2_R2278_U169, P2_R2278_U170, P2_R2278_U171, P2_R2278_U172, P2_R2278_U173, P2_R2278_U174, P2_R2278_U175, P2_R2278_U176, P2_R2278_U177, P2_R2278_U178, P2_R2278_U179, P2_R2278_U180, P2_R2278_U181, P2_R2278_U182, P2_R2278_U183, P2_R2278_U184, P2_R2278_U185, P2_R2278_U186, P2_R2278_U187, P2_R2278_U188, P2_R2278_U189, P2_R2278_U190, P2_R2278_U191, P2_R2278_U192, P2_R2278_U193, P2_R2278_U194, P2_R2278_U195, P2_R2278_U196, P2_R2278_U197, P2_R2278_U198, P2_R2278_U199, P2_R2278_U200, P2_R2278_U201, P2_R2278_U202, P2_R2278_U203, P2_R2278_U204, P2_R2278_U205, P2_R2278_U206, P2_R2278_U207, P2_R2278_U208, P2_R2278_U209, P2_R2278_U210, P2_R2278_U211, P2_R2278_U212, P2_R2278_U213, P2_R2278_U214, P2_R2278_U215, P2_R2278_U216, P2_R2278_U217, P2_R2278_U218, P2_R2278_U219, P2_R2278_U220, P2_R2278_U221, P2_R2278_U222, P2_R2278_U223, P2_R2278_U224, P2_R2278_U225, P2_R2278_U226, P2_R2278_U227, P2_R2278_U228, P2_R2278_U229, P2_R2278_U230, P2_R2278_U231, P2_R2278_U232, P2_R2278_U233, P2_R2278_U234, P2_R2278_U235, P2_R2278_U236, P2_R2278_U237, P2_R2278_U238, P2_R2278_U239, P2_R2278_U240, P2_R2278_U241, P2_R2278_U242, P2_R2278_U243, P2_R2278_U244, P2_R2278_U245, P2_R2278_U246, P2_R2278_U247, P2_R2278_U248, P2_R2278_U249, P2_R2278_U250, P2_R2278_U251, P2_R2278_U252, P2_R2278_U253, P2_R2278_U254, P2_R2278_U255, P2_R2278_U256, P2_R2278_U257, P2_R2278_U258, P2_R2278_U259, P2_R2278_U260, P2_R2278_U261, P2_R2278_U262, P2_R2278_U263, P2_R2278_U264, P2_R2278_U265, P2_R2278_U266, P2_R2278_U267, P2_R2278_U268, P2_R2278_U269, P2_R2278_U270, P2_R2278_U271, P2_R2278_U272, P2_R2278_U273, P2_R2278_U274, P2_R2278_U275, P2_R2278_U276, P2_R2278_U277, P2_R2278_U278, P2_R2278_U279, P2_R2278_U280, P2_R2278_U281, P2_R2278_U282, P2_R2278_U283, P2_R2278_U284, P2_R2278_U285, P2_R2278_U286, P2_R2278_U287, P2_R2278_U288, P2_R2278_U289, P2_R2278_U290, P2_R2278_U291, P2_R2278_U292, P2_R2278_U293, P2_R2278_U294, P2_R2278_U295, P2_R2278_U296, P2_R2278_U297, P2_R2278_U298, P2_R2278_U299, P2_R2278_U300, P2_R2278_U301, P2_R2278_U302, P2_R2278_U303, P2_R2278_U304, P2_R2278_U305, P2_R2278_U306, P2_R2278_U307, P2_R2278_U308, P2_R2278_U309, P2_R2278_U310, P2_R2278_U311, P2_R2278_U312, P2_R2278_U313, P2_R2278_U314, P2_R2278_U315, P2_R2278_U316, P2_R2278_U317, P2_R2278_U318, P2_R2278_U319, P2_R2278_U320, P2_R2278_U321, P2_R2278_U322, P2_R2278_U323, P2_R2278_U324, P2_R2278_U325, P2_R2278_U326, P2_R2278_U327, P2_R2278_U328, P2_R2278_U329, P2_R2278_U330, P2_R2278_U331, P2_R2278_U332, P2_R2278_U333, P2_R2278_U334, P2_R2278_U335, P2_R2278_U336, P2_R2278_U337, P2_R2278_U338, P2_R2278_U339, P2_R2278_U340, P2_R2278_U341, P2_R2278_U342, P2_R2278_U343, P2_R2278_U344, P2_R2278_U345, P2_R2278_U346, P2_R2278_U347, P2_R2278_U348, P2_R2278_U349, P2_R2278_U350, P2_R2278_U351, P2_R2278_U352, P2_R2278_U353, P2_R2278_U354, P2_R2278_U355, P2_R2278_U356, P2_R2278_U357, P2_R2278_U358, P2_R2278_U359, P2_R2278_U360, P2_R2278_U361, P2_R2278_U362, P2_R2278_U363, P2_R2278_U364, P2_R2278_U365, P2_R2278_U366, P2_R2278_U367, P2_R2278_U368, P2_R2278_U369, P2_R2278_U370, P2_R2278_U371, P2_R2278_U372, P2_R2278_U373, P2_R2278_U374, P2_R2278_U375, P2_R2278_U376, P2_R2278_U377, P2_R2278_U378, P2_R2278_U379, P2_R2278_U380, P2_R2278_U381, P2_R2278_U382, P2_R2278_U383, P2_R2278_U384, P2_R2278_U385, P2_R2278_U386, P2_R2278_U387, P2_R2278_U388, P2_R2278_U389, P2_R2278_U390, P2_R2278_U391, P2_R2278_U392, P2_R2278_U393, P2_R2278_U394, P2_R2278_U395, P2_R2278_U396, P2_R2278_U397, P2_R2278_U398, P2_R2278_U399, P2_R2278_U400, P2_R2278_U401, P2_R2278_U402, P2_R2278_U403, P2_R2278_U404, P2_R2278_U405, P2_R2278_U406, P2_R2278_U407, P2_R2278_U408, P2_R2278_U409, P2_R2278_U410, P2_R2278_U411, P2_R2278_U412, P2_R2278_U413, P2_R2278_U414, P2_R2278_U415, P2_R2278_U416, P2_R2278_U417, P2_R2278_U418, P2_R2278_U419, P2_R2278_U420, P2_R2278_U421, P2_R2278_U422, P2_R2278_U423, P2_R2278_U424, P2_R2278_U425, P2_R2278_U426, P2_R2278_U427, P2_R2278_U428, P2_R2278_U429, P2_R2278_U430, P2_R2278_U431, P2_R2278_U432, P2_R2278_U433, P2_R2278_U434, P2_R2278_U435, P2_R2278_U436, P2_R2278_U437, P2_R2278_U438, P2_R2278_U439, P2_R2278_U440, P2_R2278_U441, P2_R2278_U442, P2_R2278_U443, P2_R2278_U444, P2_R2278_U445, P2_R2278_U446, P2_R2278_U447, P2_R2278_U448, P2_R2278_U449, P2_R2278_U450, P2_R2278_U451, P2_R2278_U452, P2_R2278_U453, P2_R2278_U454, P2_R2278_U455, P2_R2278_U456, P2_R2278_U457, P2_R2278_U458, P2_R2278_U459, P2_R2278_U460, P2_R2278_U461, P2_R2278_U462, P2_R2278_U463, P2_R2278_U464, P2_R2278_U465, P2_R2278_U466, P2_R2278_U467, P2_R2278_U468, P2_R2278_U469, P2_R2278_U470, P2_R2278_U471, P2_R2278_U472, P2_R2278_U473, P2_R2278_U474, P2_R2278_U475, P2_R2278_U476, P2_R2278_U477, P2_R2278_U478, P2_R2278_U479, P2_R2278_U480, P2_R2278_U481, P2_R2278_U482, P2_R2278_U483, P2_R2278_U484, P2_R2278_U485, P2_R2278_U486, P2_R2278_U487, P2_R2278_U488, P2_R2278_U489, P2_R2278_U490, P2_R2278_U491, P2_R2278_U492, P2_R2278_U493, P2_R2278_U494, P2_R2278_U495, P2_R2278_U496, P2_R2278_U497, P2_R2278_U498, P2_R2278_U499, P2_R2278_U500, P2_R2278_U501, P2_R2278_U502, P2_R2278_U503, P2_R2278_U504, P2_R2278_U505, P2_R2278_U506, P2_R2278_U507, P2_R2278_U508, P2_R2278_U509, P2_R2278_U510, P2_R2278_U511, P2_R2278_U512, P2_R2278_U513, P2_R2278_U514, P2_R2278_U515, P2_R2278_U516, P2_R2278_U517, P2_R2278_U518, P2_R2278_U519, P2_R2278_U520, P2_R2278_U521, P2_R2278_U522, P2_R2278_U523, P2_R2278_U524, P2_R2278_U525, P2_R2278_U526, P2_R2278_U527, P2_R2278_U528, P2_R2278_U529, P2_R2278_U530, P2_R2278_U531, P2_R2278_U532, P2_R2278_U533, P2_R2278_U534, P2_R2278_U535, P2_R2278_U536, P2_R2278_U537, P2_R2278_U538, P2_R2278_U539, P2_R2278_U540, P2_R2278_U541, P2_R2278_U542, P2_R2278_U543, P2_R2278_U544, P2_R2278_U545, P2_R2278_U546, P2_R2278_U547, P2_R2278_U548, P2_R2278_U549, P2_R2278_U550, P2_R2278_U551, P2_R2278_U552, P2_R2278_U553, P2_R2278_U554, P2_R2278_U555, P2_R2278_U556, P2_R2278_U557, P2_R2278_U558, P2_R2278_U559, P2_R2278_U560, P2_R2278_U561, P2_R2278_U562, P2_SUB_450_U6, P2_SUB_450_U7, P2_SUB_450_U8, P2_SUB_450_U9, P2_SUB_450_U10, P2_SUB_450_U11, P2_SUB_450_U12, P2_SUB_450_U13, P2_SUB_450_U14, P2_SUB_450_U15, P2_SUB_450_U16, P2_SUB_450_U17, P2_SUB_450_U18, P2_SUB_450_U19, P2_SUB_450_U20, P2_SUB_450_U21, P2_SUB_450_U22, P2_SUB_450_U23, P2_SUB_450_U24, P2_SUB_450_U25, P2_SUB_450_U26, P2_SUB_450_U27, P2_SUB_450_U28, P2_SUB_450_U29, P2_SUB_450_U30, P2_SUB_450_U31, P2_SUB_450_U32, P2_SUB_450_U33, P2_SUB_450_U34, P2_SUB_450_U35, P2_SUB_450_U36, P2_SUB_450_U37, P2_SUB_450_U38, P2_SUB_450_U39, P2_SUB_450_U40, P2_SUB_450_U41, P2_SUB_450_U42, P2_SUB_450_U43, P2_SUB_450_U44, P2_SUB_450_U45, P2_SUB_450_U46, P2_SUB_450_U47, P2_SUB_450_U48, P2_SUB_450_U49, P2_SUB_450_U50, P2_SUB_450_U51, P2_SUB_450_U52, P2_SUB_450_U53, P2_SUB_450_U54, P2_SUB_450_U55, P2_SUB_450_U56, P2_SUB_450_U57, P2_SUB_450_U58, P2_SUB_450_U59, P2_SUB_450_U60, P2_SUB_450_U61, P2_SUB_450_U62, P2_SUB_450_U63, P2_R2088_U6, P2_R2088_U7, P2_ADD_394_U4, P2_ADD_394_U5, P2_ADD_394_U6, P2_ADD_394_U7, P2_ADD_394_U8, P2_ADD_394_U9, P2_ADD_394_U10, P2_ADD_394_U11, P2_ADD_394_U12, P2_ADD_394_U13, P2_ADD_394_U14, P2_ADD_394_U15, P2_ADD_394_U16, P2_ADD_394_U17, P2_ADD_394_U18, P2_ADD_394_U19, P2_ADD_394_U20, P2_ADD_394_U21, P2_ADD_394_U22, P2_ADD_394_U23, P2_ADD_394_U24, P2_ADD_394_U25, P2_ADD_394_U26, P2_ADD_394_U27, P2_ADD_394_U28, P2_ADD_394_U29, P2_ADD_394_U30, P2_ADD_394_U31, P2_ADD_394_U32, P2_ADD_394_U33, P2_ADD_394_U34, P2_ADD_394_U35, P2_ADD_394_U36, P2_ADD_394_U37, P2_ADD_394_U38, P2_ADD_394_U39, P2_ADD_394_U40, P2_ADD_394_U41, P2_ADD_394_U42, P2_ADD_394_U43, P2_ADD_394_U44, P2_ADD_394_U45, P2_ADD_394_U46, P2_ADD_394_U47, P2_ADD_394_U48, P2_ADD_394_U49, P2_ADD_394_U50, P2_ADD_394_U51, P2_ADD_394_U52, P2_ADD_394_U53, P2_ADD_394_U54, P2_ADD_394_U55, P2_ADD_394_U56, P2_ADD_394_U57, P2_ADD_394_U58, P2_ADD_394_U59, P2_ADD_394_U60, P2_ADD_394_U61, P2_ADD_394_U62, P2_ADD_394_U63, P2_ADD_394_U64, P2_ADD_394_U65, P2_ADD_394_U66, P2_ADD_394_U67, P2_ADD_394_U68, P2_ADD_394_U69, P2_ADD_394_U70, P2_ADD_394_U71, P2_ADD_394_U72, P2_ADD_394_U73, P2_ADD_394_U74, P2_ADD_394_U75, P2_ADD_394_U76, P2_ADD_394_U77, P2_ADD_394_U78, P2_ADD_394_U79, P2_ADD_394_U80, P2_ADD_394_U81, P2_ADD_394_U82, P2_ADD_394_U83, P2_ADD_394_U84, P2_ADD_394_U85, P2_ADD_394_U86, P2_ADD_394_U87, P2_ADD_394_U88, P2_ADD_394_U89, P2_ADD_394_U90, P2_ADD_394_U91, P2_ADD_394_U92, P2_ADD_394_U93, P2_ADD_394_U94, P2_ADD_394_U95, P2_ADD_394_U96, P2_ADD_394_U97, P2_ADD_394_U98, P2_ADD_394_U99, P2_ADD_394_U100, P2_ADD_394_U101, P2_ADD_394_U102, P2_ADD_394_U103, P2_ADD_394_U104, P2_ADD_394_U105, P2_ADD_394_U106, P2_ADD_394_U107, P2_ADD_394_U108, P2_ADD_394_U109, P2_ADD_394_U110, P2_ADD_394_U111, P2_ADD_394_U112, P2_ADD_394_U113, P2_ADD_394_U114, P2_ADD_394_U115, P2_ADD_394_U116, P2_ADD_394_U117, P2_ADD_394_U118, P2_ADD_394_U119, P2_ADD_394_U120, P2_ADD_394_U121, P2_ADD_394_U122, P2_ADD_394_U123, P2_ADD_394_U124, P2_ADD_394_U125, P2_ADD_394_U126, P2_ADD_394_U127, P2_ADD_394_U128, P2_ADD_394_U129, P2_ADD_394_U130, P2_ADD_394_U131, P2_ADD_394_U132, P2_ADD_394_U133, P2_ADD_394_U134, P2_ADD_394_U135, P2_ADD_394_U136, P2_ADD_394_U137, P2_ADD_394_U138, P2_ADD_394_U139, P2_ADD_394_U140, P2_ADD_394_U141, P2_ADD_394_U142, P2_ADD_394_U143, P2_ADD_394_U144, P2_ADD_394_U145, P2_ADD_394_U146, P2_ADD_394_U147, P2_ADD_394_U148, P2_ADD_394_U149, P2_ADD_394_U150, P2_ADD_394_U151, P2_ADD_394_U152, P2_ADD_394_U153, P2_ADD_394_U154, P2_ADD_394_U155, P2_ADD_394_U156, P2_ADD_394_U157, P2_ADD_394_U158, P2_ADD_394_U159, P2_ADD_394_U160, P2_ADD_394_U161, P2_ADD_394_U162, P2_ADD_394_U163, P2_ADD_394_U164, P2_ADD_394_U165, P2_ADD_394_U166, P2_ADD_394_U167, P2_ADD_394_U168, P2_ADD_394_U169, P2_ADD_394_U170, P2_ADD_394_U171, P2_ADD_394_U172, P2_ADD_394_U173, P2_ADD_394_U174, P2_ADD_394_U175, P2_ADD_394_U176, P2_ADD_394_U177, P2_ADD_394_U178, P2_ADD_394_U179, P2_ADD_394_U180, P2_ADD_394_U181, P2_ADD_394_U182, P2_ADD_394_U183, P2_ADD_394_U184, P2_ADD_394_U185, P2_ADD_394_U186, P2_R2267_U6, P2_R2267_U7, P2_R2267_U8, P2_R2267_U9, P2_R2267_U10, P2_R2267_U11, P2_R2267_U12, P2_R2267_U13, P2_R2267_U14, P2_R2267_U15, P2_R2267_U16, P2_R2267_U17, P2_R2267_U18, P2_R2267_U19, P2_R2267_U20, P2_R2267_U21, P2_R2267_U22, P2_R2267_U23, P2_R2267_U24, P2_R2267_U25, P2_R2267_U26, P2_R2267_U27, P2_R2267_U28, P2_R2267_U29, P2_R2267_U30, P2_R2267_U31, P2_R2267_U32, P2_R2267_U33, P2_R2267_U34, P2_R2267_U35, P2_R2267_U36, P2_R2267_U37, P2_R2267_U38, P2_R2267_U39, P2_R2267_U40, P2_R2267_U41, P2_R2267_U42, P2_R2267_U43, P2_R2267_U44, P2_R2267_U45, P2_R2267_U46, P2_R2267_U47, P2_R2267_U48, P2_R2267_U49, P2_R2267_U50, P2_R2267_U51, P2_R2267_U52, P2_R2267_U53, P2_R2267_U54, P2_R2267_U55, P2_R2267_U56, P2_R2267_U57, P2_R2267_U58, P2_R2267_U59, P2_R2267_U60, P2_R2267_U61, P2_R2267_U62, P2_R2267_U63, P2_R2267_U64, P2_R2267_U65, P2_R2267_U66, P2_R2267_U67, P2_R2267_U68, P2_R2267_U69, P2_R2267_U70, P2_R2267_U71, P2_R2267_U72, P2_R2267_U73, P2_R2267_U74, P2_R2267_U75, P2_R2267_U76, P2_R2267_U77, P2_R2267_U78, P2_R2267_U79, P2_R2267_U80, P2_R2267_U81, P2_R2267_U82, P2_R2267_U83, P2_R2267_U84, P2_R2267_U85, P2_R2267_U86, P2_R2267_U87, P2_R2267_U88, P2_R2267_U89, P2_R2267_U90, P2_R2267_U91, P2_R2267_U92, P2_R2267_U93, P2_R2267_U94, P2_R2267_U95, P2_R2267_U96, P2_R2267_U97, P2_R2267_U98, P2_R2267_U99, P2_R2267_U100, P2_R2267_U101, P2_R2267_U102, P2_R2267_U103, P2_R2267_U104, P2_R2267_U105, P2_R2267_U106, P2_R2267_U107, P2_R2267_U108, P2_R2267_U109, P2_R2267_U110, P2_R2267_U111, P2_R2267_U112, P2_R2267_U113, P2_R2267_U114, P2_R2267_U115, P2_R2267_U116, P2_R2267_U117, P2_R2267_U118, P2_R2267_U119, P2_R2267_U120, P2_R2267_U121, P2_R2267_U122, P2_R2267_U123, P2_R2267_U124, P2_R2267_U125, P2_R2267_U126, P2_R2267_U127, P2_R2267_U128, P2_R2267_U129, P2_R2267_U130, P2_R2267_U131, P2_R2267_U132, P2_R2267_U133, P2_R2267_U134, P2_R2267_U135, P2_R2267_U136, P2_R2267_U137, P2_R2267_U138, P2_R2267_U139, P2_R2267_U140, P2_R2267_U141, P2_R2267_U142, P2_R2267_U143, P2_R2267_U144, P2_R2267_U145, P2_R2267_U146, P2_R2267_U147, P2_R2267_U148, P2_R2267_U149, P2_R2267_U150, P2_R2267_U151, P2_R2267_U152, P2_R2267_U153, P2_R2267_U154, P2_R2267_U155, P2_R2267_U156, P2_R2267_U157, P2_R2267_U158, P2_R2267_U159, P2_R2267_U160, P2_R2267_U161, P2_R2267_U162, P2_R2267_U163, P2_R2267_U164, P2_R2267_U165, P2_R2267_U166, P2_ADD_371_1212_U4, P2_ADD_371_1212_U5, P2_ADD_371_1212_U6, P2_ADD_371_1212_U7, P2_ADD_371_1212_U8, P2_ADD_371_1212_U9, P2_ADD_371_1212_U10, P2_ADD_371_1212_U11, P2_ADD_371_1212_U12, P2_ADD_371_1212_U13, P2_ADD_371_1212_U14, P2_ADD_371_1212_U15, P2_ADD_371_1212_U16, P2_ADD_371_1212_U17, P2_ADD_371_1212_U18, P2_ADD_371_1212_U19, P2_ADD_371_1212_U20, P2_ADD_371_1212_U21, P2_ADD_371_1212_U22, P2_ADD_371_1212_U23, P2_ADD_371_1212_U24, P2_ADD_371_1212_U25, P2_ADD_371_1212_U26, P2_ADD_371_1212_U27, P2_ADD_371_1212_U28, P2_ADD_371_1212_U29, P2_ADD_371_1212_U30, P2_ADD_371_1212_U31, P2_ADD_371_1212_U32, P2_ADD_371_1212_U33, P2_ADD_371_1212_U34, P2_ADD_371_1212_U35, P2_ADD_371_1212_U36, P2_ADD_371_1212_U37, P2_ADD_371_1212_U38, P2_ADD_371_1212_U39, P2_ADD_371_1212_U40, P2_ADD_371_1212_U41, P2_ADD_371_1212_U42, P2_ADD_371_1212_U43, P2_ADD_371_1212_U44, P2_ADD_371_1212_U45, P2_ADD_371_1212_U46, P2_ADD_371_1212_U47, P2_ADD_371_1212_U48, P2_ADD_371_1212_U49, P2_ADD_371_1212_U50, P2_ADD_371_1212_U51, P2_ADD_371_1212_U52, P2_ADD_371_1212_U53, P2_ADD_371_1212_U54, P2_ADD_371_1212_U55, P2_ADD_371_1212_U56, P2_ADD_371_1212_U57, P2_ADD_371_1212_U58, P2_ADD_371_1212_U59, P2_ADD_371_1212_U60, P2_ADD_371_1212_U61, P2_ADD_371_1212_U62, P2_ADD_371_1212_U63, P2_ADD_371_1212_U64, P2_ADD_371_1212_U65, P2_ADD_371_1212_U66, P2_ADD_371_1212_U67, P2_ADD_371_1212_U68, P2_ADD_371_1212_U69, P2_ADD_371_1212_U70, P2_ADD_371_1212_U71, P2_ADD_371_1212_U72, P2_ADD_371_1212_U73, P2_ADD_371_1212_U74, P2_ADD_371_1212_U75, P2_ADD_371_1212_U76, P2_ADD_371_1212_U77, P2_ADD_371_1212_U78, P2_ADD_371_1212_U79, P2_ADD_371_1212_U80, P2_ADD_371_1212_U81, P2_ADD_371_1212_U82, P2_ADD_371_1212_U83, P2_ADD_371_1212_U84, P2_ADD_371_1212_U85, P2_ADD_371_1212_U86, P2_ADD_371_1212_U87, P2_ADD_371_1212_U88, P2_ADD_371_1212_U89, P2_ADD_371_1212_U90, P2_ADD_371_1212_U91, P2_ADD_371_1212_U92, P2_ADD_371_1212_U93, P2_ADD_371_1212_U94, P2_ADD_371_1212_U95, P2_ADD_371_1212_U96, P2_ADD_371_1212_U97, P2_ADD_371_1212_U98, P2_ADD_371_1212_U99, P2_ADD_371_1212_U100, P2_ADD_371_1212_U101, P2_ADD_371_1212_U102, P2_ADD_371_1212_U103, P2_ADD_371_1212_U104, P2_ADD_371_1212_U105, P2_ADD_371_1212_U106, P2_ADD_371_1212_U107, P2_ADD_371_1212_U108, P2_ADD_371_1212_U109, P2_ADD_371_1212_U110, P2_ADD_371_1212_U111, P2_ADD_371_1212_U112, P2_ADD_371_1212_U113, P2_ADD_371_1212_U114, P2_ADD_371_1212_U115, P2_ADD_371_1212_U116, P2_ADD_371_1212_U117, P2_ADD_371_1212_U118, P2_ADD_371_1212_U119, P2_ADD_371_1212_U120, P2_ADD_371_1212_U121, P2_ADD_371_1212_U122, P2_ADD_371_1212_U123, P2_ADD_371_1212_U124, P2_ADD_371_1212_U125, P2_ADD_371_1212_U126, P2_ADD_371_1212_U127, P2_ADD_371_1212_U128, P2_ADD_371_1212_U129, P2_ADD_371_1212_U130, P2_ADD_371_1212_U131, P2_ADD_371_1212_U132, P2_ADD_371_1212_U133, P2_ADD_371_1212_U134, P2_ADD_371_1212_U135, P2_ADD_371_1212_U136, P2_ADD_371_1212_U137, P2_ADD_371_1212_U138, P2_ADD_371_1212_U139, P2_ADD_371_1212_U140, P2_ADD_371_1212_U141, P2_ADD_371_1212_U142, P2_ADD_371_1212_U143, P2_ADD_371_1212_U144, P2_ADD_371_1212_U145, P2_ADD_371_1212_U146, P2_ADD_371_1212_U147, P2_ADD_371_1212_U148, P2_ADD_371_1212_U149, P2_ADD_371_1212_U150, P2_ADD_371_1212_U151, P2_ADD_371_1212_U152, P2_ADD_371_1212_U153, P2_ADD_371_1212_U154, P2_ADD_371_1212_U155, P2_ADD_371_1212_U156, P2_ADD_371_1212_U157, P2_ADD_371_1212_U158, P2_ADD_371_1212_U159, P2_ADD_371_1212_U160, P2_ADD_371_1212_U161, P2_ADD_371_1212_U162, P2_ADD_371_1212_U163, P2_ADD_371_1212_U164, P2_ADD_371_1212_U165, P2_ADD_371_1212_U166, P2_ADD_371_1212_U167, P2_ADD_371_1212_U168, P2_ADD_371_1212_U169, P2_ADD_371_1212_U170, P2_ADD_371_1212_U171, P2_ADD_371_1212_U172, P2_ADD_371_1212_U173, P2_ADD_371_1212_U174, P2_ADD_371_1212_U175, P2_ADD_371_1212_U176, P2_ADD_371_1212_U177, P2_ADD_371_1212_U178, P2_ADD_371_1212_U179, P2_ADD_371_1212_U180, P2_ADD_371_1212_U181, P2_ADD_371_1212_U182, P2_ADD_371_1212_U183, P2_ADD_371_1212_U184, P2_ADD_371_1212_U185, P2_ADD_371_1212_U186, P2_ADD_371_1212_U187, P2_ADD_371_1212_U188, P2_ADD_371_1212_U189, P2_ADD_371_1212_U190, P2_ADD_371_1212_U191, P2_ADD_371_1212_U192, P2_ADD_371_1212_U193, P2_ADD_371_1212_U194, P2_ADD_371_1212_U195, P2_ADD_371_1212_U196, P2_ADD_371_1212_U197, P2_ADD_371_1212_U198, P2_ADD_371_1212_U199, P2_ADD_371_1212_U200, P2_ADD_371_1212_U201, P2_ADD_371_1212_U202, P2_ADD_371_1212_U203, P2_ADD_371_1212_U204, P2_ADD_371_1212_U205, P2_ADD_371_1212_U206, P2_ADD_371_1212_U207, P2_ADD_371_1212_U208, P2_ADD_371_1212_U209, P2_ADD_371_1212_U210, P2_ADD_371_1212_U211, P2_ADD_371_1212_U212, P2_ADD_371_1212_U213, P2_ADD_371_1212_U214, P2_ADD_371_1212_U215, P2_ADD_371_1212_U216, P2_ADD_371_1212_U217, P2_ADD_371_1212_U218, P2_ADD_371_1212_U219, P2_ADD_371_1212_U220, P2_ADD_371_1212_U221, P2_ADD_371_1212_U222, P2_ADD_371_1212_U223, P2_ADD_371_1212_U224, P2_ADD_371_1212_U225, P2_ADD_371_1212_U226, P2_ADD_371_1212_U227, P2_ADD_371_1212_U228, P2_ADD_371_1212_U229, P2_ADD_371_1212_U230, P2_ADD_371_1212_U231, P2_ADD_371_1212_U232, P2_ADD_371_1212_U233, P2_ADD_371_1212_U234, P2_ADD_371_1212_U235, P2_ADD_371_1212_U236, P2_ADD_371_1212_U237, P2_ADD_371_1212_U238, P2_ADD_371_1212_U239, P2_ADD_371_1212_U240, P2_ADD_371_1212_U241, P2_ADD_371_1212_U242, P2_ADD_371_1212_U243, P2_ADD_371_1212_U244, P2_ADD_371_1212_U245, P2_ADD_371_1212_U246, P2_ADD_371_1212_U247, P2_ADD_371_1212_U248, P2_ADD_371_1212_U249, P2_ADD_371_1212_U250, P2_ADD_371_1212_U251, P2_ADD_371_1212_U252, P2_ADD_371_1212_U253, P2_ADD_371_1212_U254, P2_ADD_371_1212_U255, P2_ADD_371_1212_U256, P2_ADD_371_1212_U257, P2_ADD_371_1212_U258, P2_ADD_371_1212_U259, P2_ADD_371_1212_U260, P2_ADD_371_1212_U261, P2_ADD_371_1212_U262, P2_ADD_371_1212_U263, P2_ADD_371_1212_U264, P2_ADD_371_1212_U265, P2_ADD_371_1212_U266, P2_ADD_371_1212_U267, P2_ADD_371_1212_U268, P2_ADD_371_1212_U269, P2_ADD_371_1212_U270, P2_ADD_371_1212_U271, P2_ADD_371_1212_U272, P2_ADD_371_1212_U273, P2_ADD_371_1212_U274, P2_ADD_371_1212_U275, P2_ADD_371_1212_U276, P2_ADD_371_1212_U277, P2_ADD_371_1212_U278, P2_ADD_371_1212_U279, P2_ADD_371_1212_U280, P2_ADD_371_1212_U281, P2_ADD_371_1212_U282, P1_R2027_U5, P1_R2027_U6, P1_R2027_U7, P1_R2027_U8, P1_R2027_U9, P1_R2027_U10, P1_R2027_U11, P1_R2027_U12, P1_R2027_U13, P1_R2027_U14, P1_R2027_U15, P1_R2027_U16, P1_R2027_U17, P1_R2027_U18, P1_R2027_U19, P1_R2027_U20, P1_R2027_U21, P1_R2027_U22, P1_R2027_U23, P1_R2027_U24, P1_R2027_U25, P1_R2027_U26, P1_R2027_U27, P1_R2027_U28, P1_R2027_U29, P1_R2027_U30, P1_R2027_U31, P1_R2027_U32, P1_R2027_U33, P1_R2027_U34, P1_R2027_U35, P1_R2027_U36, P1_R2027_U37, P1_R2027_U38, P1_R2027_U39, P1_R2027_U40, P1_R2027_U41, P1_R2027_U42, P1_R2027_U43, P1_R2027_U44, P1_R2027_U45, P1_R2027_U46, P1_R2027_U47, P1_R2027_U48, P1_R2027_U49, P1_R2027_U50, P1_R2027_U51, P1_R2027_U52, P1_R2027_U53, P1_R2027_U54, P1_R2027_U55, P1_R2027_U56, P1_R2027_U57, P1_R2027_U58, P1_R2027_U59, P1_R2027_U60, P1_R2027_U61, P1_R2027_U62, P1_R2027_U63, P1_R2027_U64, P1_R2027_U65, P1_R2027_U66, P1_R2027_U67, P1_R2027_U68, P1_R2027_U69, P1_R2027_U70, P1_R2027_U71, P1_R2027_U72, P1_R2027_U73, P1_R2027_U74, P1_R2027_U75, P1_R2027_U76, P1_R2027_U77, P1_R2027_U78, P1_R2027_U79, P1_R2027_U80, P1_R2027_U81, P1_R2027_U82, P1_R2027_U83, P1_R2027_U84, P1_R2027_U85, P1_R2027_U86, P1_R2027_U87, P1_R2027_U88, P1_R2027_U89, P1_R2027_U90, P1_R2027_U91, P1_R2027_U92, P1_R2027_U93, P1_R2027_U94, P1_R2027_U95, P1_R2027_U96, P1_R2027_U97, P1_R2027_U98, P1_R2027_U99, P1_R2027_U100, P1_R2027_U101, P1_R2027_U102, P1_R2027_U103, P1_R2027_U104, P1_R2027_U105, P1_R2027_U106, P1_R2027_U107, P1_R2027_U108, P1_R2027_U109, P1_R2027_U110, P1_R2027_U111, P1_R2027_U112, P1_R2027_U113, P1_R2027_U114, P1_R2027_U115, P1_R2027_U116, P1_R2027_U117, P1_R2027_U118, P1_R2027_U119, P1_R2027_U120, P1_R2027_U121, P1_R2027_U122, P1_R2027_U123, P1_R2027_U124, P1_R2027_U125, P1_R2027_U126, P1_R2027_U127, P1_R2027_U128, P1_R2027_U129, P1_R2027_U130, P1_R2027_U131, P1_R2027_U132, P1_R2027_U133, P1_R2027_U134, P1_R2027_U135, P1_R2027_U136, P1_R2027_U137, P1_R2027_U138, P1_R2027_U139, P1_R2027_U140, P1_R2027_U141, P1_R2027_U142, P1_R2027_U143, P1_R2027_U144, P1_R2027_U145, P1_R2027_U146, P1_R2027_U147, P1_R2027_U148, P1_R2027_U149, P1_R2027_U150, P1_R2027_U151, P1_R2027_U152, P1_R2027_U153, P1_R2027_U154, P1_R2027_U155, P1_R2027_U156, P1_R2027_U157, P1_R2027_U158, P1_R2027_U159, P1_R2027_U160, P1_R2027_U161, P1_R2027_U162, P1_R2027_U163, P1_R2027_U164, P1_R2027_U165, P1_R2027_U166, P1_R2027_U167, P1_R2027_U168, P1_R2027_U169, P1_R2027_U170, P1_R2027_U171, P1_R2027_U172, P1_R2027_U173, P1_R2027_U174, P1_R2027_U175, P1_R2027_U176, P1_R2027_U177, P1_R2027_U178, P1_R2027_U179, P1_R2027_U180, P1_R2027_U181, P1_R2027_U182, P1_R2027_U183, P1_R2027_U184, P1_R2027_U185, P1_R2027_U186, P1_R2027_U187, P1_R2027_U188, P1_R2027_U189, P1_R2027_U190, P1_R2027_U191, P1_R2027_U192, P1_R2027_U193, P1_R2027_U194, P1_R2027_U195, P1_R2027_U196, P1_R2027_U197, P1_R2027_U198, P1_R2027_U199, P1_R2027_U200, P1_R2027_U201, P1_R2027_U202, P1_R2182_U5, P1_R2182_U6, P1_R2182_U7, P1_R2182_U8, P1_R2182_U9, P1_R2182_U10, P1_R2182_U11, P1_R2182_U12, P1_R2182_U13, P1_R2182_U14, P1_R2182_U15, P1_R2182_U16, P1_R2182_U17, P1_R2182_U18, P1_R2182_U19, P1_R2182_U20, P1_R2182_U21, P1_R2182_U22, P1_R2182_U23, P1_R2182_U24, P1_R2182_U25, P1_R2182_U26, P1_R2182_U27, P1_R2182_U28, P1_R2182_U29, P1_R2182_U30, P1_R2182_U31, P1_R2182_U32, P1_R2182_U33, P1_R2182_U34, P1_R2182_U35, P1_R2182_U36, P1_R2182_U37, P1_R2182_U38, P1_R2182_U39, P1_R2182_U40, P1_R2182_U41, P1_R2182_U42, P1_R2182_U43, P1_R2182_U44, P1_R2182_U45, P1_R2182_U46, P1_R2182_U47, P1_R2182_U48, P1_R2182_U49, P1_R2182_U50, P1_R2182_U51, P1_R2182_U52, P1_R2182_U53, P1_R2182_U54, P1_R2182_U55, P1_R2182_U56, P1_R2182_U57, P1_R2182_U58, P1_R2182_U59, P1_R2182_U60, P1_R2182_U61, P1_R2182_U62, P1_R2182_U63, P1_R2182_U64, P1_R2182_U65, P1_R2182_U66, P1_R2182_U67, P1_R2182_U68, P1_R2182_U69, P1_R2182_U70, P1_R2182_U71, P1_R2182_U72, P1_R2182_U73, P1_R2182_U74, P1_R2182_U75, P1_R2182_U76, P1_R2182_U77, P1_R2182_U78, P1_R2182_U79, P1_R2182_U80, P1_R2182_U81, P1_R2182_U82, P1_R2182_U83, P1_R2182_U84, P1_R2182_U85, P1_R2182_U86, P1_R2144_U5, P1_R2144_U6, P1_R2144_U7, P1_R2144_U8, P1_R2144_U9, P1_R2144_U10, P1_R2144_U11, P1_R2144_U12, P1_R2144_U13, P1_R2144_U14, P1_R2144_U15, P1_R2144_U16, P1_R2144_U17, P1_R2144_U18, P1_R2144_U19, P1_R2144_U20, P1_R2144_U21, P1_R2144_U22, P1_R2144_U23, P1_R2144_U24, P1_R2144_U25, P1_R2144_U26, P1_R2144_U27, P1_R2144_U28, P1_R2144_U29, P1_R2144_U30, P1_R2144_U31, P1_R2144_U32, P1_R2144_U33, P1_R2144_U34, P1_R2144_U35, P1_R2144_U36, P1_R2144_U37, P1_R2144_U38, P1_R2144_U39, P1_R2144_U40, P1_R2144_U41, P1_R2144_U42, P1_R2144_U43, P1_R2144_U44, P1_R2144_U45, P1_R2144_U46, P1_R2144_U47, P1_R2144_U48, P1_R2144_U49, P1_R2144_U50, P1_R2144_U51, P1_R2144_U52, P1_R2144_U53, P1_R2144_U54, P1_R2144_U55, P1_R2144_U56, P1_R2144_U57, P1_R2144_U58, P1_R2144_U59, P1_R2144_U60, P1_R2144_U61, P1_R2144_U62, P1_R2144_U63, P1_R2144_U64, P1_R2144_U65, P1_R2144_U66, P1_R2144_U67, P1_R2144_U68, P1_R2144_U69, P1_R2144_U70, P1_R2144_U71, P1_R2144_U72, P1_R2144_U73, P1_R2144_U74, P1_R2144_U75, P1_R2144_U76, P1_R2144_U77, P1_R2144_U78, P1_R2144_U79, P1_R2144_U80, P1_R2144_U81, P1_R2144_U82, P1_R2144_U83, P1_R2144_U84, P1_R2144_U85, P1_R2144_U86, P1_R2144_U87, P1_R2144_U88, P1_R2144_U89, P1_R2144_U90, P1_R2144_U91, P1_R2144_U92, P1_R2144_U93, P1_R2144_U94, P1_R2144_U95, P1_R2144_U96, P1_R2144_U97, P1_R2144_U98, P1_R2144_U99, P1_R2144_U100, P1_R2144_U101, P1_R2144_U102, P1_R2144_U103, P1_R2144_U104, P1_R2144_U105, P1_R2144_U106, P1_R2144_U107, P1_R2144_U108, P1_R2144_U109, P1_R2144_U110, P1_R2144_U111, P1_R2144_U112, P1_R2144_U113, P1_R2144_U114, P1_R2144_U115, P1_R2144_U116, P1_R2144_U117, P1_R2144_U118, P1_R2144_U119, P1_R2144_U120, P1_R2144_U121, P1_R2144_U122, P1_R2144_U123, P1_R2144_U124, P1_R2144_U125, P1_R2144_U126, P1_R2144_U127, P1_R2144_U128, P1_R2144_U129, P1_R2144_U130, P1_R2144_U131, P1_R2144_U132, P1_R2144_U133, P1_R2144_U134, P1_R2144_U135, P1_R2144_U136, P1_R2144_U137, P1_R2144_U138, P1_R2144_U139, P1_R2144_U140, P1_R2144_U141, P1_R2144_U142, P1_R2144_U143, P1_R2144_U144, P1_R2144_U145, P1_R2144_U146, P1_R2144_U147, P1_R2144_U148, P1_R2144_U149, P1_R2144_U150, P1_R2144_U151, P1_R2144_U152, P1_R2144_U153, P1_R2144_U154, P1_R2144_U155, P1_R2144_U156, P1_R2144_U157, P1_R2144_U158, P1_R2144_U159, P1_R2144_U160, P1_R2144_U161, P1_R2144_U162, P1_R2144_U163, P1_R2144_U164, P1_R2144_U165, P1_R2144_U166, P1_R2144_U167, P1_R2144_U168, P1_R2144_U169, P1_R2144_U170, P1_R2144_U171, P1_R2144_U172, P1_R2144_U173, P1_R2144_U174, P1_R2144_U175, P1_R2144_U176, P1_R2144_U177, P1_R2144_U178, P1_R2144_U179, P1_R2144_U180, P1_R2144_U181, P1_R2144_U182, P1_R2144_U183, P1_R2144_U184, P1_R2144_U185, P1_R2144_U186, P1_R2144_U187, P1_R2144_U188, P1_R2144_U189, P1_R2144_U190, P1_R2144_U191, P1_R2144_U192, P1_R2144_U193, P1_R2144_U194, P1_R2144_U195, P1_R2144_U196, P1_R2144_U197, P1_R2144_U198, P1_R2144_U199, P1_R2144_U200, P1_R2144_U201, P1_R2144_U202, P1_R2144_U203, P1_R2144_U204, P1_R2144_U205, P1_R2144_U206, P1_R2144_U207, P1_R2144_U208, P1_R2144_U209, P1_R2144_U210, P1_R2144_U211, P1_R2144_U212, P1_R2144_U213, P1_R2144_U214, P1_R2144_U215, P1_R2144_U216, P1_R2144_U217, P1_R2144_U218, P1_R2144_U219, P1_R2144_U220, P1_R2144_U221, P1_R2144_U222, P1_R2144_U223, P1_R2144_U224, P1_R2144_U225, P1_R2144_U226, P1_R2144_U227, P1_R2144_U228, P1_R2144_U229, P1_R2144_U230, P1_R2144_U231, P1_R2144_U232, P1_R2144_U233, P1_R2144_U234, P1_R2144_U235, P1_R2144_U236, P1_R2144_U237, P1_R2144_U238, P1_R2144_U239, P1_R2144_U240, P1_R2144_U241, P1_R2144_U242, P1_R2144_U243, P1_R2144_U244, P1_R2144_U245, P1_R2144_U246, P1_R2144_U247, P1_R2144_U248, P1_R2144_U249, P1_R2144_U250, P1_R2144_U251, P1_R2144_U252, P1_R2144_U253, P1_R2144_U254, P1_R2144_U255, P1_R2144_U256, P1_R2144_U257, P1_R2144_U258, P1_R2144_U259, P1_R2144_U260, P1_R2278_U5, P1_R2278_U6, P1_R2278_U7, P1_R2278_U8, P1_R2278_U9, P1_R2278_U10, P1_R2278_U11, P1_R2278_U12, P1_R2278_U13, P1_R2278_U14, P1_R2278_U15, P1_R2278_U16, P1_R2278_U17, P1_R2278_U18, P1_R2278_U19, P1_R2278_U20, P1_R2278_U21, P1_R2278_U22, P1_R2278_U23, P1_R2278_U24, P1_R2278_U25, P1_R2278_U26, P1_R2278_U27, P1_R2278_U28, P1_R2278_U29, P1_R2278_U30, P1_R2278_U31, P1_R2278_U32, P1_R2278_U33, P1_R2278_U34, P1_R2278_U35, P1_R2278_U36, P1_R2278_U37, P1_R2278_U38, P1_R2278_U39, P1_R2278_U40, P1_R2278_U41, P1_R2278_U42, P1_R2278_U43, P1_R2278_U44, P1_R2278_U45, P1_R2278_U46, P1_R2278_U47, P1_R2278_U48, P1_R2278_U49, P1_R2278_U50, P1_R2278_U51, P1_R2278_U52, P1_R2278_U53, P1_R2278_U54, P1_R2278_U55, P1_R2278_U56, P1_R2278_U57, P1_R2278_U58, P1_R2278_U59, P1_R2278_U60, P1_R2278_U61, P1_R2278_U62, P1_R2278_U63, P1_R2278_U64, P1_R2278_U65, P1_R2278_U66, P1_R2278_U67, P1_R2278_U68, P1_R2278_U69, P1_R2278_U70, P1_R2278_U71, P1_R2278_U72, P1_R2278_U73, P1_R2278_U74, P1_R2278_U75, P1_R2278_U76, P1_R2278_U77, P1_R2278_U78, P1_R2278_U79, P1_R2278_U80, P1_R2278_U81, P1_R2278_U82, P1_R2278_U83, P1_R2278_U84, P1_R2278_U85, P1_R2278_U86, P1_R2278_U87, P1_R2278_U88, P1_R2278_U89, P1_R2278_U90, P1_R2278_U91, P1_R2278_U92, P1_R2278_U93, P1_R2278_U94, P1_R2278_U95, P1_R2278_U96, P1_R2278_U97, P1_R2278_U98, P1_R2278_U99, P1_R2278_U100, P1_R2278_U101, P1_R2278_U102, P1_R2278_U103, P1_R2278_U104, P1_R2278_U105, P1_R2278_U106, P1_R2278_U107, P1_R2278_U108, P1_R2278_U109, P1_R2278_U110, P1_R2278_U111, P1_R2278_U112, P1_R2278_U113, P1_R2278_U114, P1_R2278_U115, P1_R2278_U116, P1_R2278_U117, P1_R2278_U118, P1_R2278_U119, P1_R2278_U120, P1_R2278_U121, P1_R2278_U122, P1_R2278_U123, P1_R2278_U124, P1_R2278_U125, P1_R2278_U126, P1_R2278_U127, P1_R2278_U128, P1_R2278_U129, P1_R2278_U130, P1_R2278_U131, P1_R2278_U132, P1_R2278_U133, P1_R2278_U134, P1_R2278_U135, P1_R2278_U136, P1_R2278_U137, P1_R2278_U138, P1_R2278_U139, P1_R2278_U140, P1_R2278_U141, P1_R2278_U142, P1_R2278_U143, P1_R2278_U144, P1_R2278_U145, P1_R2278_U146, P1_R2278_U147, P1_R2278_U148, P1_R2278_U149, P1_R2278_U150, P1_R2278_U151, P1_R2278_U152, P1_R2278_U153, P1_R2278_U154, P1_R2278_U155, P1_R2278_U156, P1_R2278_U157, P1_R2278_U158, P1_R2278_U159, P1_R2278_U160, P1_R2278_U161, P1_R2278_U162, P1_R2278_U163, P1_R2278_U164, P1_R2278_U165, P1_R2278_U166, P1_R2278_U167, P1_R2278_U168, P1_R2278_U169, P1_R2278_U170, P1_R2278_U171, P1_R2278_U172, P1_R2278_U173, P1_R2278_U174, P1_R2278_U175, P1_R2278_U176, P1_R2278_U177, P1_R2278_U178, P1_R2278_U179, P1_R2278_U180, P1_R2278_U181, P1_R2278_U182, P1_R2278_U183, P1_R2278_U184, P1_R2278_U185, P1_R2278_U186, P1_R2278_U187, P1_R2278_U188, P1_R2278_U189, P1_R2278_U190, P1_R2278_U191, P1_R2278_U192, P1_R2278_U193, P1_R2278_U194, P1_R2278_U195, P1_R2278_U196, P1_R2278_U197, P1_R2278_U198, P1_R2278_U199, P1_R2278_U200, P1_R2278_U201, P1_R2278_U202, P1_R2278_U203, P1_R2278_U204, P1_R2278_U205, P1_R2278_U206, P1_R2278_U207, P1_R2278_U208, P1_R2278_U209, P1_R2278_U210, P1_R2278_U211, P1_R2278_U212, P1_R2278_U213, P1_R2278_U214, P1_R2278_U215, P1_R2278_U216, P1_R2278_U217, P1_R2278_U218, P1_R2278_U219, P1_R2278_U220, P1_R2278_U221, P1_R2278_U222, P1_R2278_U223, P1_R2278_U224, P1_R2278_U225, P1_R2278_U226, P1_R2278_U227, P1_R2278_U228, P1_R2278_U229, P1_R2278_U230, P1_R2278_U231, P1_R2278_U232, P1_R2278_U233, P1_R2278_U234, P1_R2278_U235, P1_R2278_U236, P1_R2278_U237, P1_R2278_U238, P1_R2278_U239, P1_R2278_U240, P1_R2278_U241, P1_R2278_U242, P1_R2278_U243, P1_R2278_U244, P1_R2278_U245, P1_R2278_U246, P1_R2278_U247, P1_R2278_U248, P1_R2278_U249, P1_R2278_U250, P1_R2278_U251, P1_R2278_U252, P1_R2278_U253, P1_R2278_U254, P1_R2278_U255, P1_R2278_U256, P1_R2278_U257, P1_R2278_U258, P1_R2278_U259, P1_R2278_U260, P1_R2278_U261, P1_R2278_U262, P1_R2278_U263, P1_R2278_U264, P1_R2278_U265, P1_R2278_U266, P1_R2278_U267, P1_R2278_U268, P1_R2278_U269, P1_R2278_U270, P1_R2278_U271, P1_R2278_U272, P1_R2278_U273, P1_R2278_U274, P1_R2278_U275, P1_R2278_U276, P1_R2278_U277, P1_R2278_U278, P1_R2278_U279, P1_R2278_U280, P1_R2278_U281, P1_R2278_U282, P1_R2278_U283, P1_R2278_U284, P1_R2278_U285, P1_R2278_U286, P1_R2278_U287, P1_R2278_U288, P1_R2278_U289, P1_R2278_U290, P1_R2278_U291, P1_R2278_U292, P1_R2278_U293, P1_R2278_U294, P1_R2278_U295, P1_R2278_U296, P1_R2278_U297, P1_R2278_U298, P1_R2278_U299, P1_R2278_U300, P1_R2278_U301, P1_R2278_U302, P1_R2278_U303, P1_R2278_U304, P1_R2278_U305, P1_R2278_U306, P1_R2278_U307, P1_R2278_U308, P1_R2278_U309, P1_R2278_U310, P1_R2278_U311, P1_R2278_U312, P1_R2278_U313, P1_R2278_U314, P1_R2278_U315, P1_R2278_U316, P1_R2278_U317, P1_R2278_U318, P1_R2278_U319, P1_R2278_U320, P1_R2278_U321, P1_R2278_U322, P1_R2278_U323, P1_R2278_U324, P1_R2278_U325, P1_R2278_U326, P1_R2278_U327, P1_R2278_U328, P1_R2278_U329, P1_R2278_U330, P1_R2278_U331, P1_R2278_U332, P1_R2278_U333, P1_R2278_U334, P1_R2278_U335, P1_R2278_U336, P1_R2278_U337, P1_R2278_U338, P1_R2278_U339, P1_R2278_U340, P1_R2278_U341, P1_R2278_U342, P1_R2278_U343, P1_R2278_U344, P1_R2278_U345, P1_R2278_U346, P1_R2278_U347, P1_R2278_U348, P1_R2278_U349, P1_R2278_U350, P1_R2278_U351, P1_R2278_U352, P1_R2278_U353, P1_R2278_U354, P1_R2278_U355, P1_R2278_U356, P1_R2278_U357, P1_R2278_U358, P1_R2278_U359, P1_R2278_U360, P1_R2278_U361, P1_R2278_U362, P1_R2278_U363, P1_R2278_U364, P1_R2278_U365, P1_R2278_U366, P1_R2278_U367, P1_R2278_U368, P1_R2278_U369, P1_R2278_U370, P1_R2278_U371, P1_R2278_U372, P1_R2278_U373, P1_R2278_U374, P1_R2278_U375, P1_R2278_U376, P1_R2278_U377, P1_R2278_U378, P1_R2278_U379, P1_R2278_U380, P1_R2278_U381, P1_R2278_U382, P1_R2278_U383, P1_R2278_U384, P1_R2278_U385, P1_R2278_U386, P1_R2278_U387, P1_R2278_U388, P1_R2278_U389, P1_R2278_U390, P1_R2278_U391, P1_R2278_U392, P1_R2278_U393, P1_R2278_U394, P1_R2278_U395, P1_R2278_U396, P1_R2278_U397, P1_R2278_U398, P1_R2278_U399, P1_R2278_U400, P1_R2278_U401, P1_R2278_U402, P1_R2278_U403, P1_R2278_U404, P1_R2278_U405, P1_R2278_U406, P1_R2278_U407, P1_R2278_U408, P1_R2278_U409, P1_R2278_U410, P1_R2278_U411, P1_R2278_U412, P1_R2278_U413, P1_R2278_U414, P1_R2278_U415, P1_R2278_U416, P1_R2278_U417, P1_R2278_U418, P1_R2278_U419, P1_R2278_U420, P1_R2278_U421, P1_R2278_U422, P1_R2278_U423, P1_R2278_U424, P1_R2278_U425, P1_R2278_U426, P1_R2278_U427, P1_R2278_U428, P1_R2278_U429, P1_R2278_U430, P1_R2278_U431, P1_R2278_U432, P1_R2278_U433, P1_R2278_U434, P1_R2278_U435, P1_R2278_U436, P1_R2278_U437, P1_R2278_U438, P1_R2278_U439, P1_R2278_U440, P1_R2278_U441, P1_R2278_U442, P1_R2278_U443, P1_R2278_U444, P1_R2278_U445, P1_R2278_U446, P1_R2278_U447, P1_R2278_U448, P1_R2278_U449, P1_R2278_U450, P1_R2278_U451, P1_R2278_U452, P1_R2278_U453, P1_R2278_U454, P1_R2278_U455, P1_R2278_U456, P1_R2278_U457, P1_R2278_U458, P1_R2278_U459, P1_R2278_U460, P1_R2278_U461, P1_R2278_U462, P1_R2278_U463, P1_R2278_U464, P1_R2278_U465, P1_R2278_U466, P1_R2278_U467, P1_R2278_U468, P1_R2278_U469, P1_R2278_U470, P1_R2278_U471, P1_R2278_U472, P1_R2278_U473, P1_R2278_U474, P1_R2278_U475, P1_R2278_U476, P1_R2278_U477, P1_R2278_U478, P1_R2278_U479, P1_R2278_U480, P1_R2278_U481, P1_R2278_U482, P1_R2278_U483, P1_R2278_U484, P1_R2278_U485, P1_R2278_U486, P1_R2278_U487, P1_R2278_U488, P1_R2278_U489, P1_R2278_U490, P1_R2278_U491, P1_R2278_U492, P1_R2278_U493, P1_R2278_U494, P1_R2278_U495, P1_R2278_U496, P1_R2278_U497, P1_R2278_U498, P1_R2278_U499, P1_R2278_U500, P1_R2278_U501, P1_R2278_U502, P1_R2278_U503, P1_R2278_U504, P1_R2278_U505, P1_R2278_U506, P1_R2278_U507, P1_R2278_U508, P1_R2278_U509, P1_R2278_U510, P1_R2278_U511, P1_R2278_U512, P1_R2278_U513, P1_R2278_U514, P1_R2278_U515, P1_R2278_U516, P1_R2278_U517, P1_R2278_U518, P1_R2278_U519, P1_R2278_U520, P1_R2278_U521, P1_R2278_U522, P1_R2278_U523, P1_R2278_U524, P1_R2278_U525, P1_R2278_U526, P1_R2278_U527, P1_R2278_U528, P1_R2278_U529, P1_R2278_U530, P1_R2278_U531, P1_R2278_U532, P1_R2278_U533, P1_R2278_U534, P1_R2278_U535, P1_R2278_U536, P1_R2278_U537, P1_R2278_U538, P1_R2278_U539, P1_R2278_U540, P1_R2278_U541, P1_R2278_U542, P1_R2278_U543, P1_R2278_U544, P1_R2278_U545, P1_R2278_U546, P1_R2278_U547, P1_R2278_U548, P1_R2278_U549, P1_R2278_U550, P1_R2278_U551, P1_R2278_U552, P1_R2278_U553, P1_R2278_U554, P1_R2278_U555, P1_R2278_U556, P1_R2278_U557, P1_R2278_U558, P1_R2278_U559, P1_R2278_U560, P1_R2278_U561, P1_R2278_U562, P1_R2278_U563, P1_R2278_U564, P1_R2278_U565, P1_R2278_U566, P1_R2278_U567, P1_R2278_U568, P1_R2278_U569, P1_R2278_U570, P1_R2278_U571, P1_R2278_U572, P1_R2278_U573, P1_R2278_U574, P1_R2278_U575, P1_R2278_U576, P1_R2278_U577, P1_R2278_U578, P1_R2278_U579, P1_R2278_U580, P1_R2278_U581, P1_R2278_U582, P1_R2278_U583, P1_R2278_U584, P1_R2278_U585, P1_R2278_U586, P1_R2278_U587, P1_R2278_U588, P1_R2278_U589, P1_R2278_U590, P1_R2278_U591, P1_R2278_U592, P1_R2278_U593, P1_R2278_U594, P1_R2278_U595, P1_R2278_U596, P1_R2278_U597, P1_R2278_U598, P1_R2278_U599, P1_R2278_U600, P1_R2278_U601, P1_R2278_U602, P1_R2278_U603, P1_R2278_U604, P1_R2278_U605, P1_R2278_U606, P1_R2278_U607, P1_R2278_U608, P1_R2278_U609, P1_R2278_U610, P1_R2358_U5, P1_R2358_U6, P1_R2358_U7, P1_R2358_U8, P1_R2358_U9, P1_R2358_U10, P1_R2358_U11, P1_R2358_U12, P1_R2358_U13, P1_R2358_U14, P1_R2358_U15, P1_R2358_U16, P1_R2358_U17, P1_R2358_U18, P1_R2358_U19, P1_R2358_U20, P1_R2358_U21, P1_R2358_U22, P1_R2358_U23, P1_R2358_U24, P1_R2358_U25, P1_R2358_U26, P1_R2358_U27, P1_R2358_U28, P1_R2358_U29, P1_R2358_U30, P1_R2358_U31, P1_R2358_U32, P1_R2358_U33, P1_R2358_U34, P1_R2358_U35, P1_R2358_U36, P1_R2358_U37, P1_R2358_U38, P1_R2358_U39, P1_R2358_U40, P1_R2358_U41, P1_R2358_U42, P1_R2358_U43, P1_R2358_U44, P1_R2358_U45, P1_R2358_U46, P1_R2358_U47, P1_R2358_U48, P1_R2358_U49, P1_R2358_U50, P1_R2358_U51, P1_R2358_U52, P1_R2358_U53, P1_R2358_U54, P1_R2358_U55, P1_R2358_U56, P1_R2358_U57, P1_R2358_U58, P1_R2358_U59, P1_R2358_U60, P1_R2358_U61, P1_R2358_U62, P1_R2358_U63, P1_R2358_U64, P1_R2358_U65, P1_R2358_U66, P1_R2358_U67, P1_R2358_U68, P1_R2358_U69, P1_R2358_U70, P1_R2358_U71, P1_R2358_U72, P1_R2358_U73, P1_R2358_U74, P1_R2358_U75, P1_R2358_U76, P1_R2358_U77, P1_R2358_U78, P1_R2358_U79, P1_R2358_U80, P1_R2358_U81, P1_R2358_U82, P1_R2358_U83, P1_R2358_U84, P1_R2358_U85, P1_R2358_U86, P1_R2358_U87, P1_R2358_U88, P1_R2358_U89, P1_R2358_U90, P1_R2358_U91, P1_R2358_U92, P1_R2358_U93, P1_R2358_U94, P1_R2358_U95, P1_R2358_U96, P1_R2358_U97, P1_R2358_U98, P1_R2358_U99, P1_R2358_U100, P1_R2358_U101, P1_R2358_U102, P1_R2358_U103, P1_R2358_U104, P1_R2358_U105, P1_R2358_U106, P1_R2358_U107, P1_R2358_U108, P1_R2358_U109, P1_R2358_U110, P1_R2358_U111, P1_R2358_U112, P1_R2358_U113, P1_R2358_U114, P1_R2358_U115, P1_R2358_U116, P1_R2358_U117, P1_R2358_U118, P1_R2358_U119, P1_R2358_U120, P1_R2358_U121, P1_R2358_U122, P1_R2358_U123, P1_R2358_U124, P1_R2358_U125, P1_R2358_U126, P1_R2358_U127, P1_R2358_U128, P1_R2358_U129, P1_R2358_U130, P1_R2358_U131, P1_R2358_U132, P1_R2358_U133, P1_R2358_U134, P1_R2358_U135, P1_R2358_U136, P1_R2358_U137, P1_R2358_U138, P1_R2358_U139, P1_R2358_U140, P1_R2358_U141, P1_R2358_U142, P1_R2358_U143, P1_R2358_U144, P1_R2358_U145, P1_R2358_U146, P1_R2358_U147, P1_R2358_U148, P1_R2358_U149, P1_R2358_U150, P1_R2358_U151, P1_R2358_U152, P1_R2358_U153, P1_R2358_U154, P1_R2358_U155, P1_R2358_U156, P1_R2358_U157, P1_R2358_U158, P1_R2358_U159, P1_R2358_U160, P1_R2358_U161, P1_R2358_U162, P1_R2358_U163, P1_R2358_U164, P1_R2358_U165, P1_R2358_U166, P1_R2358_U167, P1_R2358_U168, P1_R2358_U169, P1_R2358_U170, P1_R2358_U171, P1_R2358_U172, P1_R2358_U173, P1_R2358_U174, P1_R2358_U175, P1_R2358_U176, P1_R2358_U177, P1_R2358_U178, P1_R2358_U179, P1_R2358_U180, P1_R2358_U181, P1_R2358_U182, P1_R2358_U183, P1_R2358_U184, P1_R2358_U185, P1_R2358_U186, P1_R2358_U187, P1_R2358_U188, P1_R2358_U189, P1_R2358_U190, P1_R2358_U191, P1_R2358_U192, P1_R2358_U193, P1_R2358_U194, P1_R2358_U195, P1_R2358_U196, P1_R2358_U197, P1_R2358_U198, P1_R2358_U199, P1_R2358_U200, P1_R2358_U201, P1_R2358_U202, P1_R2358_U203, P1_R2358_U204, P1_R2358_U205, P1_R2358_U206, P1_R2358_U207, P1_R2358_U208, P1_R2358_U209, P1_R2358_U210, P1_R2358_U211, P1_R2358_U212, P1_R2358_U213, P1_R2358_U214, P1_R2358_U215, P1_R2358_U216, P1_R2358_U217, P1_R2358_U218, P1_R2358_U219, P1_R2358_U220, P1_R2358_U221, P1_R2358_U222, P1_R2358_U223, P1_R2358_U224, P1_R2358_U225, P1_R2358_U226, P1_R2358_U227, P1_R2358_U228, P1_R2358_U229, P1_R2358_U230, P1_R2358_U231, P1_R2358_U232, P1_R2358_U233, P1_R2358_U234, P1_R2358_U235, P1_R2358_U236, P1_R2358_U237, P1_R2358_U238, P1_R2358_U239, P1_R2358_U240, P1_R2358_U241, P1_R2358_U242, P1_R2358_U243, P1_R2358_U244, P1_R2358_U245, P1_R2358_U246, P1_R2358_U247, P1_R2358_U248, P1_R2358_U249, P1_R2358_U250, P1_R2358_U251, P1_R2358_U252, P1_R2358_U253, P1_R2358_U254, P1_R2358_U255, P1_R2358_U256, P1_R2358_U257, P1_R2358_U258, P1_R2358_U259, P1_R2358_U260, P1_R2358_U261, P1_R2358_U262, P1_R2358_U263, P1_R2358_U264, P1_R2358_U265, P1_R2358_U266, P1_R2358_U267, P1_R2358_U268, P1_R2358_U269, P1_R2358_U270, P1_R2358_U271, P1_R2358_U272, P1_R2358_U273, P1_R2358_U274, P1_R2358_U275, P1_R2358_U276, P1_R2358_U277, P1_R2358_U278, P1_R2358_U279, P1_R2358_U280, P1_R2358_U281, P1_R2358_U282, P1_R2358_U283, P1_R2358_U284, P1_R2358_U285, P1_R2358_U286, P1_R2358_U287, P1_R2358_U288, P1_R2358_U289, P1_R2358_U290, P1_R2358_U291, P1_R2358_U292, P1_R2358_U293, P1_R2358_U294, P1_R2358_U295, P1_R2358_U296, P1_R2358_U297, P1_R2358_U298, P1_R2358_U299, P1_R2358_U300, P1_R2358_U301, P1_R2358_U302, P1_R2358_U303, P1_R2358_U304, P1_R2358_U305, P1_R2358_U306, P1_R2358_U307, P1_R2358_U308, P1_R2358_U309, P1_R2358_U310, P1_R2358_U311, P1_R2358_U312, P1_R2358_U313, P1_R2358_U314, P1_R2358_U315, P1_R2358_U316, P1_R2358_U317, P1_R2358_U318, P1_R2358_U319, P1_R2358_U320, P1_R2358_U321, P1_R2358_U322, P1_R2358_U323, P1_R2358_U324, P1_R2358_U325, P1_R2358_U326, P1_R2358_U327, P1_R2358_U328, P1_R2358_U329, P1_R2358_U330, P1_R2358_U331, P1_R2358_U332, P1_R2358_U333, P1_R2358_U334, P1_R2358_U335, P1_R2358_U336, P1_R2358_U337, P1_R2358_U338, P1_R2358_U339, P1_R2358_U340, P1_R2358_U341, P1_R2358_U342, P1_R2358_U343, P1_R2358_U344, P1_R2358_U345, P1_R2358_U346, P1_R2358_U347, P1_R2358_U348, P1_R2358_U349, P1_R2358_U350, P1_R2358_U351, P1_R2358_U352, P1_R2358_U353, P1_R2358_U354, P1_R2358_U355, P1_R2358_U356, P1_R2358_U357, P1_R2358_U358, P1_R2358_U359, P1_R2358_U360, P1_R2358_U361, P1_R2358_U362, P1_R2358_U363, P1_R2358_U364, P1_R2358_U365, P1_R2358_U366, P1_R2358_U367, P1_R2358_U368, P1_R2358_U369, P1_R2358_U370, P1_R2358_U371, P1_R2358_U372, P1_R2358_U373, P1_R2358_U374, P1_R2358_U375, P1_R2358_U376, P1_R2358_U377, P1_R2358_U378, P1_R2358_U379, P1_R2358_U380, P1_R2358_U381, P1_R2358_U382, P1_R2358_U383, P1_R2358_U384, P1_R2358_U385, P1_R2358_U386, P1_R2358_U387, P1_R2358_U388, P1_R2358_U389, P1_R2358_U390, P1_R2358_U391, P1_R2358_U392, P1_R2358_U393, P1_R2358_U394, P1_R2358_U395, P1_R2358_U396, P1_R2358_U397, P1_R2358_U398, P1_R2358_U399, P1_R2358_U400, P1_R2358_U401, P1_R2358_U402, P1_R2358_U403, P1_R2358_U404, P1_R2358_U405, P1_R2358_U406, P1_R2358_U407, P1_R2358_U408, P1_R2358_U409, P1_R2358_U410, P1_R2358_U411, P1_R2358_U412, P1_R2358_U413, P1_R2358_U414, P1_R2358_U415, P1_R2358_U416, P1_R2358_U417, P1_R2358_U418, P1_R2358_U419, P1_R2358_U420, P1_R2358_U421, P1_R2358_U422, P1_R2358_U423, P1_R2358_U424, P1_R2358_U425, P1_R2358_U426, P1_R2358_U427, P1_R2358_U428, P1_R2358_U429, P1_R2358_U430, P1_R2358_U431, P1_R2358_U432, P1_R2358_U433, P1_R2358_U434, P1_R2358_U435, P1_R2358_U436, P1_R2358_U437, P1_R2358_U438, P1_R2358_U439, P1_R2358_U440, P1_R2358_U441, P1_R2358_U442, P1_R2358_U443, P1_R2358_U444, P1_R2358_U445, P1_R2358_U446, P1_R2358_U447, P1_R2358_U448, P1_R2358_U449, P1_R2358_U450, P1_R2358_U451, P1_R2358_U452, P1_R2358_U453, P1_R2358_U454, P1_R2358_U455, P1_R2358_U456, P1_R2358_U457, P1_R2358_U458, P1_R2358_U459, P1_R2358_U460, P1_R2358_U461, P1_R2358_U462, P1_R2358_U463, P1_R2358_U464, P1_R2358_U465, P1_R2358_U466, P1_R2358_U467, P1_R2358_U468, P1_R2358_U469, P1_R2358_U470, P1_R2358_U471, P1_R2358_U472, P1_R2358_U473, P1_R2358_U474, P1_R2358_U475, P1_R2358_U476, P1_R2358_U477, P1_R2358_U478, P1_R2358_U479, P1_R2358_U480, P1_R2358_U481, P1_R2358_U482, P1_R2358_U483, P1_R2358_U484, P1_R2358_U485, P1_R2358_U486, P1_R2358_U487, P1_R2358_U488, P1_R2358_U489, P1_R2358_U490, P1_R2358_U491, P1_R2358_U492, P1_R2358_U493, P1_R2358_U494, P1_R2358_U495, P1_R2358_U496, P1_R2358_U497, P1_R2358_U498, P1_R2358_U499, P1_R2358_U500, P1_R2358_U501, P1_R2358_U502, P1_R2358_U503, P1_R2358_U504, P1_R2358_U505, P1_R2358_U506, P1_R2358_U507, P1_R2358_U508, P1_R2358_U509, P1_R2358_U510, P1_R2358_U511, P1_R2358_U512, P1_R2358_U513, P1_R2358_U514, P1_R2358_U515, P1_R2358_U516, P1_R2358_U517, P1_R2358_U518, P1_R2358_U519, P1_R2358_U520, P1_R2358_U521, P1_R2358_U522, P1_R2358_U523, P1_R2358_U524, P1_R2358_U525, P1_R2358_U526, P1_R2358_U527, P1_R2358_U528, P1_R2358_U529, P1_R2358_U530, P1_R2358_U531, P1_R2358_U532, P1_R2358_U533, P1_R2358_U534, P1_R2358_U535, P1_R2358_U536, P1_R2358_U537, P1_R2358_U538, P1_R2358_U539, P1_R2358_U540, P1_R2358_U541, P1_R2358_U542, P1_R2358_U543, P1_R2358_U544, P1_R2358_U545, P1_R2358_U546, P1_R2358_U547, P1_R2358_U548, P1_R2358_U549, P1_R2358_U550, P1_R2358_U551, P1_R2358_U552, P1_R2358_U553, P1_R2358_U554, P1_R2358_U555, P1_R2358_U556, P1_R2358_U557, P1_R2358_U558, P1_R2358_U559, P1_R2358_U560, P1_R2358_U561, P1_R2358_U562, P1_R2358_U563, P1_R2358_U564, P1_R2358_U565, P1_R2358_U566, P1_R2358_U567, P1_R2358_U568, P1_R2358_U569, P1_R2358_U570, P1_R2358_U571, P1_R2358_U572, P1_R2358_U573, P1_R2358_U574, P1_R2358_U575, P1_R2358_U576, P1_R2358_U577, P1_R2358_U578, P1_R2358_U579, P1_R2358_U580, P1_R2358_U581, P1_R2358_U582, P1_R2358_U583, P1_R2358_U584, P1_R2358_U585, P1_R2358_U586, P1_R2358_U587, P1_R2358_U588, P1_R2358_U589, P1_R2358_U590, P1_R2358_U591, P1_R2358_U592, P1_R2358_U593, P1_R2358_U594, P1_R2358_U595, P1_R2358_U596, P1_R2358_U597, P1_R2358_U598, P1_R2358_U599, P1_R2358_U600, P1_R2358_U601, P1_R2358_U602, P1_R2358_U603, P1_R2358_U604, P1_R2358_U605, P1_R2358_U606, P1_R2358_U607, P1_R2358_U608, P1_R2358_U609, P1_R2358_U610, P1_R2358_U611, P1_LT_589_U6, P1_LT_589_U7, P1_LT_589_U8, P1_R584_U6, P1_R584_U7, P1_R584_U8, P1_R584_U9, P1_R2099_U4, P1_R2099_U5, P1_R2099_U6, P1_R2099_U7, P1_R2099_U8, P1_R2099_U9, P1_R2099_U10, P1_R2099_U11, P1_R2099_U12, P1_R2099_U13, P1_R2099_U14, P1_R2099_U15, P1_R2099_U16, P1_R2099_U17, P1_R2099_U18, P1_R2099_U19, P1_R2099_U20, P1_R2099_U21, P1_R2099_U22, P1_R2099_U23, P1_R2099_U24, P1_R2099_U25, P1_R2099_U26, P1_R2099_U27, P1_R2099_U28, P1_R2099_U29, P1_R2099_U30, P1_R2099_U31, P1_R2099_U32, P1_R2099_U33, P1_R2099_U34, P1_R2099_U35, P1_R2099_U36, P1_R2099_U37, P1_R2099_U38, P1_R2099_U39, P1_R2099_U40, P1_R2099_U41, P1_R2099_U42, P1_R2099_U43, P1_R2099_U44, P1_R2099_U45, P1_R2099_U46, P1_R2099_U47, P1_R2099_U48, P1_R2099_U49, P1_R2099_U50, P1_R2099_U51, P1_R2099_U52, P1_R2099_U53, P1_R2099_U54, P1_R2099_U55, P1_R2099_U56, P1_R2099_U57, P1_R2099_U58, P1_R2099_U59, P1_R2099_U60, P1_R2099_U61, P1_R2099_U62, P1_R2099_U63, P1_R2099_U64, P1_R2099_U65, P1_R2099_U66, P1_R2099_U67, P1_R2099_U68, P1_R2099_U69, P1_R2099_U70, P1_R2099_U71, P1_R2099_U72, P1_R2099_U73, P1_R2099_U74, P1_R2099_U75, P1_R2099_U76, P1_R2099_U77, P1_R2099_U78, P1_R2099_U79, P1_R2099_U80, P1_R2099_U81, P1_R2099_U82, P1_R2099_U83, P1_R2099_U84, P1_R2099_U85, P1_R2099_U86, P1_R2099_U87, P1_R2099_U88, P1_R2099_U89, P1_R2099_U90, P1_R2099_U91, P1_R2099_U92, P1_R2099_U93, P1_R2099_U94, P1_R2099_U95, P1_R2099_U96, P1_R2099_U97, P1_R2099_U98, P1_R2099_U99, P1_R2099_U100, P1_R2099_U101, P1_R2099_U102, P1_R2099_U103, P1_R2099_U104, P1_R2099_U105, P1_R2099_U106, P1_R2099_U107, P1_R2099_U108, P1_R2099_U109, P1_R2099_U110, P1_R2099_U111, P1_R2099_U112, P1_R2099_U113, P1_R2099_U114, P1_R2099_U115, P1_R2099_U116, P1_R2099_U117, P1_R2099_U118, P1_R2099_U119, P1_R2099_U120, P1_R2099_U121, P1_R2099_U122, P1_R2099_U123, P1_R2099_U124, P1_R2099_U125, P1_R2099_U126, P1_R2099_U127, P1_R2099_U128, P1_R2099_U129, P1_R2099_U130, P1_R2099_U131, P1_R2099_U132, P1_R2099_U133, P1_R2099_U134, P1_R2099_U135, P1_R2099_U136, P1_R2099_U137, P1_R2099_U138, P1_R2099_U139, P1_R2099_U140, P1_R2099_U141, P1_R2099_U142, P1_R2099_U143, P1_R2099_U144, P1_R2099_U145, P1_R2099_U146, P1_R2099_U147, P1_R2099_U148, P1_R2099_U149, P1_R2099_U150, P1_R2099_U151, P1_R2099_U152, P1_R2099_U153, P1_R2099_U154, P1_R2099_U155, P1_R2099_U156, P1_R2099_U157, P1_R2099_U158, P1_R2099_U159, P1_R2099_U160, P1_R2099_U161, P1_R2099_U162, P1_R2099_U163, P1_R2099_U164, P1_R2099_U165, P1_R2099_U166, P1_R2099_U167, P1_R2099_U168, P1_R2099_U169, P1_R2099_U170, P1_R2099_U171, P1_R2099_U172, P1_R2099_U173, P1_R2099_U174, P1_R2099_U175, P1_R2099_U176, P1_R2099_U177, P1_R2099_U178, P1_R2099_U179, P1_R2099_U180, P1_R2099_U181, P1_R2099_U182, P1_R2099_U183, P1_R2099_U184, P1_R2099_U185, P1_R2099_U186, P1_R2099_U187, P1_R2099_U188, P1_R2099_U189, P1_R2099_U190, P1_R2099_U191, P1_R2099_U192, P1_R2099_U193, P1_R2099_U194, P1_R2099_U195, P1_R2099_U196, P1_R2099_U197, P1_R2099_U198, P1_R2099_U199, P1_R2099_U200, P1_R2099_U201, P1_R2099_U202, P1_R2099_U203, P1_R2099_U204, P1_R2099_U205, P1_R2099_U206, P1_R2099_U207, P1_R2099_U208, P1_R2099_U209, P1_R2099_U210, P1_R2099_U211, P1_R2099_U212, P1_R2099_U213, P1_R2099_U214, P1_R2099_U215, P1_R2099_U216, P1_R2099_U217, P1_R2099_U218, P1_R2099_U219, P1_R2099_U220, P1_R2099_U221, P1_R2099_U222, P1_R2099_U223, P1_R2099_U224, P1_R2099_U225, P1_R2099_U226, P1_R2099_U227, P1_R2099_U228, P1_R2099_U229, P1_R2099_U230, P1_R2099_U231, P1_R2099_U232, P1_R2099_U233, P1_R2099_U234, P1_R2099_U235, P1_R2099_U236, P1_R2099_U237, P1_R2099_U238, P1_R2099_U239, P1_R2099_U240, P1_R2099_U241, P1_R2099_U242, P1_R2099_U243, P1_R2099_U244, P1_R2099_U245, P1_R2099_U246, P1_R2099_U247, P1_R2099_U248, P1_R2099_U249, P1_R2099_U250, P1_R2099_U251, P1_R2099_U252, P1_R2099_U253, P1_R2099_U254, P1_R2099_U255, P1_R2099_U256, P1_R2099_U257, P1_R2099_U258, P1_R2099_U259, P1_R2099_U260, P1_R2099_U261, P1_R2099_U262, P1_R2099_U263, P1_R2099_U264, P1_R2099_U265, P1_R2099_U266, P1_R2099_U267, P1_R2099_U268, P1_R2099_U269, P1_R2099_U270, P1_R2099_U271, P1_R2099_U272, P1_R2099_U273, P1_R2099_U274, P1_R2099_U275, P1_R2099_U276, P1_R2099_U277, P1_R2099_U278, P1_R2099_U279, P1_R2099_U280, P1_R2099_U281, P1_R2099_U282, P1_R2099_U283, P1_R2099_U284, P1_R2099_U285, P1_R2099_U286, P1_R2099_U287, P1_R2099_U288, P1_R2099_U289, P1_R2099_U290, P1_R2099_U291, P1_R2099_U292, P1_R2099_U293, P1_R2099_U294, P1_R2099_U295, P1_R2099_U296, P1_R2099_U297, P1_R2099_U298, P1_R2099_U299, P1_R2099_U300, P1_R2099_U301, P1_R2099_U302, P1_R2099_U303, P1_R2099_U304, P1_R2099_U305, P1_R2099_U306, P1_R2099_U307, P1_R2099_U308, P1_R2099_U309, P1_R2099_U310, P1_R2099_U311, P1_R2099_U312, P1_R2099_U313, P1_R2099_U314, P1_R2099_U315, P1_R2099_U316, P1_R2099_U317, P1_R2099_U318, P1_R2099_U319, P1_R2099_U320, P1_R2099_U321, P1_R2099_U322, P1_R2099_U323, P1_R2099_U324, P1_R2099_U325, P1_R2099_U326, P1_R2099_U327, P1_R2099_U328, P1_R2099_U329, P1_R2099_U330, P1_R2099_U331, P1_R2099_U332, P1_R2099_U333, P1_R2099_U334, P1_R2099_U335, P1_R2099_U336, P1_R2099_U337, P1_R2099_U338, P1_R2099_U339, P1_R2099_U340, P1_R2099_U341, P1_R2099_U342, P1_R2099_U343, P1_R2099_U344, P1_R2099_U345, P1_R2099_U346, P1_R2099_U347, P1_R2099_U348, P1_R2099_U349, P1_R2167_U6, P1_R2167_U7, P1_R2167_U8, P1_R2167_U9, P1_R2167_U10, P1_R2167_U11, P1_R2167_U12, P1_R2167_U13, P1_R2167_U14, P1_R2167_U15, P1_R2167_U16, P1_R2167_U17, P1_R2167_U18, P1_R2167_U19, P1_R2167_U20, P1_R2167_U21, P1_R2167_U22, P1_R2167_U23, P1_R2167_U24, P1_R2167_U25, P1_R2167_U26, P1_R2167_U27, P1_R2167_U28, P1_R2167_U29, P1_R2167_U30, P1_R2167_U31, P1_R2167_U32, P1_R2167_U33, P1_R2167_U34, P1_R2167_U35, P1_R2167_U36, P1_R2167_U37, P1_R2167_U38, P1_R2167_U39, P1_R2167_U40, P1_R2167_U41, P1_R2167_U42, P1_R2167_U43, P1_R2167_U44, P1_R2167_U45, P1_R2167_U46, P1_R2167_U47, P1_R2167_U48, P1_R2167_U49, P1_R2167_U50, P1_R2337_U4, P1_R2337_U5, P1_R2337_U6, P1_R2337_U7, P1_R2337_U8, P1_R2337_U9, P1_R2337_U10, P1_R2337_U11, P1_R2337_U12, P1_R2337_U13, P1_R2337_U14, P1_R2337_U15, P1_R2337_U16, P1_R2337_U17, P1_R2337_U18, P1_R2337_U19, P1_R2337_U20, P1_R2337_U21, P1_R2337_U22, P1_R2337_U23, P1_R2337_U24, P1_R2337_U25, P1_R2337_U26, P1_R2337_U27, P1_R2337_U28, P1_R2337_U29, P1_R2337_U30, P1_R2337_U31, P1_R2337_U32, P1_R2337_U33, P1_R2337_U34, P1_R2337_U35, P1_R2337_U36, P1_R2337_U37, P1_R2337_U38, P1_R2337_U39, P1_R2337_U40, P1_R2337_U41, P1_R2337_U42, P1_R2337_U43, P1_R2337_U44, P1_R2337_U45, P1_R2337_U46, P1_R2337_U47, P1_R2337_U48, P1_R2337_U49, P1_R2337_U50, P1_R2337_U51, P1_R2337_U52, P1_R2337_U53, P1_R2337_U54, P1_R2337_U55, P1_R2337_U56, P1_R2337_U57, P1_R2337_U58, P1_R2337_U59, P1_R2337_U60, P1_R2337_U61, P1_R2337_U62, P1_R2337_U63, P1_R2337_U64, P1_R2337_U65, P1_R2337_U66, P1_R2337_U67, P1_R2337_U68, P1_R2337_U69, P1_R2337_U70, P1_R2337_U71, P1_R2337_U72, P1_R2337_U73, P1_R2337_U74, P1_R2337_U75, P1_R2337_U76, P1_R2337_U77, P1_R2337_U78, P1_R2337_U79, P1_R2337_U80, P1_R2337_U81, P1_R2337_U82, P1_R2337_U83, P1_R2337_U84, P1_R2337_U85, P1_R2337_U86, P1_R2337_U87, P1_R2337_U88, P1_R2337_U89, P1_R2337_U90, P1_R2337_U91, P1_R2337_U92, P1_R2337_U93, P1_R2337_U94, P1_R2337_U95, P1_R2337_U96, P1_R2337_U97, P1_R2337_U98, P1_R2337_U99, P1_R2337_U100, P1_R2337_U101, P1_R2337_U102, P1_R2337_U103, P1_R2337_U104, P1_R2337_U105, P1_R2337_U106, P1_R2337_U107, P1_R2337_U108, P1_R2337_U109, P1_R2337_U110, P1_R2337_U111, P1_R2337_U112, P1_R2337_U113, P1_R2337_U114, P1_R2337_U115, P1_R2337_U116, P1_R2337_U117, P1_R2337_U118, P1_R2337_U119, P1_R2337_U120, P1_R2337_U121, P1_R2337_U122, P1_R2337_U123, P1_R2337_U124, P1_R2337_U125, P1_R2337_U126, P1_R2337_U127, P1_R2337_U128, P1_R2337_U129, P1_R2337_U130, P1_R2337_U131, P1_R2337_U132, P1_R2337_U133, P1_R2337_U134, P1_R2337_U135, P1_R2337_U136, P1_R2337_U137, P1_R2337_U138, P1_R2337_U139, P1_R2337_U140, P1_R2337_U141, P1_R2337_U142, P1_R2337_U143, P1_R2337_U144, P1_R2337_U145, P1_R2337_U146, P1_R2337_U147, P1_R2337_U148, P1_R2337_U149, P1_R2337_U150, P1_R2337_U151, P1_R2337_U152, P1_R2337_U153, P1_R2337_U154, P1_R2337_U155, P1_R2337_U156, P1_R2337_U157, P1_R2337_U158, P1_R2337_U159, P1_R2337_U160, P1_R2337_U161, P1_R2337_U162, P1_R2337_U163, P1_R2337_U164, P1_R2337_U165, P1_R2337_U166, P1_R2337_U167, P1_R2337_U168, P1_R2337_U169, P1_R2337_U170, P1_R2337_U171, P1_R2337_U172, P1_R2337_U173, P1_R2337_U174, P1_R2337_U175, P1_R2337_U176, P1_R2337_U177, P1_R2337_U178, P1_R2337_U179, P1_R2337_U180, P1_R2337_U181, P1_R2337_U182, P1_SUB_357_U6, P1_SUB_357_U7, P1_SUB_357_U8, P1_SUB_357_U9, P1_SUB_357_U10, P1_SUB_357_U11, P1_SUB_357_U12, P1_SUB_357_U13, P1_LT_563_1260_U6, P1_LT_563_1260_U7, P1_LT_563_1260_U8, P1_LT_563_1260_U9, P1_SUB_580_U6, P1_SUB_580_U7, P1_SUB_580_U8, P1_SUB_580_U9, P1_SUB_580_U10, P1_R2096_U4, P1_R2096_U5, P1_R2096_U6, P1_R2096_U7, P1_R2096_U8, P1_R2096_U9, P1_R2096_U10, P1_R2096_U11, P1_R2096_U12, P1_R2096_U13, P1_R2096_U14, P1_R2096_U15, P1_R2096_U16, P1_R2096_U17, P1_R2096_U18, P1_R2096_U19, P1_R2096_U20, P1_R2096_U21, P1_R2096_U22, P1_R2096_U23, P1_R2096_U24, P1_R2096_U25, P1_R2096_U26, P1_R2096_U27, P1_R2096_U28, P1_R2096_U29, P1_R2096_U30, P1_R2096_U31, P1_R2096_U32, P1_R2096_U33, P1_R2096_U34, P1_R2096_U35, P1_R2096_U36, P1_R2096_U37, P1_R2096_U38, P1_R2096_U39, P1_R2096_U40, P1_R2096_U41, P1_R2096_U42, P1_R2096_U43, P1_R2096_U44, P1_R2096_U45, P1_R2096_U46, P1_R2096_U47, P1_R2096_U48, P1_R2096_U49, P1_R2096_U50, P1_R2096_U51, P1_R2096_U52, P1_R2096_U53, P1_R2096_U54, P1_R2096_U55, P1_R2096_U56, P1_R2096_U57, P1_R2096_U58, P1_R2096_U59, P1_R2096_U60, P1_R2096_U61, P1_R2096_U62, P1_R2096_U63, P1_R2096_U64, P1_R2096_U65, P1_R2096_U66, P1_R2096_U67, P1_R2096_U68, P1_R2096_U69, P1_R2096_U70, P1_R2096_U71, P1_R2096_U72, P1_R2096_U73, P1_R2096_U74, P1_R2096_U75, P1_R2096_U76, P1_R2096_U77, P1_R2096_U78, P1_R2096_U79, P1_R2096_U80, P1_R2096_U81, P1_R2096_U82, P1_R2096_U83, P1_R2096_U84, P1_R2096_U85, P1_R2096_U86, P1_R2096_U87, P1_R2096_U88, P1_R2096_U89, P1_R2096_U90, P1_R2096_U91, P1_R2096_U92, P1_R2096_U93, P1_R2096_U94, P1_R2096_U95, P1_R2096_U96, P1_R2096_U97, P1_R2096_U98, P1_R2096_U99, P1_R2096_U100, P1_R2096_U101, P1_R2096_U102, P1_R2096_U103, P1_R2096_U104, P1_R2096_U105, P1_R2096_U106, P1_R2096_U107, P1_R2096_U108, P1_R2096_U109, P1_R2096_U110, P1_R2096_U111, P1_R2096_U112, P1_R2096_U113, P1_R2096_U114, P1_R2096_U115, P1_R2096_U116, P1_R2096_U117, P1_R2096_U118, P1_R2096_U119, P1_R2096_U120, P1_R2096_U121, P1_R2096_U122, P1_R2096_U123, P1_R2096_U124, P1_R2096_U125, P1_R2096_U126, P1_R2096_U127, P1_R2096_U128, P1_R2096_U129, P1_R2096_U130, P1_R2096_U131, P1_R2096_U132, P1_R2096_U133, P1_R2096_U134, P1_R2096_U135, P1_R2096_U136, P1_R2096_U137, P1_R2096_U138, P1_R2096_U139, P1_R2096_U140, P1_R2096_U141, P1_R2096_U142, P1_R2096_U143, P1_R2096_U144, P1_R2096_U145, P1_R2096_U146, P1_R2096_U147, P1_R2096_U148, P1_R2096_U149, P1_R2096_U150, P1_R2096_U151, P1_R2096_U152, P1_R2096_U153, P1_R2096_U154, P1_R2096_U155, P1_R2096_U156, P1_R2096_U157, P1_R2096_U158, P1_R2096_U159, P1_R2096_U160, P1_R2096_U161, P1_R2096_U162, P1_R2096_U163, P1_R2096_U164, P1_R2096_U165, P1_R2096_U166, P1_R2096_U167, P1_R2096_U168, P1_R2096_U169, P1_R2096_U170, P1_R2096_U171, P1_R2096_U172, P1_R2096_U173, P1_R2096_U174, P1_R2096_U175, P1_R2096_U176, P1_R2096_U177, P1_R2096_U178, P1_R2096_U179, P1_R2096_U180, P1_R2096_U181, P1_R2096_U182, P1_LT_563_U6, P1_LT_563_U7, P1_LT_563_U8, P1_LT_563_U9, P1_LT_563_U10, P1_LT_563_U11, P1_LT_563_U12, P1_LT_563_U13, P1_LT_563_U14, P1_LT_563_U15, P1_LT_563_U16, P1_LT_563_U17, P1_LT_563_U18, P1_LT_563_U19, P1_LT_563_U20, P1_LT_563_U21, P1_LT_563_U22, P1_LT_563_U23, P1_LT_563_U24, P1_LT_563_U25, P1_LT_563_U26, P1_LT_563_U27, P1_LT_563_U28, P1_R2238_U6, P1_R2238_U7, P1_R2238_U8, P1_R2238_U9, P1_R2238_U10, P1_R2238_U11, P1_R2238_U12, P1_R2238_U13, P1_R2238_U14, P1_R2238_U15, P1_R2238_U16, P1_R2238_U17, P1_R2238_U18, P1_R2238_U19, P1_R2238_U20, P1_R2238_U21, P1_R2238_U22, P1_R2238_U23, P1_R2238_U24, P1_R2238_U25, P1_R2238_U26, P1_R2238_U27, P1_R2238_U28, P1_R2238_U29, P1_R2238_U30, P1_R2238_U31, P1_R2238_U32, P1_R2238_U33, P1_R2238_U34, P1_R2238_U35, P1_R2238_U36, P1_R2238_U37, P1_R2238_U38, P1_R2238_U39, P1_R2238_U40, P1_R2238_U41, P1_R2238_U42, P1_R2238_U43, P1_R2238_U44, P1_R2238_U45, P1_R2238_U46, P1_R2238_U47, P1_R2238_U48, P1_R2238_U49, P1_R2238_U50, P1_R2238_U51, P1_R2238_U52, P1_R2238_U53, P1_R2238_U54, P1_R2238_U55, P1_R2238_U56, P1_R2238_U57, P1_R2238_U58, P1_R2238_U59, P1_R2238_U60, P1_R2238_U61, P1_R2238_U62, P1_R2238_U63, P1_R2238_U64, P1_R2238_U65, P1_R2238_U66, P1_SUB_450_U6, P1_SUB_450_U7, P1_SUB_450_U8, P1_SUB_450_U9, P1_SUB_450_U10, P1_SUB_450_U11, P1_SUB_450_U12, P1_SUB_450_U13, P1_SUB_450_U14, P1_SUB_450_U15, P1_SUB_450_U16, P1_SUB_450_U17, P1_SUB_450_U18, P1_SUB_450_U19, P1_SUB_450_U20, P1_SUB_450_U21, P1_SUB_450_U22, P1_SUB_450_U23, P1_SUB_450_U24, P1_SUB_450_U25, P1_SUB_450_U26, P1_SUB_450_U27, P1_SUB_450_U28, P1_SUB_450_U29, P1_SUB_450_U30, P1_SUB_450_U31, P1_SUB_450_U32, P1_SUB_450_U33, P1_SUB_450_U34, P1_SUB_450_U35, P1_SUB_450_U36, P1_SUB_450_U37, P1_SUB_450_U38, P1_SUB_450_U39, P1_SUB_450_U40, P1_SUB_450_U41, P1_SUB_450_U42, P1_SUB_450_U43, P1_SUB_450_U44, P1_SUB_450_U45, P1_SUB_450_U46, P1_SUB_450_U47, P1_SUB_450_U48, P1_SUB_450_U49, P1_SUB_450_U50, P1_SUB_450_U51, P1_SUB_450_U52, P1_SUB_450_U53, P1_SUB_450_U54, P1_SUB_450_U55, P1_SUB_450_U56, P1_SUB_450_U57, P1_SUB_450_U58, P1_SUB_450_U59, P1_SUB_450_U60, P1_SUB_450_U61, P1_SUB_450_U62, P1_SUB_450_U63, P1_SUB_450_U64, P1_SUB_450_U65, P1_SUB_450_U66, P1_ADD_371_U4, P1_ADD_371_U5, P1_ADD_371_U6, P1_ADD_371_U7, P1_ADD_371_U8, P1_ADD_371_U9, P1_ADD_371_U10, P1_ADD_371_U11, P1_ADD_371_U12, P1_ADD_371_U13, P1_ADD_371_U14, P1_ADD_371_U15, P1_ADD_371_U16, P1_ADD_371_U17, P1_ADD_371_U18, P1_ADD_371_U19, P1_ADD_371_U20, P1_ADD_371_U21, P1_ADD_371_U22, P1_ADD_371_U23, P1_ADD_371_U24, P1_ADD_371_U25, P1_ADD_371_U26, P1_ADD_371_U27, P1_ADD_371_U28, P1_ADD_371_U29, P1_ADD_371_U30, P1_ADD_371_U31, P1_ADD_371_U32, P1_ADD_371_U33, P1_ADD_371_U34, P1_ADD_371_U35, P1_ADD_371_U36, P1_ADD_371_U37, P1_ADD_371_U38, P1_ADD_371_U39, P1_ADD_371_U40, P1_ADD_371_U41, P1_ADD_371_U42, P1_ADD_371_U43, P1_ADD_371_U44, P1_ADD_405_U4, P1_ADD_405_U5, P1_ADD_405_U6, P1_ADD_405_U7, P1_ADD_405_U8, P1_ADD_405_U9, P1_ADD_405_U10, P1_ADD_405_U11, P1_ADD_405_U12, P1_ADD_405_U13, P1_ADD_405_U14, P1_ADD_405_U15, P1_ADD_405_U16, P1_ADD_405_U17, P1_ADD_405_U18, P1_ADD_405_U19, P1_ADD_405_U20, P1_ADD_405_U21, P1_ADD_405_U22, P1_ADD_405_U23, P1_ADD_405_U24, P1_ADD_405_U25, P1_ADD_405_U26, P1_ADD_405_U27, P1_ADD_405_U28, P1_ADD_405_U29, P1_ADD_405_U30, P1_ADD_405_U31, P1_ADD_405_U32, P1_ADD_405_U33, P1_ADD_405_U34, P1_ADD_405_U35, P1_ADD_405_U36, P1_ADD_405_U37, P1_ADD_405_U38, P1_ADD_405_U39, P1_ADD_405_U40, P1_ADD_405_U41, P1_ADD_405_U42, P1_ADD_405_U43, P1_ADD_405_U44, P1_ADD_405_U45, P1_ADD_405_U46, P1_ADD_405_U47, P1_ADD_405_U48, P1_ADD_405_U49, P1_ADD_405_U50, P1_ADD_405_U51, P1_ADD_405_U52, P1_ADD_405_U53, P1_ADD_405_U54, P1_ADD_405_U55, P1_ADD_405_U56, P1_ADD_405_U57, P1_ADD_405_U58, P1_ADD_405_U59, P1_ADD_405_U60, P1_ADD_405_U61, P1_ADD_405_U62, P1_ADD_405_U63, P1_ADD_405_U64, P1_ADD_405_U65, P1_ADD_405_U66, P1_ADD_405_U67, P1_ADD_405_U68, P1_ADD_405_U69, P1_ADD_405_U70, P1_ADD_405_U71, P1_ADD_405_U72, P1_ADD_405_U73, P1_ADD_405_U74, P1_ADD_405_U75, P1_ADD_405_U76, P1_ADD_405_U77, P1_ADD_405_U78, P1_ADD_405_U79, P1_ADD_405_U80, P1_ADD_405_U81, P1_ADD_405_U82, P1_ADD_405_U83, P1_ADD_405_U84, P1_ADD_405_U85, P1_ADD_405_U86, P1_ADD_405_U87, P1_ADD_405_U88, P1_ADD_405_U89, P1_ADD_405_U90, P1_ADD_405_U91, P1_ADD_405_U92, P1_ADD_405_U93, P1_ADD_405_U94, P1_ADD_405_U95, P1_ADD_405_U96, P1_ADD_405_U97, P1_ADD_405_U98, P1_ADD_405_U99, P1_ADD_405_U100, P1_ADD_405_U101, P1_ADD_405_U102, P1_ADD_405_U103, P1_ADD_405_U104, P1_ADD_405_U105, P1_ADD_405_U106, P1_ADD_405_U107, P1_ADD_405_U108, P1_ADD_405_U109, P1_ADD_405_U110, P1_ADD_405_U111, P1_ADD_405_U112, P1_ADD_405_U113, P1_ADD_405_U114, P1_ADD_405_U115, P1_ADD_405_U116, P1_ADD_405_U117, P1_ADD_405_U118, P1_ADD_405_U119, P1_ADD_405_U120, P1_ADD_405_U121, P1_ADD_405_U122, P1_ADD_405_U123, P1_ADD_405_U124, P1_ADD_405_U125, P1_ADD_405_U126, P1_ADD_405_U127, P1_ADD_405_U128, P1_ADD_405_U129, P1_ADD_405_U130, P1_ADD_405_U131, P1_ADD_405_U132, P1_ADD_405_U133, P1_ADD_405_U134, P1_ADD_405_U135, P1_ADD_405_U136, P1_ADD_405_U137, P1_ADD_405_U138, P1_ADD_405_U139, P1_ADD_405_U140, P1_ADD_405_U141, P1_ADD_405_U142, P1_ADD_405_U143, P1_ADD_405_U144, P1_ADD_405_U145, P1_ADD_405_U146, P1_ADD_405_U147, P1_ADD_405_U148, P1_ADD_405_U149, P1_ADD_405_U150, P1_ADD_405_U151, P1_ADD_405_U152, P1_ADD_405_U153, P1_ADD_405_U154, P1_ADD_405_U155, P1_ADD_405_U156, P1_ADD_405_U157, P1_ADD_405_U158, P1_ADD_405_U159, P1_ADD_405_U160, P1_ADD_405_U161, P1_ADD_405_U162, P1_ADD_405_U163, P1_ADD_405_U164, P1_ADD_405_U165, P1_ADD_405_U166, P1_ADD_405_U167, P1_ADD_405_U168, P1_ADD_405_U169, P1_ADD_405_U170, P1_ADD_405_U171, P1_ADD_405_U172, P1_ADD_405_U173, P1_ADD_405_U174, P1_ADD_405_U175, P1_ADD_405_U176, P1_ADD_405_U177, P1_ADD_405_U178, P1_ADD_405_U179, P1_ADD_405_U180, P1_ADD_405_U181, P1_ADD_405_U182, P1_ADD_405_U183, P1_ADD_405_U184, P1_ADD_405_U185, P1_ADD_405_U186, P1_GTE_485_U6, P1_GTE_485_U7, P1_ADD_515_U4, P1_ADD_515_U5, P1_ADD_515_U6, P1_ADD_515_U7, P1_ADD_515_U8, P1_ADD_515_U9, P1_ADD_515_U10, P1_ADD_515_U11, P1_ADD_515_U12, P1_ADD_515_U13, P1_ADD_515_U14, P1_ADD_515_U15, P1_ADD_515_U16, P1_ADD_515_U17, P1_ADD_515_U18, P1_ADD_515_U19, P1_ADD_515_U20, P1_ADD_515_U21, P1_ADD_515_U22, P1_ADD_515_U23, P1_ADD_515_U24, P1_ADD_515_U25, P1_ADD_515_U26, P1_ADD_515_U27, P1_ADD_515_U28, P1_ADD_515_U29, P1_ADD_515_U30, P1_ADD_515_U31, P1_ADD_515_U32, P1_ADD_515_U33, P1_ADD_515_U34, P1_ADD_515_U35, P1_ADD_515_U36, P1_ADD_515_U37, P1_ADD_515_U38, P1_ADD_515_U39, P1_ADD_515_U40, P1_ADD_515_U41, P1_ADD_515_U42, P1_ADD_515_U43, P1_ADD_515_U44, P1_ADD_515_U45, P1_ADD_515_U46, P1_ADD_515_U47, P1_ADD_515_U48, P1_ADD_515_U49, P1_ADD_515_U50, P1_ADD_515_U51, P1_ADD_515_U52, P1_ADD_515_U53, P1_ADD_515_U54, P1_ADD_515_U55, P1_ADD_515_U56, P1_ADD_515_U57, P1_ADD_515_U58, P1_ADD_515_U59, P1_ADD_515_U60, P1_ADD_515_U61, P1_ADD_515_U62, P1_ADD_515_U63, P1_ADD_515_U64, P1_ADD_515_U65, P1_ADD_515_U66, P1_ADD_515_U67, P1_ADD_515_U68, P1_ADD_515_U69, P1_ADD_515_U70, P1_ADD_515_U71, P1_ADD_515_U72, P1_ADD_515_U73, P1_ADD_515_U74, P1_ADD_515_U75, P1_ADD_515_U76, P1_ADD_515_U77, P1_ADD_515_U78, P1_ADD_515_U79, P1_ADD_515_U80, P1_ADD_515_U81, P1_ADD_515_U82, P1_ADD_515_U83, P1_ADD_515_U84, P1_ADD_515_U85, P1_ADD_515_U86, P1_ADD_515_U87, P1_ADD_515_U88, P1_ADD_515_U89, P1_ADD_515_U90, P1_ADD_515_U91, P1_ADD_515_U92, P1_ADD_515_U93, P1_ADD_515_U94, P1_ADD_515_U95, P1_ADD_515_U96, P1_ADD_515_U97, P1_ADD_515_U98, P1_ADD_515_U99, P1_ADD_515_U100, P1_ADD_515_U101, P1_ADD_515_U102, P1_ADD_515_U103, P1_ADD_515_U104, P1_ADD_515_U105, P1_ADD_515_U106, P1_ADD_515_U107, P1_ADD_515_U108, P1_ADD_515_U109, P1_ADD_515_U110, P1_ADD_515_U111, P1_ADD_515_U112, P1_ADD_515_U113, P1_ADD_515_U114, P1_ADD_515_U115, P1_ADD_515_U116, P1_ADD_515_U117, P1_ADD_515_U118, P1_ADD_515_U119, P1_ADD_515_U120, P1_ADD_515_U121, P1_ADD_515_U122, P1_ADD_515_U123, P1_ADD_515_U124, P1_ADD_515_U125, P1_ADD_515_U126, P1_ADD_515_U127, P1_ADD_515_U128, P1_ADD_515_U129, P1_ADD_515_U130, P1_ADD_515_U131, P1_ADD_515_U132, P1_ADD_515_U133, P1_ADD_515_U134, P1_ADD_515_U135, P1_ADD_515_U136, P1_ADD_515_U137, P1_ADD_515_U138, P1_ADD_515_U139, P1_ADD_515_U140, P1_ADD_515_U141, P1_ADD_515_U142, P1_ADD_515_U143, P1_ADD_515_U144, P1_ADD_515_U145, P1_ADD_515_U146, P1_ADD_515_U147, P1_ADD_515_U148, P1_ADD_515_U149, P1_ADD_515_U150, P1_ADD_515_U151, P1_ADD_515_U152, P1_ADD_515_U153, P1_ADD_515_U154, P1_ADD_515_U155, P1_ADD_515_U156, P1_ADD_515_U157, P1_ADD_515_U158, P1_ADD_515_U159, P1_ADD_515_U160, P1_ADD_515_U161, P1_ADD_515_U162, P1_ADD_515_U163, P1_ADD_515_U164, P1_ADD_515_U165, P1_ADD_515_U166, P1_ADD_515_U167, P1_ADD_515_U168, P1_ADD_515_U169, P1_ADD_515_U170, P1_ADD_515_U171, P1_ADD_515_U172, P1_ADD_515_U173, P1_ADD_515_U174, P1_ADD_515_U175, P1_ADD_515_U176, P1_ADD_515_U177, P1_ADD_515_U178, P1_ADD_515_U179, P1_ADD_515_U180, P1_ADD_515_U181, P1_ADD_515_U182; 
assign U209 = READY2 & READY22_REG_SCAN_IN; 
assign U210 = READY1 & READY11_REG_SCAN_IN; 
assign U211 = READY12_REG_SCAN_IN & READY21_REG_SCAN_IN; 
assign U377 = ~(P2_BE_N_REG_2__SCAN_IN | P2_BE_N_REG_1__SCAN_IN | P2_BE_N_REG_0__SCAN_IN | P2_ADS_N_REG_SCAN_IN); 
assign U378 = ~(P2_BE_N_REG_3__SCAN_IN | P2_D_C_N_REG_SCAN_IN); 
assign U379 = ~(P3_BE_N_REG_1__SCAN_IN | P3_BE_N_REG_0__SCAN_IN | P3_W_R_N_REG_SCAN_IN | P3_D_C_N_REG_SCAN_IN | P3_ADS_N_REG_SCAN_IN); 
assign U380 = ~(P3_BE_N_REG_3__SCAN_IN | P3_BE_N_REG_2__SCAN_IN); 
assign U381 = ~(P1_BE_N_REG_3__SCAN_IN | P1_BE_N_REG_1__SCAN_IN | P1_BE_N_REG_0__SCAN_IN | P1_D_C_N_REG_SCAN_IN | P1_ADS_N_REG_SCAN_IN); 
assign U383 = ~P1_BE_N_REG_2__SCAN_IN; 
assign P3_U2453 = P3_STATE2_REG_2__SCAN_IN & P3_STATE2_REG_1__SCAN_IN; 
assign P3_U2464 = P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P3_U2481 = ~(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_U2501 = ~(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P3_U2631 = ~P3_STATEBS16_REG_SCAN_IN; 
assign P3_U3075 = ~P3_REQUESTPENDING_REG_SCAN_IN; 
assign P3_U3076 = ~P3_STATE_REG_1__SCAN_IN; 
assign P3_U3079 = ~P3_STATE_REG_2__SCAN_IN; 
assign P3_U3081 = ~P3_REIP_REG_1__SCAN_IN; 
assign P3_U3083 = P3_STATE_REG_2__SCAN_IN | P3_STATE_REG_1__SCAN_IN; 
assign P3_U3084 = ~HOLD; 
assign P3_U3085 = ~P3_STATE_REG_0__SCAN_IN; 
assign P3_U3088 = HOLD | P3_REQUESTPENDING_REG_SCAN_IN; 
assign P3_U3089 = ~P3_STATE2_REG_1__SCAN_IN; 
assign P3_U3090 = ~P3_STATE2_REG_2__SCAN_IN; 
assign P3_U3091 = P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P3_U3093 = ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P3_U3094 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P3_U3095 = ~(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P3_U3097 = ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P3_U3100 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P3_U3121 = ~P3_STATE2_REG_0__SCAN_IN; 
assign P3_U3123 = P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_1__SCAN_IN; 
assign P3_U3125 = P3_STATE2_REG_2__SCAN_IN | P3_STATE2_REG_1__SCAN_IN; 
assign P3_U3128 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN; 
assign P3_U3129 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign P3_U3130 = ~(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P3_U3131 = ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P3_U3133 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign P3_U3135 = P3_STATE2_REG_3__SCAN_IN | P3_STATE2_REG_2__SCAN_IN; 
assign P3_U3207 = ~P3_FLUSH_REG_SCAN_IN; 
assign P3_U3240 = ~P3_REIP_REG_0__SCAN_IN; 
assign P3_U3256 = ~P3_EBX_REG_31__SCAN_IN; 
assign P3_U3263 = ~P3_CODEFETCH_REG_SCAN_IN; 
assign P3_U3264 = ~P3_READREQUEST_REG_SCAN_IN; 
assign P3_U3291 = ~(P3_DATAWIDTH_REG_1__SCAN_IN | P3_REIP_REG_1__SCAN_IN); 
assign P3_U3312 = P3_STATE_REG_0__SCAN_IN & P3_REQUESTPENDING_REG_SCAN_IN; 
assign P3_U3365 = P3_STATE2_REG_3__SCAN_IN & P3_STATE2_REG_0__SCAN_IN; 
assign P3_U3386 = P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign P3_U3404 = P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P3_U3457 = P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign P3_U3563 = ~(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_U3581 = ~(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_U3616 = ~(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_U3634 = ~(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_U3653 = P3_STATE2_REG_0__SCAN_IN & P3_FLUSH_REG_SCAN_IN; 
assign P3_U4136 = ~(P3_DATAWIDTH_REG_2__SCAN_IN | P3_DATAWIDTH_REG_3__SCAN_IN | P3_DATAWIDTH_REG_4__SCAN_IN | P3_DATAWIDTH_REG_5__SCAN_IN); 
assign P3_U4137 = ~(P3_DATAWIDTH_REG_6__SCAN_IN | P3_DATAWIDTH_REG_7__SCAN_IN | P3_DATAWIDTH_REG_8__SCAN_IN | P3_DATAWIDTH_REG_9__SCAN_IN); 
assign P3_U4139 = ~(P3_DATAWIDTH_REG_10__SCAN_IN | P3_DATAWIDTH_REG_11__SCAN_IN | P3_DATAWIDTH_REG_12__SCAN_IN | P3_DATAWIDTH_REG_13__SCAN_IN); 
assign P3_U4140 = ~(P3_DATAWIDTH_REG_14__SCAN_IN | P3_DATAWIDTH_REG_15__SCAN_IN | P3_DATAWIDTH_REG_16__SCAN_IN | P3_DATAWIDTH_REG_17__SCAN_IN); 
assign P3_U4142 = ~(P3_DATAWIDTH_REG_18__SCAN_IN | P3_DATAWIDTH_REG_19__SCAN_IN | P3_DATAWIDTH_REG_20__SCAN_IN | P3_DATAWIDTH_REG_21__SCAN_IN); 
assign P3_U4143 = ~(P3_DATAWIDTH_REG_22__SCAN_IN | P3_DATAWIDTH_REG_23__SCAN_IN | P3_DATAWIDTH_REG_24__SCAN_IN | P3_DATAWIDTH_REG_25__SCAN_IN); 
assign P3_U4145 = ~(P3_DATAWIDTH_REG_26__SCAN_IN | P3_DATAWIDTH_REG_27__SCAN_IN); 
assign P3_U4146 = ~(P3_DATAWIDTH_REG_28__SCAN_IN | P3_DATAWIDTH_REG_29__SCAN_IN); 
assign P3_U4147 = ~(P3_DATAWIDTH_REG_30__SCAN_IN | P3_DATAWIDTH_REG_31__SCAN_IN); 
assign P3_U4149 = ~(P3_DATAWIDTH_REG_0__SCAN_IN | P3_DATAWIDTH_REG_1__SCAN_IN | P3_REIP_REG_0__SCAN_IN); 
assign P3_U4284 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_U4286 = ~BS16; 
assign P3_U4450 = NA | P3_STATE_REG_0__SCAN_IN; 
assign P3_U4624 = P3_FLUSH_REG_SCAN_IN | P3_MORE_REG_SCAN_IN; 
assign P3_U5503 = ~(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P3_U7366 = ~(P3_DATAWIDTH_REG_0__SCAN_IN & P3_DATAWIDTH_REG_1__SCAN_IN); 
assign P3_U7367 = P3_REIP_REG_0__SCAN_IN | P3_REIP_REG_1__SCAN_IN; 
assign P3_U7383 = ~(P3_STATE_REG_0__SCAN_IN & P3_ADS_N_REG_SCAN_IN); 
assign P3_U7935 = P3_STATE_REG_1__SCAN_IN | P3_STATE_REG_0__SCAN_IN; 
assign P3_U7956 = P3_STATE2_REG_0__SCAN_IN | P3_STATEBS16_REG_SCAN_IN; 
assign P3_U7987 = ~(P3_INSTADDRPOINTER_REG_0__SCAN_IN & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_U8004 = P3_DATAWIDTH_REG_0__SCAN_IN | P3_DATAWIDTH_REG_1__SCAN_IN; 
assign P3_U8008 = ~(P3_REIP_REG_0__SCAN_IN & P3_REIP_REG_1__SCAN_IN); 
assign P2_U2448 = P2_STATE2_REG_2__SCAN_IN & P2_STATE2_REG_1__SCAN_IN; 
assign P2_U2464 = P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P2_U2478 = ~(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P2_U2503 = ~(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P2_U3244 = ~P2_STATE_REG_2__SCAN_IN; 
assign P2_U3256 = ~P2_REQUESTPENDING_REG_SCAN_IN; 
assign P2_U3258 = ~P2_STATE_REG_1__SCAN_IN; 
assign P2_U3263 = P2_STATE_REG_2__SCAN_IN | P2_STATE_REG_1__SCAN_IN; 
assign P2_U3264 = ~HOLD; 
assign P2_U3266 = ~P2_STATE_REG_0__SCAN_IN; 
assign P2_U3268 = HOLD | P2_REQUESTPENDING_REG_SCAN_IN; 
assign P2_U3269 = ~P2_STATE2_REG_1__SCAN_IN; 
assign P2_U3270 = ~P2_STATE2_REG_2__SCAN_IN; 
assign P2_U3271 = ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P2_U3272 = ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P2_U3273 = ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U3275 = P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P2_U3276 = ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P2_U3277 = ~(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P2_U3284 = ~P2_STATE2_REG_0__SCAN_IN; 
assign P2_U3300 = ~P2_STATE2_REG_3__SCAN_IN; 
assign P2_U3302 = ~P2_STATEBS16_REG_SCAN_IN; 
assign P2_U3303 = P2_STATE2_REG_3__SCAN_IN | P2_STATE2_REG_1__SCAN_IN; 
assign P2_U3307 = ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN; 
assign P2_U3308 = ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign P2_U3309 = ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign P2_U3310 = ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P2_U3311 = ~(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P2_U3313 = P2_STATE2_REG_3__SCAN_IN | P2_STATE2_REG_2__SCAN_IN; 
assign P2_U3327 = ~P2_INSTQUEUE_REG_15__7__SCAN_IN; 
assign P2_U3328 = ~P2_INSTQUEUE_REG_15__6__SCAN_IN; 
assign P2_U3329 = ~P2_INSTQUEUE_REG_15__5__SCAN_IN; 
assign P2_U3330 = ~P2_INSTQUEUE_REG_15__4__SCAN_IN; 
assign P2_U3331 = ~P2_INSTQUEUE_REG_15__3__SCAN_IN; 
assign P2_U3332 = ~P2_INSTQUEUE_REG_15__2__SCAN_IN; 
assign P2_U3333 = ~P2_INSTQUEUE_REG_15__1__SCAN_IN; 
assign P2_U3334 = ~P2_INSTQUEUE_REG_15__0__SCAN_IN; 
assign P2_U3341 = ~P2_INSTQUEUE_REG_14__7__SCAN_IN; 
assign P2_U3342 = ~P2_INSTQUEUE_REG_14__6__SCAN_IN; 
assign P2_U3343 = ~P2_INSTQUEUE_REG_14__5__SCAN_IN; 
assign P2_U3344 = ~P2_INSTQUEUE_REG_14__4__SCAN_IN; 
assign P2_U3345 = ~P2_INSTQUEUE_REG_14__3__SCAN_IN; 
assign P2_U3346 = ~P2_INSTQUEUE_REG_14__2__SCAN_IN; 
assign P2_U3347 = ~P2_INSTQUEUE_REG_14__1__SCAN_IN; 
assign P2_U3348 = ~P2_INSTQUEUE_REG_14__0__SCAN_IN; 
assign P2_U3357 = ~P2_INSTQUEUE_REG_13__7__SCAN_IN; 
assign P2_U3358 = ~P2_INSTQUEUE_REG_13__6__SCAN_IN; 
assign P2_U3359 = ~P2_INSTQUEUE_REG_13__5__SCAN_IN; 
assign P2_U3360 = ~P2_INSTQUEUE_REG_13__4__SCAN_IN; 
assign P2_U3361 = ~P2_INSTQUEUE_REG_13__3__SCAN_IN; 
assign P2_U3362 = ~P2_INSTQUEUE_REG_13__2__SCAN_IN; 
assign P2_U3363 = ~P2_INSTQUEUE_REG_13__1__SCAN_IN; 
assign P2_U3364 = ~P2_INSTQUEUE_REG_13__0__SCAN_IN; 
assign P2_U3368 = ~P2_INSTQUEUE_REG_12__7__SCAN_IN; 
assign P2_U3369 = ~P2_INSTQUEUE_REG_12__6__SCAN_IN; 
assign P2_U3370 = ~P2_INSTQUEUE_REG_12__5__SCAN_IN; 
assign P2_U3371 = ~P2_INSTQUEUE_REG_12__4__SCAN_IN; 
assign P2_U3372 = ~P2_INSTQUEUE_REG_12__3__SCAN_IN; 
assign P2_U3373 = ~P2_INSTQUEUE_REG_12__2__SCAN_IN; 
assign P2_U3374 = ~P2_INSTQUEUE_REG_12__1__SCAN_IN; 
assign P2_U3375 = ~P2_INSTQUEUE_REG_12__0__SCAN_IN; 
assign P2_U3382 = ~P2_INSTQUEUE_REG_11__7__SCAN_IN; 
assign P2_U3383 = ~P2_INSTQUEUE_REG_11__6__SCAN_IN; 
assign P2_U3384 = ~P2_INSTQUEUE_REG_11__5__SCAN_IN; 
assign P2_U3385 = ~P2_INSTQUEUE_REG_11__4__SCAN_IN; 
assign P2_U3386 = ~P2_INSTQUEUE_REG_11__3__SCAN_IN; 
assign P2_U3387 = ~P2_INSTQUEUE_REG_11__2__SCAN_IN; 
assign P2_U3388 = ~P2_INSTQUEUE_REG_11__1__SCAN_IN; 
assign P2_U3389 = ~P2_INSTQUEUE_REG_11__0__SCAN_IN; 
assign P2_U3393 = ~P2_INSTQUEUE_REG_10__7__SCAN_IN; 
assign P2_U3394 = ~P2_INSTQUEUE_REG_10__6__SCAN_IN; 
assign P2_U3395 = ~P2_INSTQUEUE_REG_10__5__SCAN_IN; 
assign P2_U3396 = ~P2_INSTQUEUE_REG_10__4__SCAN_IN; 
assign P2_U3397 = ~P2_INSTQUEUE_REG_10__3__SCAN_IN; 
assign P2_U3398 = ~P2_INSTQUEUE_REG_10__2__SCAN_IN; 
assign P2_U3399 = ~P2_INSTQUEUE_REG_10__1__SCAN_IN; 
assign P2_U3400 = ~P2_INSTQUEUE_REG_10__0__SCAN_IN; 
assign P2_U3405 = ~P2_INSTQUEUE_REG_9__7__SCAN_IN; 
assign P2_U3406 = ~P2_INSTQUEUE_REG_9__6__SCAN_IN; 
assign P2_U3407 = ~P2_INSTQUEUE_REG_9__5__SCAN_IN; 
assign P2_U3408 = ~P2_INSTQUEUE_REG_9__4__SCAN_IN; 
assign P2_U3409 = ~P2_INSTQUEUE_REG_9__3__SCAN_IN; 
assign P2_U3410 = ~P2_INSTQUEUE_REG_9__2__SCAN_IN; 
assign P2_U3411 = ~P2_INSTQUEUE_REG_9__1__SCAN_IN; 
assign P2_U3412 = ~P2_INSTQUEUE_REG_9__0__SCAN_IN; 
assign P2_U3416 = ~P2_INSTQUEUE_REG_8__7__SCAN_IN; 
assign P2_U3417 = ~P2_INSTQUEUE_REG_8__6__SCAN_IN; 
assign P2_U3418 = ~P2_INSTQUEUE_REG_8__5__SCAN_IN; 
assign P2_U3419 = ~P2_INSTQUEUE_REG_8__4__SCAN_IN; 
assign P2_U3420 = ~P2_INSTQUEUE_REG_8__3__SCAN_IN; 
assign P2_U3421 = ~P2_INSTQUEUE_REG_8__2__SCAN_IN; 
assign P2_U3422 = ~P2_INSTQUEUE_REG_8__1__SCAN_IN; 
assign P2_U3423 = ~P2_INSTQUEUE_REG_8__0__SCAN_IN; 
assign P2_U3431 = ~P2_INSTQUEUE_REG_7__7__SCAN_IN; 
assign P2_U3432 = ~P2_INSTQUEUE_REG_7__6__SCAN_IN; 
assign P2_U3433 = ~P2_INSTQUEUE_REG_7__5__SCAN_IN; 
assign P2_U3434 = ~P2_INSTQUEUE_REG_7__4__SCAN_IN; 
assign P2_U3435 = ~P2_INSTQUEUE_REG_7__3__SCAN_IN; 
assign P2_U3436 = ~P2_INSTQUEUE_REG_7__2__SCAN_IN; 
assign P2_U3437 = ~P2_INSTQUEUE_REG_7__1__SCAN_IN; 
assign P2_U3438 = ~P2_INSTQUEUE_REG_7__0__SCAN_IN; 
assign P2_U3442 = ~P2_INSTQUEUE_REG_6__7__SCAN_IN; 
assign P2_U3443 = ~P2_INSTQUEUE_REG_6__6__SCAN_IN; 
assign P2_U3444 = ~P2_INSTQUEUE_REG_6__5__SCAN_IN; 
assign P2_U3445 = ~P2_INSTQUEUE_REG_6__4__SCAN_IN; 
assign P2_U3446 = ~P2_INSTQUEUE_REG_6__3__SCAN_IN; 
assign P2_U3447 = ~P2_INSTQUEUE_REG_6__2__SCAN_IN; 
assign P2_U3448 = ~P2_INSTQUEUE_REG_6__1__SCAN_IN; 
assign P2_U3449 = ~P2_INSTQUEUE_REG_6__0__SCAN_IN; 
assign P2_U3454 = ~P2_INSTQUEUE_REG_5__7__SCAN_IN; 
assign P2_U3455 = ~P2_INSTQUEUE_REG_5__6__SCAN_IN; 
assign P2_U3456 = ~P2_INSTQUEUE_REG_5__5__SCAN_IN; 
assign P2_U3457 = ~P2_INSTQUEUE_REG_5__4__SCAN_IN; 
assign P2_U3458 = ~P2_INSTQUEUE_REG_5__3__SCAN_IN; 
assign P2_U3459 = ~P2_INSTQUEUE_REG_5__2__SCAN_IN; 
assign P2_U3460 = ~P2_INSTQUEUE_REG_5__1__SCAN_IN; 
assign P2_U3461 = ~P2_INSTQUEUE_REG_5__0__SCAN_IN; 
assign P2_U3465 = ~P2_INSTQUEUE_REG_4__7__SCAN_IN; 
assign P2_U3466 = ~P2_INSTQUEUE_REG_4__6__SCAN_IN; 
assign P2_U3467 = ~P2_INSTQUEUE_REG_4__5__SCAN_IN; 
assign P2_U3468 = ~P2_INSTQUEUE_REG_4__4__SCAN_IN; 
assign P2_U3469 = ~P2_INSTQUEUE_REG_4__3__SCAN_IN; 
assign P2_U3470 = ~P2_INSTQUEUE_REG_4__2__SCAN_IN; 
assign P2_U3471 = ~P2_INSTQUEUE_REG_4__1__SCAN_IN; 
assign P2_U3472 = ~P2_INSTQUEUE_REG_4__0__SCAN_IN; 
assign P2_U3477 = ~P2_INSTQUEUE_REG_3__7__SCAN_IN; 
assign P2_U3478 = ~P2_INSTQUEUE_REG_3__6__SCAN_IN; 
assign P2_U3479 = ~P2_INSTQUEUE_REG_3__5__SCAN_IN; 
assign P2_U3480 = ~P2_INSTQUEUE_REG_3__4__SCAN_IN; 
assign P2_U3481 = ~P2_INSTQUEUE_REG_3__3__SCAN_IN; 
assign P2_U3482 = ~P2_INSTQUEUE_REG_3__2__SCAN_IN; 
assign P2_U3483 = ~P2_INSTQUEUE_REG_3__1__SCAN_IN; 
assign P2_U3484 = ~P2_INSTQUEUE_REG_3__0__SCAN_IN; 
assign P2_U3488 = ~P2_INSTQUEUE_REG_2__7__SCAN_IN; 
assign P2_U3489 = ~P2_INSTQUEUE_REG_2__6__SCAN_IN; 
assign P2_U3490 = ~P2_INSTQUEUE_REG_2__5__SCAN_IN; 
assign P2_U3491 = ~P2_INSTQUEUE_REG_2__4__SCAN_IN; 
assign P2_U3492 = ~P2_INSTQUEUE_REG_2__3__SCAN_IN; 
assign P2_U3493 = ~P2_INSTQUEUE_REG_2__2__SCAN_IN; 
assign P2_U3494 = ~P2_INSTQUEUE_REG_2__1__SCAN_IN; 
assign P2_U3495 = ~P2_INSTQUEUE_REG_2__0__SCAN_IN; 
assign P2_U3500 = ~P2_INSTQUEUE_REG_1__7__SCAN_IN; 
assign P2_U3501 = ~P2_INSTQUEUE_REG_1__6__SCAN_IN; 
assign P2_U3502 = ~P2_INSTQUEUE_REG_1__5__SCAN_IN; 
assign P2_U3503 = ~P2_INSTQUEUE_REG_1__4__SCAN_IN; 
assign P2_U3504 = ~P2_INSTQUEUE_REG_1__3__SCAN_IN; 
assign P2_U3505 = ~P2_INSTQUEUE_REG_1__2__SCAN_IN; 
assign P2_U3506 = ~P2_INSTQUEUE_REG_1__1__SCAN_IN; 
assign P2_U3507 = ~P2_INSTQUEUE_REG_1__0__SCAN_IN; 
assign P2_U3511 = ~P2_INSTQUEUE_REG_0__7__SCAN_IN; 
assign P2_U3512 = ~P2_INSTQUEUE_REG_0__6__SCAN_IN; 
assign P2_U3513 = ~P2_INSTQUEUE_REG_0__5__SCAN_IN; 
assign P2_U3514 = ~P2_INSTQUEUE_REG_0__4__SCAN_IN; 
assign P2_U3515 = ~P2_INSTQUEUE_REG_0__3__SCAN_IN; 
assign P2_U3516 = ~P2_INSTQUEUE_REG_0__2__SCAN_IN; 
assign P2_U3517 = ~P2_INSTQUEUE_REG_0__1__SCAN_IN; 
assign P2_U3518 = ~P2_INSTQUEUE_REG_0__0__SCAN_IN; 
assign P2_U3519 = ~P2_FLUSH_REG_SCAN_IN; 
assign P2_U3532 = ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P2_U3544 = ~P2_EBX_REG_31__SCAN_IN; 
assign P2_U3551 = ~P2_CODEFETCH_REG_SCAN_IN; 
assign P2_U3552 = ~P2_READREQUEST_REG_SCAN_IN; 
assign P2_U3573 = P2_STATE2_REG_1__SCAN_IN | P2_STATE2_REG_0__SCAN_IN; 
assign P2_U3606 = ~(P2_DATAWIDTH_REG_1__SCAN_IN | P2_REIP_REG_1__SCAN_IN); 
assign P2_U3692 = P2_STATE_REG_0__SCAN_IN & P2_REQUESTPENDING_REG_SCAN_IN; 
assign P2_U3719 = ~(P2_STATE2_REG_2__SCAN_IN | P2_STATE2_REG_1__SCAN_IN); 
assign P2_U3867 = P2_STATE2_REG_0__SCAN_IN & P2_FLUSH_REG_SCAN_IN; 
assign P2_U3989 = P2_STATE2_REG_1__SCAN_IN & P2_STATEBS16_REG_SCAN_IN; 
assign P2_U3990 = ~(P2_STATE2_REG_2__SCAN_IN | P2_STATE2_REG_1__SCAN_IN); 
assign P2_U4169 = ~(P2_DATAWIDTH_REG_2__SCAN_IN | P2_DATAWIDTH_REG_3__SCAN_IN | P2_DATAWIDTH_REG_4__SCAN_IN | P2_DATAWIDTH_REG_5__SCAN_IN); 
assign P2_U4170 = ~(P2_DATAWIDTH_REG_6__SCAN_IN | P2_DATAWIDTH_REG_7__SCAN_IN | P2_DATAWIDTH_REG_8__SCAN_IN | P2_DATAWIDTH_REG_9__SCAN_IN); 
assign P2_U4172 = ~(P2_DATAWIDTH_REG_10__SCAN_IN | P2_DATAWIDTH_REG_11__SCAN_IN | P2_DATAWIDTH_REG_12__SCAN_IN | P2_DATAWIDTH_REG_13__SCAN_IN); 
assign P2_U4173 = ~(P2_DATAWIDTH_REG_14__SCAN_IN | P2_DATAWIDTH_REG_15__SCAN_IN | P2_DATAWIDTH_REG_16__SCAN_IN | P2_DATAWIDTH_REG_17__SCAN_IN); 
assign P2_U4175 = ~(P2_DATAWIDTH_REG_18__SCAN_IN | P2_DATAWIDTH_REG_19__SCAN_IN | P2_DATAWIDTH_REG_20__SCAN_IN | P2_DATAWIDTH_REG_21__SCAN_IN); 
assign P2_U4176 = ~(P2_DATAWIDTH_REG_22__SCAN_IN | P2_DATAWIDTH_REG_23__SCAN_IN | P2_DATAWIDTH_REG_24__SCAN_IN | P2_DATAWIDTH_REG_25__SCAN_IN); 
assign P2_U4178 = ~(P2_DATAWIDTH_REG_26__SCAN_IN | P2_DATAWIDTH_REG_27__SCAN_IN); 
assign P2_U4179 = ~(P2_DATAWIDTH_REG_28__SCAN_IN | P2_DATAWIDTH_REG_29__SCAN_IN); 
assign P2_U4180 = ~(P2_DATAWIDTH_REG_30__SCAN_IN | P2_DATAWIDTH_REG_31__SCAN_IN); 
assign P2_U4182 = ~(P2_DATAWIDTH_REG_0__SCAN_IN | P2_DATAWIDTH_REG_1__SCAN_IN | P2_REIP_REG_0__SCAN_IN); 
assign P2_U4183 = ~(P2_DATAWIDTH_REG_1__SCAN_IN | P2_REIP_REG_1__SCAN_IN); 
assign P2_U4401 = ~BS16; 
assign P2_U4591 = ~(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P2_U4615 = P2_FLUSH_REG_SCAN_IN | P2_MORE_REG_SCAN_IN; 
assign P2_U6835 = ~(P2_DATAWIDTH_REG_0__SCAN_IN & P2_DATAWIDTH_REG_1__SCAN_IN); 
assign P2_U6851 = P2_STATE2_REG_2__SCAN_IN | P2_STATE2_REG_1__SCAN_IN; 
assign P2_U6856 = ~(P2_STATE_REG_0__SCAN_IN & P2_ADS_N_REG_SCAN_IN); 
assign P2_U7006 = P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P2_U7423 = ~(P2_STATE2_REG_3__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P2_U7425 = ~(P2_STATE2_REG_3__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P2_U7428 = ~(P2_STATE2_REG_3__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P2_U7430 = ~(P2_STATE2_REG_3__SCAN_IN & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P2_U7594 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_9__SCAN_IN); 
assign P2_U7598 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_8__SCAN_IN); 
assign P2_U7602 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_7__SCAN_IN); 
assign P2_U7606 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_6__SCAN_IN); 
assign P2_U7610 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_5__SCAN_IN); 
assign P2_U7614 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_4__SCAN_IN); 
assign P2_U7618 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_31__SCAN_IN); 
assign P2_U7622 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_30__SCAN_IN); 
assign P2_U7626 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_3__SCAN_IN); 
assign P2_U7630 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_29__SCAN_IN); 
assign P2_U7634 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_28__SCAN_IN); 
assign P2_U7638 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_27__SCAN_IN); 
assign P2_U7642 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_26__SCAN_IN); 
assign P2_U7646 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_25__SCAN_IN); 
assign P2_U7650 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_24__SCAN_IN); 
assign P2_U7654 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_23__SCAN_IN); 
assign P2_U7658 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_22__SCAN_IN); 
assign P2_U7662 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_21__SCAN_IN); 
assign P2_U7666 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_20__SCAN_IN); 
assign P2_U7670 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_2__SCAN_IN); 
assign P2_U7674 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_19__SCAN_IN); 
assign P2_U7678 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_18__SCAN_IN); 
assign P2_U7682 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_17__SCAN_IN); 
assign P2_U7686 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_16__SCAN_IN); 
assign P2_U7690 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_15__SCAN_IN); 
assign P2_U7694 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_14__SCAN_IN); 
assign P2_U7698 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_13__SCAN_IN); 
assign P2_U7702 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_12__SCAN_IN); 
assign P2_U7706 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_11__SCAN_IN); 
assign P2_U7710 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_10__SCAN_IN); 
assign P2_U7714 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_1__SCAN_IN); 
assign P2_U7719 = ~(P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_0__SCAN_IN); 
assign P2_U7898 = ~(P2_DATAWIDTH_REG_0__SCAN_IN & P2_REIP_REG_0__SCAN_IN); 
assign P2_U7908 = NA | P2_STATE_REG_0__SCAN_IN; 
assign P2_U7915 = P2_STATE_REG_1__SCAN_IN | P2_STATE_REG_0__SCAN_IN; 
assign P2_U7923 = P2_INSTQUEUE_REG_3__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7924 = P2_INSTQUEUE_REG_0__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7926 = P2_INSTQUEUE_REG_1__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7929 = P2_INSTQUEUE_REG_4__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7931 = P2_INSTQUEUE_REG_7__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7933 = P2_INSTQUEUE_REG_5__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7935 = P2_INSTQUEUE_REG_6__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7937 = P2_INSTQUEUE_REG_2__1__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7939 = P2_INSTQUEUE_REG_3__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7940 = P2_INSTQUEUE_REG_0__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7942 = P2_INSTQUEUE_REG_1__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7945 = P2_INSTQUEUE_REG_4__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7947 = P2_INSTQUEUE_REG_7__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7949 = P2_INSTQUEUE_REG_5__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7951 = P2_INSTQUEUE_REG_6__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7953 = P2_INSTQUEUE_REG_2__0__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7955 = P2_INSTQUEUE_REG_3__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7956 = P2_INSTQUEUE_REG_0__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7958 = P2_INSTQUEUE_REG_1__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7961 = P2_INSTQUEUE_REG_4__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7963 = P2_INSTQUEUE_REG_7__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7965 = P2_INSTQUEUE_REG_5__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7967 = P2_INSTQUEUE_REG_6__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7969 = P2_INSTQUEUE_REG_2__4__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7971 = P2_INSTQUEUE_REG_3__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7972 = P2_INSTQUEUE_REG_0__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7974 = P2_INSTQUEUE_REG_1__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7977 = P2_INSTQUEUE_REG_4__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7979 = P2_INSTQUEUE_REG_7__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7981 = P2_INSTQUEUE_REG_5__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7983 = P2_INSTQUEUE_REG_6__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7985 = P2_INSTQUEUE_REG_2__6__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7987 = P2_INSTQUEUE_REG_3__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7988 = P2_INSTQUEUE_REG_0__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7990 = P2_INSTQUEUE_REG_1__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7993 = P2_INSTQUEUE_REG_4__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7995 = P2_INSTQUEUE_REG_7__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7997 = P2_INSTQUEUE_REG_5__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U7999 = P2_INSTQUEUE_REG_6__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8001 = P2_INSTQUEUE_REG_2__5__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8003 = P2_INSTQUEUE_REG_3__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8004 = P2_INSTQUEUE_REG_0__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8006 = P2_INSTQUEUE_REG_1__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8009 = P2_INSTQUEUE_REG_4__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8011 = P2_INSTQUEUE_REG_7__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8013 = P2_INSTQUEUE_REG_5__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8015 = P2_INSTQUEUE_REG_6__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8017 = P2_INSTQUEUE_REG_2__2__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8019 = P2_INSTQUEUE_REG_3__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8020 = P2_INSTQUEUE_REG_0__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8022 = P2_INSTQUEUE_REG_1__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8025 = P2_INSTQUEUE_REG_4__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8027 = P2_INSTQUEUE_REG_7__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8029 = P2_INSTQUEUE_REG_5__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8031 = P2_INSTQUEUE_REG_6__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8033 = P2_INSTQUEUE_REG_2__3__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8035 = P2_INSTQUEUE_REG_3__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8036 = P2_INSTQUEUE_REG_0__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8038 = P2_INSTQUEUE_REG_1__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8041 = P2_INSTQUEUE_REG_4__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8043 = P2_INSTQUEUE_REG_7__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8045 = P2_INSTQUEUE_REG_5__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8047 = P2_INSTQUEUE_REG_6__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8049 = P2_INSTQUEUE_REG_2__7__SCAN_IN | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U8350 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P2_U8362 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P2_U8364 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P2_U8366 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P2_U8368 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P2_U8370 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P2_U8372 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P2_U8374 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P2_U8376 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P2_U8378 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P2_U8380 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P2_U8382 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P2_U8384 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P2_U8386 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P2_U8388 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P2_U8390 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P2_U8392 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P2_U8394 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P2_U8396 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P2_U8398 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P2_U8400 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P2_U8402 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P2_U8404 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P2_U8406 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P2_U8408 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P2_U8410 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P2_U8412 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P2_U8414 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P2_U8416 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P2_U8418 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P2_U8420 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P2_U8422 = ~(P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P1_U2352 = ~(P1_STATE2_REG_2__SCAN_IN | P1_STATEBS16_REG_SCAN_IN); 
assign P1_U2427 = ~(P1_STATE2_REG_3__SCAN_IN | P1_STATE2_REG_1__SCAN_IN); 
assign P1_U2428 = P1_STATE2_REG_2__SCAN_IN & P1_STATE2_REG_1__SCAN_IN; 
assign P1_U2453 = P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_U2469 = ~(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_U2478 = P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P1_U2488 = ~(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P1_U2510 = ~(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P1_U3247 = ~P1_REQUESTPENDING_REG_SCAN_IN; 
assign P1_U3248 = ~P1_STATE_REG_1__SCAN_IN; 
assign P1_U3251 = ~P1_STATE_REG_2__SCAN_IN; 
assign P1_U3253 = ~P1_REIP_REG_1__SCAN_IN; 
assign P1_U3255 = P1_STATE_REG_2__SCAN_IN | P1_STATE_REG_1__SCAN_IN; 
assign P1_U3256 = ~HOLD; 
assign P1_U3258 = ~P1_STATE_REG_0__SCAN_IN; 
assign P1_U3261 = HOLD | P1_REQUESTPENDING_REG_SCAN_IN; 
assign P1_U3262 = ~P1_STATE2_REG_1__SCAN_IN; 
assign P1_U3263 = ~P1_STATE2_REG_2__SCAN_IN; 
assign P1_U3264 = ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P1_U3265 = ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P1_U3266 = ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_U3268 = P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_U3269 = P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_U3270 = ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P1_U3275 = ~(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U3294 = ~P1_STATE2_REG_0__SCAN_IN; 
assign P1_U3296 = ~P1_STATE2_REG_3__SCAN_IN; 
assign P1_U3298 = P1_STATE2_REG_2__SCAN_IN | P1_STATE2_REG_1__SCAN_IN; 
assign P1_U3301 = ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN; 
assign P1_U3302 = ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign P1_U3303 = ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign P1_U3304 = ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P1_U3305 = ~(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P1_U3307 = P1_STATE2_REG_3__SCAN_IN | P1_STATE2_REG_2__SCAN_IN; 
assign P1_U3308 = ~P1_STATEBS16_REG_SCAN_IN; 
assign P1_U3387 = ~P1_FLUSH_REG_SCAN_IN; 
assign P1_U3413 = ~P1_REIP_REG_0__SCAN_IN; 
assign P1_U3429 = ~P1_EBX_REG_31__SCAN_IN; 
assign P1_U3435 = ~P1_CODEFETCH_REG_SCAN_IN; 
assign P1_U3436 = ~P1_READREQUEST_REG_SCAN_IN; 
assign P1_U3480 = ~(P1_DATAWIDTH_REG_1__SCAN_IN | P1_REIP_REG_1__SCAN_IN); 
assign P1_U3496 = P1_STATE_REG_0__SCAN_IN & P1_REQUESTPENDING_REG_SCAN_IN; 
assign P1_U3497 = ~(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_U3498 = P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_U3499 = ~(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U3500 = P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_U3501 = ~(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U3502 = P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P1_U3503 = ~(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U3504 = P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_U3505 = ~(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U3506 = P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P1_U3507 = P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P1_U3520 = ~(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U3521 = P1_INSTQUEUE_REG_5__5__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_U3522 = ~(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U3523 = P1_INSTQUEUE_REG_6__5__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P1_U3524 = P1_INSTQUEUE_REG_8__5__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P1_U3525 = ~(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U3526 = P1_INSTQUEUE_REG_10__5__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P1_U3527 = P1_INSTQUEUE_REG_12__5__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P1_U3528 = ~(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U3529 = P1_INSTQUEUE_REG_9__5__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_U3534 = ~(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_U3535 = P1_INSTQUEUE_REG_3__6__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_U3540 = ~(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_U3541 = P1_INSTQUEUE_REG_1__4__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_U3542 = ~(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U3543 = P1_INSTQUEUE_REG_4__4__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P1_U3544 = ~(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U3545 = P1_INSTQUEUE_REG_12__4__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P1_U3546 = P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_U3547 = P1_INSTQUEUE_REG_13__4__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P1_U3548 = ~(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U3549 = P1_INSTQUEUE_REG_6__4__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P1_U3550 = P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P1_U3551 = P1_INSTQUEUE_REG_14__4__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P1_U3552 = ~(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U3553 = P1_INSTQUEUE_REG_9__4__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P1_U3584 = P1_STATE2_REG_3__SCAN_IN & P1_STATE2_REG_0__SCAN_IN; 
assign P1_U3731 = P1_STATE2_REG_0__SCAN_IN & P1_FLUSH_REG_SCAN_IN; 
assign P1_U3864 = P1_STATE2_REG_1__SCAN_IN & P1_STATEBS16_REG_SCAN_IN; 
assign P1_U3950 = ~(P1_DATAWIDTH_REG_2__SCAN_IN | P1_DATAWIDTH_REG_3__SCAN_IN | P1_DATAWIDTH_REG_4__SCAN_IN | P1_DATAWIDTH_REG_5__SCAN_IN); 
assign P1_U3951 = ~(P1_DATAWIDTH_REG_6__SCAN_IN | P1_DATAWIDTH_REG_7__SCAN_IN | P1_DATAWIDTH_REG_8__SCAN_IN | P1_DATAWIDTH_REG_9__SCAN_IN); 
assign P1_U3953 = ~(P1_DATAWIDTH_REG_10__SCAN_IN | P1_DATAWIDTH_REG_11__SCAN_IN | P1_DATAWIDTH_REG_12__SCAN_IN | P1_DATAWIDTH_REG_13__SCAN_IN); 
assign P1_U3954 = ~(P1_DATAWIDTH_REG_14__SCAN_IN | P1_DATAWIDTH_REG_15__SCAN_IN | P1_DATAWIDTH_REG_16__SCAN_IN | P1_DATAWIDTH_REG_17__SCAN_IN); 
assign P1_U3956 = ~(P1_DATAWIDTH_REG_18__SCAN_IN | P1_DATAWIDTH_REG_19__SCAN_IN | P1_DATAWIDTH_REG_20__SCAN_IN | P1_DATAWIDTH_REG_21__SCAN_IN); 
assign P1_U3957 = ~(P1_DATAWIDTH_REG_22__SCAN_IN | P1_DATAWIDTH_REG_23__SCAN_IN | P1_DATAWIDTH_REG_24__SCAN_IN | P1_DATAWIDTH_REG_25__SCAN_IN); 
assign P1_U3959 = ~(P1_DATAWIDTH_REG_26__SCAN_IN | P1_DATAWIDTH_REG_27__SCAN_IN); 
assign P1_U3960 = ~(P1_DATAWIDTH_REG_28__SCAN_IN | P1_DATAWIDTH_REG_29__SCAN_IN); 
assign P1_U3961 = ~(P1_DATAWIDTH_REG_30__SCAN_IN | P1_DATAWIDTH_REG_31__SCAN_IN); 
assign P1_U3963 = ~(P1_DATAWIDTH_REG_0__SCAN_IN | P1_DATAWIDTH_REG_1__SCAN_IN | P1_REIP_REG_0__SCAN_IN); 
assign P1_U4174 = ~P1_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P1_U4179 = ~BS16; 
assign P1_U4362 = NA | P1_STATE_REG_0__SCAN_IN; 
assign P1_U4414 = ~(P1_INSTQUEUE_REG_15__5__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U4510 = P1_FLUSH_REG_SCAN_IN | P1_MORE_REG_SCAN_IN; 
assign P1_U5477 = ~(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U6598 = ~(P1_DATAWIDTH_REG_0__SCAN_IN & P1_DATAWIDTH_REG_1__SCAN_IN); 
assign P1_U6599 = P1_REIP_REG_0__SCAN_IN | P1_REIP_REG_1__SCAN_IN; 
assign P1_U6613 = ~(P1_STATE_REG_0__SCAN_IN & P1_ADS_N_REG_SCAN_IN); 
assign P1_U7648 = P1_STATE_REG_1__SCAN_IN | P1_STATE_REG_0__SCAN_IN; 
assign P1_U7664 = ~(P1_INSTQUEUE_REG_15__4__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U7687 = P1_STATE2_REG_0__SCAN_IN | P1_STATEBS16_REG_SCAN_IN; 
assign P1_U7714 = ~(P1_INSTADDRPOINTER_REG_0__SCAN_IN & P1_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P1_U7748 = P1_DATAWIDTH_REG_0__SCAN_IN | P1_DATAWIDTH_REG_1__SCAN_IN; 
assign P1_U7752 = ~(P1_REIP_REG_0__SCAN_IN & P1_REIP_REG_1__SCAN_IN); 
assign LT_782_120_U7 = ~P3_DATAO_REG_31__SCAN_IN; 
assign LT_782_U7 = ~P1_DATAO_REG_31__SCAN_IN; 
assign LT_748_U6 = ~P2_ADDRESS_REG_29__SCAN_IN; 
assign R170_U7 = P2_ADDRESS_REG_22__SCAN_IN | P2_ADDRESS_REG_17__SCAN_IN | P2_ADDRESS_REG_9__SCAN_IN | P2_ADDRESS_REG_7__SCAN_IN; 
assign R170_U9 = P2_ADDRESS_REG_18__SCAN_IN | P2_ADDRESS_REG_16__SCAN_IN | P2_ADDRESS_REG_8__SCAN_IN | P2_ADDRESS_REG_0__SCAN_IN; 
assign R170_U11 = P2_ADDRESS_REG_28__SCAN_IN | P2_ADDRESS_REG_26__SCAN_IN | P2_ADDRESS_REG_21__SCAN_IN | P2_ADDRESS_REG_6__SCAN_IN; 
assign R170_U13 = P2_ADDRESS_REG_27__SCAN_IN | P2_ADDRESS_REG_20__SCAN_IN | P2_ADDRESS_REG_13__SCAN_IN | P2_ADDRESS_REG_3__SCAN_IN; 
assign R165_U7 = P1_ADDRESS_REG_22__SCAN_IN | P1_ADDRESS_REG_17__SCAN_IN | P1_ADDRESS_REG_9__SCAN_IN | P1_ADDRESS_REG_7__SCAN_IN; 
assign R165_U9 = P1_ADDRESS_REG_18__SCAN_IN | P1_ADDRESS_REG_16__SCAN_IN | P1_ADDRESS_REG_8__SCAN_IN | P1_ADDRESS_REG_0__SCAN_IN; 
assign R165_U11 = P1_ADDRESS_REG_28__SCAN_IN | P1_ADDRESS_REG_26__SCAN_IN | P1_ADDRESS_REG_21__SCAN_IN | P1_ADDRESS_REG_6__SCAN_IN; 
assign R165_U13 = P1_ADDRESS_REG_27__SCAN_IN | P1_ADDRESS_REG_20__SCAN_IN | P1_ADDRESS_REG_13__SCAN_IN | P1_ADDRESS_REG_3__SCAN_IN; 
assign LT_782_119_U7 = ~P2_DATAO_REG_31__SCAN_IN; 
assign P3_ADD_526_U5 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P3_ADD_526_U6 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_526_U7 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_526_U8 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_526_U9 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_526_U10 = ~(P3_INSTADDRPOINTER_REG_0__SCAN_IN & P3_INSTADDRPOINTER_REG_1__SCAN_IN & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_526_U11 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_526_U12 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_526_U14 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_526_U15 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_526_U18 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_526_U19 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_526_U20 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_526_U21 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_526_U23 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_526_U24 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_526_U26 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_526_U28 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_526_U29 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_526_U30 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_526_U32 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_526_U33 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_526_U35 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_526_U37 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_526_U38 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_526_U39 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_526_U41 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_526_U42 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_526_U44 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_526_U45 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_526_U47 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_526_U50 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_526_U82 = P3_INSTADDRPOINTER_REG_3__SCAN_IN & P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_526_U83 = P3_INSTADDRPOINTER_REG_5__SCAN_IN & P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_526_U84 = P3_INSTADDRPOINTER_REG_7__SCAN_IN & P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_526_U85 = P3_INSTADDRPOINTER_REG_9__SCAN_IN & P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_526_U86 = P3_INSTADDRPOINTER_REG_11__SCAN_IN & P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_526_U87 = P3_INSTADDRPOINTER_REG_13__SCAN_IN & P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_526_U88 = P3_INSTADDRPOINTER_REG_15__SCAN_IN & P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_526_U89 = P3_INSTADDRPOINTER_REG_17__SCAN_IN & P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_526_U90 = P3_INSTADDRPOINTER_REG_19__SCAN_IN & P3_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_526_U91 = P3_INSTADDRPOINTER_REG_21__SCAN_IN & P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_526_U92 = P3_INSTADDRPOINTER_REG_23__SCAN_IN & P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_526_U93 = P3_INSTADDRPOINTER_REG_25__SCAN_IN & P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_526_U94 = P3_INSTADDRPOINTER_REG_27__SCAN_IN & P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_526_U98 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_ADD_526_U100 = ~(P3_INSTADDRPOINTER_REG_0__SCAN_IN & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_552_U5 = ~P3_EBX_REG_0__SCAN_IN; 
assign P3_ADD_552_U6 = ~P3_EBX_REG_2__SCAN_IN; 
assign P3_ADD_552_U7 = ~P3_EBX_REG_1__SCAN_IN; 
assign P3_ADD_552_U8 = ~P3_EBX_REG_4__SCAN_IN; 
assign P3_ADD_552_U9 = ~P3_EBX_REG_3__SCAN_IN; 
assign P3_ADD_552_U10 = ~(P3_EBX_REG_0__SCAN_IN & P3_EBX_REG_1__SCAN_IN & P3_EBX_REG_2__SCAN_IN); 
assign P3_ADD_552_U11 = ~P3_EBX_REG_6__SCAN_IN; 
assign P3_ADD_552_U12 = ~P3_EBX_REG_5__SCAN_IN; 
assign P3_ADD_552_U14 = ~P3_EBX_REG_8__SCAN_IN; 
assign P3_ADD_552_U15 = ~P3_EBX_REG_7__SCAN_IN; 
assign P3_ADD_552_U18 = ~P3_EBX_REG_9__SCAN_IN; 
assign P3_ADD_552_U19 = ~P3_EBX_REG_10__SCAN_IN; 
assign P3_ADD_552_U20 = ~P3_EBX_REG_12__SCAN_IN; 
assign P3_ADD_552_U21 = ~P3_EBX_REG_11__SCAN_IN; 
assign P3_ADD_552_U23 = ~P3_EBX_REG_14__SCAN_IN; 
assign P3_ADD_552_U24 = ~P3_EBX_REG_13__SCAN_IN; 
assign P3_ADD_552_U26 = ~P3_EBX_REG_15__SCAN_IN; 
assign P3_ADD_552_U28 = ~P3_EBX_REG_16__SCAN_IN; 
assign P3_ADD_552_U29 = ~P3_EBX_REG_18__SCAN_IN; 
assign P3_ADD_552_U30 = ~P3_EBX_REG_17__SCAN_IN; 
assign P3_ADD_552_U32 = ~P3_EBX_REG_20__SCAN_IN; 
assign P3_ADD_552_U33 = ~P3_EBX_REG_19__SCAN_IN; 
assign P3_ADD_552_U35 = ~P3_EBX_REG_21__SCAN_IN; 
assign P3_ADD_552_U37 = ~P3_EBX_REG_22__SCAN_IN; 
assign P3_ADD_552_U38 = ~P3_EBX_REG_24__SCAN_IN; 
assign P3_ADD_552_U39 = ~P3_EBX_REG_23__SCAN_IN; 
assign P3_ADD_552_U41 = ~P3_EBX_REG_26__SCAN_IN; 
assign P3_ADD_552_U42 = ~P3_EBX_REG_25__SCAN_IN; 
assign P3_ADD_552_U44 = ~P3_EBX_REG_27__SCAN_IN; 
assign P3_ADD_552_U45 = ~P3_EBX_REG_28__SCAN_IN; 
assign P3_ADD_552_U47 = ~P3_EBX_REG_29__SCAN_IN; 
assign P3_ADD_552_U50 = ~P3_EBX_REG_30__SCAN_IN; 
assign P3_ADD_552_U82 = P3_EBX_REG_3__SCAN_IN & P3_EBX_REG_4__SCAN_IN; 
assign P3_ADD_552_U83 = P3_EBX_REG_5__SCAN_IN & P3_EBX_REG_6__SCAN_IN; 
assign P3_ADD_552_U84 = P3_EBX_REG_7__SCAN_IN & P3_EBX_REG_8__SCAN_IN; 
assign P3_ADD_552_U85 = P3_EBX_REG_9__SCAN_IN & P3_EBX_REG_10__SCAN_IN; 
assign P3_ADD_552_U86 = P3_EBX_REG_11__SCAN_IN & P3_EBX_REG_12__SCAN_IN; 
assign P3_ADD_552_U87 = P3_EBX_REG_13__SCAN_IN & P3_EBX_REG_14__SCAN_IN; 
assign P3_ADD_552_U88 = P3_EBX_REG_15__SCAN_IN & P3_EBX_REG_16__SCAN_IN; 
assign P3_ADD_552_U89 = P3_EBX_REG_17__SCAN_IN & P3_EBX_REG_18__SCAN_IN; 
assign P3_ADD_552_U90 = P3_EBX_REG_19__SCAN_IN & P3_EBX_REG_20__SCAN_IN; 
assign P3_ADD_552_U91 = P3_EBX_REG_21__SCAN_IN & P3_EBX_REG_22__SCAN_IN; 
assign P3_ADD_552_U92 = P3_EBX_REG_23__SCAN_IN & P3_EBX_REG_24__SCAN_IN; 
assign P3_ADD_552_U93 = P3_EBX_REG_25__SCAN_IN & P3_EBX_REG_26__SCAN_IN; 
assign P3_ADD_552_U94 = P3_EBX_REG_27__SCAN_IN & P3_EBX_REG_28__SCAN_IN; 
assign P3_ADD_552_U98 = ~P3_EBX_REG_31__SCAN_IN; 
assign P3_ADD_552_U100 = ~(P3_EBX_REG_0__SCAN_IN & P3_EBX_REG_1__SCAN_IN); 
assign P3_ADD_546_U5 = ~P3_EAX_REG_0__SCAN_IN; 
assign P3_ADD_546_U6 = ~P3_EAX_REG_2__SCAN_IN; 
assign P3_ADD_546_U7 = ~P3_EAX_REG_1__SCAN_IN; 
assign P3_ADD_546_U8 = ~P3_EAX_REG_4__SCAN_IN; 
assign P3_ADD_546_U9 = ~P3_EAX_REG_3__SCAN_IN; 
assign P3_ADD_546_U10 = ~(P3_EAX_REG_0__SCAN_IN & P3_EAX_REG_1__SCAN_IN & P3_EAX_REG_2__SCAN_IN); 
assign P3_ADD_546_U11 = ~P3_EAX_REG_6__SCAN_IN; 
assign P3_ADD_546_U12 = ~P3_EAX_REG_5__SCAN_IN; 
assign P3_ADD_546_U14 = ~P3_EAX_REG_8__SCAN_IN; 
assign P3_ADD_546_U15 = ~P3_EAX_REG_7__SCAN_IN; 
assign P3_ADD_546_U18 = ~P3_EAX_REG_9__SCAN_IN; 
assign P3_ADD_546_U19 = ~P3_EAX_REG_10__SCAN_IN; 
assign P3_ADD_546_U20 = ~P3_EAX_REG_12__SCAN_IN; 
assign P3_ADD_546_U21 = ~P3_EAX_REG_11__SCAN_IN; 
assign P3_ADD_546_U23 = ~P3_EAX_REG_14__SCAN_IN; 
assign P3_ADD_546_U24 = ~P3_EAX_REG_13__SCAN_IN; 
assign P3_ADD_546_U26 = ~P3_EAX_REG_15__SCAN_IN; 
assign P3_ADD_546_U28 = ~P3_EAX_REG_16__SCAN_IN; 
assign P3_ADD_546_U29 = ~P3_EAX_REG_18__SCAN_IN; 
assign P3_ADD_546_U30 = ~P3_EAX_REG_17__SCAN_IN; 
assign P3_ADD_546_U32 = ~P3_EAX_REG_20__SCAN_IN; 
assign P3_ADD_546_U33 = ~P3_EAX_REG_19__SCAN_IN; 
assign P3_ADD_546_U35 = ~P3_EAX_REG_21__SCAN_IN; 
assign P3_ADD_546_U37 = ~P3_EAX_REG_22__SCAN_IN; 
assign P3_ADD_546_U38 = ~P3_EAX_REG_24__SCAN_IN; 
assign P3_ADD_546_U39 = ~P3_EAX_REG_23__SCAN_IN; 
assign P3_ADD_546_U41 = ~P3_EAX_REG_26__SCAN_IN; 
assign P3_ADD_546_U42 = ~P3_EAX_REG_25__SCAN_IN; 
assign P3_ADD_546_U44 = ~P3_EAX_REG_27__SCAN_IN; 
assign P3_ADD_546_U45 = ~P3_EAX_REG_28__SCAN_IN; 
assign P3_ADD_546_U47 = ~P3_EAX_REG_29__SCAN_IN; 
assign P3_ADD_546_U50 = ~P3_EAX_REG_30__SCAN_IN; 
assign P3_ADD_546_U82 = P3_EAX_REG_3__SCAN_IN & P3_EAX_REG_4__SCAN_IN; 
assign P3_ADD_546_U83 = P3_EAX_REG_5__SCAN_IN & P3_EAX_REG_6__SCAN_IN; 
assign P3_ADD_546_U84 = P3_EAX_REG_7__SCAN_IN & P3_EAX_REG_8__SCAN_IN; 
assign P3_ADD_546_U85 = P3_EAX_REG_9__SCAN_IN & P3_EAX_REG_10__SCAN_IN; 
assign P3_ADD_546_U86 = P3_EAX_REG_11__SCAN_IN & P3_EAX_REG_12__SCAN_IN; 
assign P3_ADD_546_U87 = P3_EAX_REG_13__SCAN_IN & P3_EAX_REG_14__SCAN_IN; 
assign P3_ADD_546_U88 = P3_EAX_REG_15__SCAN_IN & P3_EAX_REG_16__SCAN_IN; 
assign P3_ADD_546_U89 = P3_EAX_REG_17__SCAN_IN & P3_EAX_REG_18__SCAN_IN; 
assign P3_ADD_546_U90 = P3_EAX_REG_19__SCAN_IN & P3_EAX_REG_20__SCAN_IN; 
assign P3_ADD_546_U91 = P3_EAX_REG_21__SCAN_IN & P3_EAX_REG_22__SCAN_IN; 
assign P3_ADD_546_U92 = P3_EAX_REG_23__SCAN_IN & P3_EAX_REG_24__SCAN_IN; 
assign P3_ADD_546_U93 = P3_EAX_REG_25__SCAN_IN & P3_EAX_REG_26__SCAN_IN; 
assign P3_ADD_546_U94 = P3_EAX_REG_27__SCAN_IN & P3_EAX_REG_28__SCAN_IN; 
assign P3_ADD_546_U98 = ~P3_EAX_REG_31__SCAN_IN; 
assign P3_ADD_546_U100 = ~(P3_EAX_REG_0__SCAN_IN & P3_EAX_REG_1__SCAN_IN); 
assign P3_ADD_476_U4 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_476_U5 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_476_U6 = ~(P3_INSTADDRPOINTER_REG_1__SCAN_IN & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_476_U7 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_476_U9 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_476_U11 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_476_U13 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_476_U15 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_476_U17 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_476_U18 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_476_U21 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_476_U23 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_476_U25 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_476_U27 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_476_U29 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_476_U31 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_476_U33 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_476_U35 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_476_U37 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_476_U39 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_476_U41 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_476_U43 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_476_U45 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_476_U47 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_476_U49 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_476_U51 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_476_U53 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_476_U55 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_476_U57 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_476_U59 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_476_U61 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_476_U92 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_ADD_531_U5 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P3_ADD_531_U6 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_531_U7 = ~(P3_INSTADDRPOINTER_REG_0__SCAN_IN & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_531_U8 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_531_U10 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_531_U12 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_531_U14 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_531_U16 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_531_U18 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_531_U20 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_531_U21 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_531_U24 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_531_U26 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_531_U28 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_531_U30 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_531_U32 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_531_U34 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_531_U36 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_531_U38 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_531_U40 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_531_U42 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_531_U44 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_531_U46 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_531_U48 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_531_U50 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_531_U52 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_531_U54 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_531_U56 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_531_U58 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_531_U60 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_531_U62 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_531_U64 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_531_U96 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_SUB_320_U72 = ~P3_PHYADDRPOINTER_REG_0__SCAN_IN; 
assign P3_ADD_505_U5 = ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P3_ADD_505_U7 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P3_ADD_505_U8 = ~(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P3_ADD_505_U9 = ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P3_ADD_505_U11 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P3_ADD_505_U13 = ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P3_ADD_318_U4 = ~P3_PHYADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_318_U5 = ~P3_PHYADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_318_U6 = ~(P3_PHYADDRPOINTER_REG_1__SCAN_IN & P3_PHYADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_318_U7 = ~P3_PHYADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_318_U9 = ~P3_PHYADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_318_U11 = ~P3_PHYADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_318_U13 = ~P3_PHYADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_318_U15 = ~P3_PHYADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_318_U17 = ~P3_PHYADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_318_U18 = ~P3_PHYADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_318_U21 = ~P3_PHYADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_318_U23 = ~P3_PHYADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_318_U25 = ~P3_PHYADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_318_U27 = ~P3_PHYADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_318_U29 = ~P3_PHYADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_318_U31 = ~P3_PHYADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_318_U33 = ~P3_PHYADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_318_U35 = ~P3_PHYADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_318_U37 = ~P3_PHYADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_318_U39 = ~P3_PHYADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_318_U41 = ~P3_PHYADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_318_U43 = ~P3_PHYADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_318_U45 = ~P3_PHYADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_318_U47 = ~P3_PHYADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_318_U49 = ~P3_PHYADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_318_U51 = ~P3_PHYADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_318_U53 = ~P3_PHYADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_318_U55 = ~P3_PHYADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_318_U57 = ~P3_PHYADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_318_U59 = ~P3_PHYADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_318_U61 = ~P3_PHYADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_318_U92 = ~P3_PHYADDRPOINTER_REG_31__SCAN_IN; 
assign P3_SUB_370_U8 = ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P3_SUB_370_U10 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign P3_SUB_370_U11 = ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P3_SUB_370_U12 = ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P3_SUB_370_U13 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P3_SUB_370_U14 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign P3_SUB_370_U15 = ~P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign P3_SUB_370_U17 = ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P3_SUB_370_U18 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN; 
assign P3_SUB_370_U29 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P3_ADD_315_U4 = ~P3_PHYADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_315_U5 = ~P3_PHYADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_315_U6 = ~(P3_PHYADDRPOINTER_REG_2__SCAN_IN & P3_PHYADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_315_U7 = ~P3_PHYADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_315_U9 = ~P3_PHYADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_315_U11 = ~P3_PHYADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_315_U13 = ~P3_PHYADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_315_U15 = ~P3_PHYADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_315_U16 = ~P3_PHYADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_315_U19 = ~P3_PHYADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_315_U21 = ~P3_PHYADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_315_U23 = ~P3_PHYADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_315_U25 = ~P3_PHYADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_315_U27 = ~P3_PHYADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_315_U29 = ~P3_PHYADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_315_U31 = ~P3_PHYADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_315_U33 = ~P3_PHYADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_315_U35 = ~P3_PHYADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_315_U37 = ~P3_PHYADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_315_U39 = ~P3_PHYADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_315_U41 = ~P3_PHYADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_315_U43 = ~P3_PHYADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_315_U45 = ~P3_PHYADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_315_U47 = ~P3_PHYADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_315_U49 = ~P3_PHYADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_315_U51 = ~P3_PHYADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_315_U53 = ~P3_PHYADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_315_U55 = ~P3_PHYADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_315_U57 = ~P3_PHYADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_315_U59 = ~P3_PHYADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_315_U89 = ~P3_PHYADDRPOINTER_REG_31__SCAN_IN; 
assign P3_ADD_360_1242_U21 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_360_1242_U23 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_360_1242_U25 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P3_ADD_360_1242_U26 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_360_1242_U30 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_360_1242_U31 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_360_1242_U34 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_360_1242_U35 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_360_1242_U38 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_360_1242_U39 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_360_1242_U42 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_360_1242_U43 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_360_1242_U44 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_360_1242_U47 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_360_1242_U48 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_360_1242_U49 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_360_1242_U51 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_360_1242_U52 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_360_1242_U54 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_360_1242_U55 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_360_1242_U57 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_360_1242_U59 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_360_1242_U61 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_360_1242_U62 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_360_1242_U64 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_360_1242_U65 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_360_1242_U67 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_360_1242_U69 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_360_1242_U70 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_360_1242_U72 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_360_1242_U74 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_360_1242_U97 = P3_INSTADDRPOINTER_REG_9__SCAN_IN & P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_360_1242_U98 = P3_INSTADDRPOINTER_REG_11__SCAN_IN & P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_360_1242_U99 = P3_INSTADDRPOINTER_REG_13__SCAN_IN & P3_INSTADDRPOINTER_REG_14__SCAN_IN & P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_360_1242_U100 = P3_INSTADDRPOINTER_REG_16__SCAN_IN & P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_360_1242_U101 = P3_INSTADDRPOINTER_REG_18__SCAN_IN & P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_360_1242_U102 = P3_INSTADDRPOINTER_REG_22__SCAN_IN & P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_360_1242_U103 = P3_INSTADDRPOINTER_REG_24__SCAN_IN & P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_360_1242_U104 = P3_INSTADDRPOINTER_REG_27__SCAN_IN & P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_360_1242_U116 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_ADD_467_U4 = ~P3_REIP_REG_1__SCAN_IN; 
assign P3_ADD_467_U5 = ~P3_REIP_REG_2__SCAN_IN; 
assign P3_ADD_467_U6 = ~(P3_REIP_REG_1__SCAN_IN & P3_REIP_REG_2__SCAN_IN); 
assign P3_ADD_467_U7 = ~P3_REIP_REG_3__SCAN_IN; 
assign P3_ADD_467_U9 = ~P3_REIP_REG_4__SCAN_IN; 
assign P3_ADD_467_U11 = ~P3_REIP_REG_5__SCAN_IN; 
assign P3_ADD_467_U13 = ~P3_REIP_REG_6__SCAN_IN; 
assign P3_ADD_467_U15 = ~P3_REIP_REG_7__SCAN_IN; 
assign P3_ADD_467_U17 = ~P3_REIP_REG_8__SCAN_IN; 
assign P3_ADD_467_U18 = ~P3_REIP_REG_9__SCAN_IN; 
assign P3_ADD_467_U21 = ~P3_REIP_REG_10__SCAN_IN; 
assign P3_ADD_467_U23 = ~P3_REIP_REG_11__SCAN_IN; 
assign P3_ADD_467_U25 = ~P3_REIP_REG_12__SCAN_IN; 
assign P3_ADD_467_U27 = ~P3_REIP_REG_13__SCAN_IN; 
assign P3_ADD_467_U29 = ~P3_REIP_REG_14__SCAN_IN; 
assign P3_ADD_467_U31 = ~P3_REIP_REG_15__SCAN_IN; 
assign P3_ADD_467_U33 = ~P3_REIP_REG_16__SCAN_IN; 
assign P3_ADD_467_U35 = ~P3_REIP_REG_17__SCAN_IN; 
assign P3_ADD_467_U37 = ~P3_REIP_REG_18__SCAN_IN; 
assign P3_ADD_467_U39 = ~P3_REIP_REG_19__SCAN_IN; 
assign P3_ADD_467_U41 = ~P3_REIP_REG_20__SCAN_IN; 
assign P3_ADD_467_U43 = ~P3_REIP_REG_21__SCAN_IN; 
assign P3_ADD_467_U45 = ~P3_REIP_REG_22__SCAN_IN; 
assign P3_ADD_467_U47 = ~P3_REIP_REG_23__SCAN_IN; 
assign P3_ADD_467_U49 = ~P3_REIP_REG_24__SCAN_IN; 
assign P3_ADD_467_U51 = ~P3_REIP_REG_25__SCAN_IN; 
assign P3_ADD_467_U53 = ~P3_REIP_REG_26__SCAN_IN; 
assign P3_ADD_467_U55 = ~P3_REIP_REG_27__SCAN_IN; 
assign P3_ADD_467_U57 = ~P3_REIP_REG_28__SCAN_IN; 
assign P3_ADD_467_U59 = ~P3_REIP_REG_29__SCAN_IN; 
assign P3_ADD_467_U61 = ~P3_REIP_REG_30__SCAN_IN; 
assign P3_ADD_467_U92 = ~P3_REIP_REG_31__SCAN_IN; 
assign P3_ADD_430_U4 = ~P3_REIP_REG_1__SCAN_IN; 
assign P3_ADD_430_U5 = ~P3_REIP_REG_2__SCAN_IN; 
assign P3_ADD_430_U6 = ~(P3_REIP_REG_1__SCAN_IN & P3_REIP_REG_2__SCAN_IN); 
assign P3_ADD_430_U7 = ~P3_REIP_REG_3__SCAN_IN; 
assign P3_ADD_430_U9 = ~P3_REIP_REG_4__SCAN_IN; 
assign P3_ADD_430_U11 = ~P3_REIP_REG_5__SCAN_IN; 
assign P3_ADD_430_U13 = ~P3_REIP_REG_6__SCAN_IN; 
assign P3_ADD_430_U15 = ~P3_REIP_REG_7__SCAN_IN; 
assign P3_ADD_430_U17 = ~P3_REIP_REG_8__SCAN_IN; 
assign P3_ADD_430_U18 = ~P3_REIP_REG_9__SCAN_IN; 
assign P3_ADD_430_U21 = ~P3_REIP_REG_10__SCAN_IN; 
assign P3_ADD_430_U23 = ~P3_REIP_REG_11__SCAN_IN; 
assign P3_ADD_430_U25 = ~P3_REIP_REG_12__SCAN_IN; 
assign P3_ADD_430_U27 = ~P3_REIP_REG_13__SCAN_IN; 
assign P3_ADD_430_U29 = ~P3_REIP_REG_14__SCAN_IN; 
assign P3_ADD_430_U31 = ~P3_REIP_REG_15__SCAN_IN; 
assign P3_ADD_430_U33 = ~P3_REIP_REG_16__SCAN_IN; 
assign P3_ADD_430_U35 = ~P3_REIP_REG_17__SCAN_IN; 
assign P3_ADD_430_U37 = ~P3_REIP_REG_18__SCAN_IN; 
assign P3_ADD_430_U39 = ~P3_REIP_REG_19__SCAN_IN; 
assign P3_ADD_430_U41 = ~P3_REIP_REG_20__SCAN_IN; 
assign P3_ADD_430_U43 = ~P3_REIP_REG_21__SCAN_IN; 
assign P3_ADD_430_U45 = ~P3_REIP_REG_22__SCAN_IN; 
assign P3_ADD_430_U47 = ~P3_REIP_REG_23__SCAN_IN; 
assign P3_ADD_430_U49 = ~P3_REIP_REG_24__SCAN_IN; 
assign P3_ADD_430_U51 = ~P3_REIP_REG_25__SCAN_IN; 
assign P3_ADD_430_U53 = ~P3_REIP_REG_26__SCAN_IN; 
assign P3_ADD_430_U55 = ~P3_REIP_REG_27__SCAN_IN; 
assign P3_ADD_430_U57 = ~P3_REIP_REG_28__SCAN_IN; 
assign P3_ADD_430_U59 = ~P3_REIP_REG_29__SCAN_IN; 
assign P3_ADD_430_U61 = ~P3_REIP_REG_30__SCAN_IN; 
assign P3_ADD_430_U92 = ~P3_REIP_REG_31__SCAN_IN; 
assign P3_ADD_380_U5 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P3_ADD_380_U6 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_380_U7 = ~(P3_INSTADDRPOINTER_REG_0__SCAN_IN & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_380_U8 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_380_U10 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_380_U12 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_380_U14 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_380_U16 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_380_U18 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_380_U20 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_380_U21 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_380_U24 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_380_U26 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_380_U28 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_380_U30 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_380_U32 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_380_U34 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_380_U36 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_380_U38 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_380_U40 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_380_U42 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_380_U44 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_380_U46 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_380_U48 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_380_U50 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_380_U52 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_380_U54 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_380_U56 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_380_U58 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_380_U60 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_380_U62 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_380_U64 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_380_U96 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_ADD_344_U5 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P3_ADD_344_U6 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_344_U7 = ~(P3_INSTADDRPOINTER_REG_0__SCAN_IN & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_344_U8 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_344_U10 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_344_U12 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_344_U14 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_344_U16 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_344_U18 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_344_U20 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_344_U21 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_344_U24 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_344_U26 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_344_U28 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_344_U30 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_344_U32 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_344_U34 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_344_U36 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_344_U38 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_344_U40 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_344_U42 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_344_U44 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_344_U46 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_344_U48 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_344_U50 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_344_U52 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_344_U54 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_344_U56 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_344_U58 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_344_U60 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_344_U62 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_344_U64 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_344_U96 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_LT_563_U7 = ~P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign P3_LT_563_U9 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign P3_LT_563_U11 = ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P3_LT_563_U12 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign P3_ADD_339_U4 = ~P3_PHYADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_339_U5 = ~P3_PHYADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_339_U6 = ~(P3_PHYADDRPOINTER_REG_1__SCAN_IN & P3_PHYADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_339_U7 = ~P3_PHYADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_339_U9 = ~P3_PHYADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_339_U11 = ~P3_PHYADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_339_U13 = ~P3_PHYADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_339_U15 = ~P3_PHYADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_339_U17 = ~P3_PHYADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_339_U18 = ~P3_PHYADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_339_U21 = ~P3_PHYADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_339_U23 = ~P3_PHYADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_339_U25 = ~P3_PHYADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_339_U27 = ~P3_PHYADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_339_U29 = ~P3_PHYADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_339_U31 = ~P3_PHYADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_339_U33 = ~P3_PHYADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_339_U35 = ~P3_PHYADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_339_U37 = ~P3_PHYADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_339_U39 = ~P3_PHYADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_339_U41 = ~P3_PHYADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_339_U43 = ~P3_PHYADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_339_U45 = ~P3_PHYADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_339_U47 = ~P3_PHYADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_339_U49 = ~P3_PHYADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_339_U51 = ~P3_PHYADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_339_U53 = ~P3_PHYADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_339_U55 = ~P3_PHYADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_339_U57 = ~P3_PHYADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_339_U59 = ~P3_PHYADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_339_U61 = ~P3_PHYADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_339_U92 = ~P3_PHYADDRPOINTER_REG_31__SCAN_IN; 
assign P3_LTE_597_U6 = ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P3_SUB_580_U7 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_SUB_580_U8 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P3_ADD_541_U4 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_541_U5 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_541_U6 = ~(P3_INSTADDRPOINTER_REG_1__SCAN_IN & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_541_U7 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_541_U9 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_541_U11 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_541_U13 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_541_U15 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_541_U17 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_541_U18 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_541_U21 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_541_U23 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_541_U25 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_541_U27 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_541_U29 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_541_U31 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_541_U33 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_541_U35 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_541_U37 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_541_U39 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_541_U41 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_541_U43 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_541_U45 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_541_U47 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_541_U49 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_541_U51 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_541_U53 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_541_U55 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_541_U57 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_541_U59 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_541_U61 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_541_U92 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_SUB_355_U8 = ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P3_SUB_355_U10 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign P3_SUB_355_U11 = ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P3_SUB_355_U12 = ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P3_SUB_355_U13 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P3_SUB_355_U14 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign P3_SUB_355_U15 = ~P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign P3_SUB_355_U17 = ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P3_SUB_355_U18 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN; 
assign P3_SUB_355_U29 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P3_SUB_450_U8 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign P3_SUB_450_U9 = ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P3_SUB_450_U10 = ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P3_SUB_450_U11 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P3_SUB_450_U12 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign P3_SUB_450_U13 = ~P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign P3_SUB_450_U15 = ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P3_SUB_450_U26 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P3_SUB_450_U27 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN; 
assign P3_SUB_357_1258_U4 = P3_INSTADDRPOINTER_REG_27__SCAN_IN & P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_SUB_357_1258_U23 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_SUB_357_1258_U25 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_SUB_357_1258_U27 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_SUB_357_1258_U29 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P3_SUB_357_1258_U33 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_SUB_357_1258_U34 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_SUB_357_1258_U36 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_SUB_357_1258_U38 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_SUB_357_1258_U40 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_SUB_357_1258_U41 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_SUB_357_1258_U42 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_SUB_357_1258_U43 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_SUB_357_1258_U44 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_SUB_357_1258_U45 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_SUB_357_1258_U46 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_SUB_357_1258_U47 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_SUB_357_1258_U48 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_SUB_357_1258_U49 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_SUB_357_1258_U50 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_SUB_357_1258_U51 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P3_SUB_357_1258_U52 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_SUB_357_1258_U53 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_SUB_357_1258_U54 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_SUB_357_1258_U55 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_SUB_357_1258_U56 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_SUB_357_1258_U57 = ~(P3_INSTADDRPOINTER_REG_19__SCAN_IN & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_SUB_357_1258_U58 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P3_SUB_357_1258_U59 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P3_SUB_357_1258_U60 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P3_SUB_357_1258_U101 = P3_INSTADDRPOINTER_REG_16__SCAN_IN & P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_SUB_357_1258_U108 = P3_INSTADDRPOINTER_REG_30__SCAN_IN & P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_SUB_357_1258_U191 = ~(P3_INSTADDRPOINTER_REG_12__SCAN_IN & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_SUB_357_1258_U217 = ~(P3_INSTADDRPOINTER_REG_25__SCAN_IN & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_486_U5 = ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P3_ADD_486_U7 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P3_ADD_486_U8 = ~(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P3_ADD_486_U9 = ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P3_ADD_486_U11 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P3_ADD_486_U13 = ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P3_SUB_485_U8 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign P3_SUB_485_U9 = ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P3_SUB_485_U10 = ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P3_SUB_485_U11 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P3_SUB_485_U12 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign P3_SUB_485_U13 = ~P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign P3_SUB_485_U15 = ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P3_SUB_485_U26 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P3_SUB_485_U27 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN; 
assign P3_ADD_515_U4 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_515_U5 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_515_U6 = ~(P3_INSTADDRPOINTER_REG_1__SCAN_IN & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_515_U7 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_515_U9 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_515_U11 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_515_U13 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_515_U15 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_515_U17 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_515_U18 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_515_U21 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_515_U23 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_515_U25 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_515_U27 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_515_U29 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_515_U31 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_515_U33 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_515_U35 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_515_U37 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_515_U39 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_515_U41 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_515_U43 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_515_U45 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_515_U47 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_515_U49 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_515_U51 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_515_U53 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_515_U55 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_515_U57 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_515_U59 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_515_U61 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_515_U92 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_ADD_394_U4 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P3_ADD_394_U6 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_394_U7 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_394_U9 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_394_U11 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_394_U13 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_394_U15 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_394_U17 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_394_U18 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_394_U21 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_394_U23 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_394_U25 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_394_U27 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_394_U29 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_394_U31 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_394_U33 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_394_U35 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_394_U37 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_394_U39 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_394_U41 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_394_U43 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_394_U45 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_394_U47 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_394_U49 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_394_U51 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_394_U53 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_394_U55 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_394_U57 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_394_U59 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_394_U61 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_394_U62 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_394_U94 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_ADD_394_U96 = ~(P3_INSTADDRPOINTER_REG_0__SCAN_IN & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_394_U126 = ~(P3_INSTADDRPOINTER_REG_0__SCAN_IN & P3_INSTADDRPOINTER_REG_1__SCAN_IN & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_SUB_414_U21 = P3_EBX_REG_0__SCAN_IN | P3_EBX_REG_1__SCAN_IN | P3_EBX_REG_2__SCAN_IN; 
assign P3_SUB_414_U25 = ~P3_EBX_REG_8__SCAN_IN; 
assign P3_SUB_414_U26 = ~P3_EBX_REG_6__SCAN_IN; 
assign P3_SUB_414_U27 = ~P3_EBX_REG_4__SCAN_IN; 
assign P3_SUB_414_U39 = ~P3_EBX_REG_29__SCAN_IN; 
assign P3_SUB_414_U40 = ~P3_EBX_REG_28__SCAN_IN; 
assign P3_SUB_414_U41 = ~P3_EBX_REG_26__SCAN_IN; 
assign P3_SUB_414_U42 = ~P3_EBX_REG_24__SCAN_IN; 
assign P3_SUB_414_U43 = ~P3_EBX_REG_22__SCAN_IN; 
assign P3_SUB_414_U44 = ~P3_EBX_REG_20__SCAN_IN; 
assign P3_SUB_414_U45 = ~P3_EBX_REG_18__SCAN_IN; 
assign P3_SUB_414_U46 = ~P3_EBX_REG_16__SCAN_IN; 
assign P3_SUB_414_U47 = ~P3_EBX_REG_14__SCAN_IN; 
assign P3_SUB_414_U48 = ~P3_EBX_REG_12__SCAN_IN; 
assign P3_SUB_414_U49 = ~P3_EBX_REG_10__SCAN_IN; 
assign P3_SUB_414_U52 = ~P3_EBX_REG_9__SCAN_IN; 
assign P3_SUB_414_U54 = ~P3_EBX_REG_7__SCAN_IN; 
assign P3_SUB_414_U56 = ~P3_EBX_REG_5__SCAN_IN; 
assign P3_SUB_414_U58 = ~P3_EBX_REG_3__SCAN_IN; 
assign P3_SUB_414_U60 = ~P3_EBX_REG_31__SCAN_IN; 
assign P3_SUB_414_U61 = ~P3_EBX_REG_30__SCAN_IN; 
assign P3_SUB_414_U63 = ~P3_EBX_REG_27__SCAN_IN; 
assign P3_SUB_414_U65 = ~P3_EBX_REG_25__SCAN_IN; 
assign P3_SUB_414_U67 = ~P3_EBX_REG_23__SCAN_IN; 
assign P3_SUB_414_U69 = ~P3_EBX_REG_21__SCAN_IN; 
assign P3_SUB_414_U71 = ~P3_EBX_REG_1__SCAN_IN; 
assign P3_SUB_414_U72 = ~P3_EBX_REG_0__SCAN_IN; 
assign P3_SUB_414_U73 = ~P3_EBX_REG_19__SCAN_IN; 
assign P3_SUB_414_U75 = ~P3_EBX_REG_17__SCAN_IN; 
assign P3_SUB_414_U77 = ~P3_EBX_REG_15__SCAN_IN; 
assign P3_SUB_414_U79 = ~P3_EBX_REG_13__SCAN_IN; 
assign P3_SUB_414_U81 = ~P3_EBX_REG_11__SCAN_IN; 
assign P3_SUB_414_U104 = P3_EBX_REG_0__SCAN_IN | P3_EBX_REG_1__SCAN_IN; 
assign P3_ADD_441_U4 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_441_U5 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_441_U6 = ~(P3_INSTADDRPOINTER_REG_1__SCAN_IN & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_441_U7 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_441_U9 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_441_U11 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_441_U13 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_441_U15 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_441_U17 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_441_U18 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_441_U21 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_441_U23 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_441_U25 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_441_U27 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_441_U29 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_441_U31 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_441_U33 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_441_U35 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_441_U37 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_441_U39 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_441_U41 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_441_U43 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_441_U45 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_441_U47 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_441_U49 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_441_U51 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_441_U53 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_441_U55 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_441_U57 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_441_U59 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_441_U61 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_441_U92 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_ADD_349_U5 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P3_ADD_349_U6 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_349_U7 = ~(P3_INSTADDRPOINTER_REG_0__SCAN_IN & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_349_U8 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_349_U10 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_349_U12 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_349_U14 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_349_U16 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_349_U18 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_349_U20 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_349_U21 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_349_U24 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_349_U26 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_349_U28 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_349_U30 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_349_U32 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_349_U34 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_349_U36 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_349_U38 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_349_U40 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_349_U42 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_349_U44 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_349_U46 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_349_U48 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_349_U50 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_349_U52 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_349_U54 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_349_U56 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_349_U58 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_349_U60 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_349_U62 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_349_U64 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_349_U96 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_ADD_405_U4 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P3_ADD_405_U6 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_405_U7 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_405_U9 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_405_U11 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_405_U13 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_405_U15 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_405_U17 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_405_U18 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_405_U21 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_405_U23 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_405_U25 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_405_U27 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_405_U29 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_405_U31 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_405_U33 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_405_U35 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_405_U37 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_405_U39 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_405_U41 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_405_U43 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_405_U45 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_405_U47 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_405_U49 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_405_U51 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_405_U53 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_405_U55 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_405_U57 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_405_U59 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_405_U61 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_405_U62 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_405_U94 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_ADD_405_U96 = ~(P3_INSTADDRPOINTER_REG_0__SCAN_IN & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_405_U126 = ~(P3_INSTADDRPOINTER_REG_0__SCAN_IN & P3_INSTADDRPOINTER_REG_1__SCAN_IN & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_553_U5 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P3_ADD_553_U6 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_553_U7 = ~(P3_INSTADDRPOINTER_REG_0__SCAN_IN & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_553_U8 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_553_U10 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_553_U12 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_553_U14 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_553_U16 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_553_U18 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_553_U20 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_553_U21 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_553_U24 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_553_U26 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_553_U28 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_553_U30 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_553_U32 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_553_U34 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_553_U36 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_553_U38 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_553_U40 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_553_U42 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_553_U44 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_553_U46 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_553_U48 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_553_U50 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_553_U52 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_553_U54 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_553_U56 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_553_U58 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_553_U60 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_553_U62 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_553_U64 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_553_U96 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_ADD_558_U5 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P3_ADD_558_U6 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_558_U7 = ~(P3_INSTADDRPOINTER_REG_0__SCAN_IN & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_558_U8 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_558_U10 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_558_U12 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_558_U14 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_558_U16 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_558_U18 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_558_U20 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_558_U21 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_558_U24 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_558_U26 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_558_U28 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_558_U30 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_558_U32 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_558_U34 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_558_U36 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_558_U38 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_558_U40 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_558_U42 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_558_U44 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_558_U46 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_558_U48 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_558_U50 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_558_U52 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_558_U54 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_558_U56 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_558_U58 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_558_U60 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_558_U62 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_558_U64 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_558_U96 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_ADD_385_U5 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P3_ADD_385_U6 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_385_U7 = ~(P3_INSTADDRPOINTER_REG_0__SCAN_IN & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_385_U8 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_385_U10 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_385_U12 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_385_U14 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_385_U16 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_385_U18 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_385_U20 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_385_U21 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_385_U24 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_385_U26 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_385_U28 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_385_U30 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_385_U32 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_385_U34 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_385_U36 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_385_U38 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_385_U40 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_385_U42 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_385_U44 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_385_U46 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_385_U48 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_385_U50 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_385_U52 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_385_U54 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_385_U56 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_385_U58 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_385_U60 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_385_U62 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_385_U64 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_385_U96 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_ADD_547_U5 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P3_ADD_547_U6 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_547_U7 = ~(P3_INSTADDRPOINTER_REG_0__SCAN_IN & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_547_U8 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_547_U10 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_547_U12 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_547_U14 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_547_U16 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_547_U18 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_547_U20 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_547_U21 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_547_U24 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_547_U26 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_547_U28 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_547_U30 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_547_U32 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_547_U34 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_547_U36 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_547_U38 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_547_U40 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_547_U42 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_547_U44 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_547_U46 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_547_U48 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_547_U50 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_547_U52 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_547_U54 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_547_U56 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_547_U58 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_547_U60 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_547_U62 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_547_U64 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_547_U96 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_SUB_412_U8 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign P3_SUB_412_U9 = ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P3_SUB_412_U10 = ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P3_SUB_412_U11 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P3_SUB_412_U12 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign P3_SUB_412_U13 = ~P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign P3_SUB_412_U15 = ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P3_SUB_412_U26 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P3_SUB_412_U27 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN; 
assign P3_ADD_371_1212_U22 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_371_1212_U23 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_371_1212_U27 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_371_1212_U28 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_371_1212_U32 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P3_ADD_371_1212_U33 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_371_1212_U37 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_371_1212_U38 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_371_1212_U41 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_371_1212_U42 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_371_1212_U45 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_371_1212_U46 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_371_1212_U47 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_371_1212_U50 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_371_1212_U51 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_371_1212_U52 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_371_1212_U54 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_371_1212_U55 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_371_1212_U57 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_371_1212_U58 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_371_1212_U60 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_371_1212_U61 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_371_1212_U63 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_371_1212_U64 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_371_1212_U66 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_371_1212_U67 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_371_1212_U69 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_371_1212_U71 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_371_1212_U72 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_371_1212_U74 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_371_1212_U76 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_371_1212_U99 = P3_INSTADDRPOINTER_REG_9__SCAN_IN & P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_371_1212_U100 = P3_INSTADDRPOINTER_REG_11__SCAN_IN & P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_371_1212_U101 = P3_INSTADDRPOINTER_REG_13__SCAN_IN & P3_INSTADDRPOINTER_REG_14__SCAN_IN & P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_371_1212_U102 = P3_INSTADDRPOINTER_REG_16__SCAN_IN & P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_371_1212_U103 = P3_INSTADDRPOINTER_REG_18__SCAN_IN & P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_371_1212_U104 = P3_INSTADDRPOINTER_REG_20__SCAN_IN & P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_371_1212_U105 = P3_INSTADDRPOINTER_REG_22__SCAN_IN & P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_371_1212_U106 = P3_INSTADDRPOINTER_REG_24__SCAN_IN & P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_371_1212_U107 = P3_INSTADDRPOINTER_REG_27__SCAN_IN & P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_371_1212_U116 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_SUB_504_U8 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign P3_SUB_504_U9 = ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P3_SUB_504_U10 = ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P3_SUB_504_U11 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P3_SUB_504_U12 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign P3_SUB_504_U13 = ~P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign P3_SUB_504_U15 = ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P3_SUB_504_U26 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P3_SUB_504_U27 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN; 
assign P3_SUB_401_U8 = ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P3_SUB_401_U10 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign P3_SUB_401_U11 = ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P3_SUB_401_U12 = ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P3_SUB_401_U13 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P3_SUB_401_U14 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign P3_SUB_401_U15 = ~P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign P3_SUB_401_U17 = ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P3_SUB_401_U18 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN; 
assign P3_SUB_401_U29 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P3_SUB_390_U8 = ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P3_SUB_390_U10 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign P3_SUB_390_U11 = ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P3_SUB_390_U12 = ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P3_SUB_390_U13 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P3_SUB_390_U14 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign P3_SUB_390_U15 = ~P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign P3_SUB_390_U17 = ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P3_SUB_390_U18 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN; 
assign P3_SUB_390_U29 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P3_ADD_495_U4 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P3_ADD_495_U5 = ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P3_ADD_495_U6 = ~(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P3_ADD_495_U7 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P3_ADD_495_U11 = ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P3_ADD_494_U4 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_494_U5 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_494_U6 = ~(P3_INSTADDRPOINTER_REG_1__SCAN_IN & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_494_U7 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_494_U9 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_494_U11 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_494_U13 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_494_U15 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_494_U17 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_494_U18 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_494_U21 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_494_U23 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_494_U25 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_494_U27 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_494_U29 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_494_U31 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_494_U33 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_494_U35 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_494_U37 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_494_U39 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_494_U41 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_494_U43 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_494_U45 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_494_U47 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_494_U49 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_494_U51 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_494_U53 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_494_U55 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_494_U57 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_494_U59 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_494_U61 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_494_U92 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_ADD_536_U4 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P3_ADD_536_U5 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_536_U6 = ~(P3_INSTADDRPOINTER_REG_1__SCAN_IN & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_536_U7 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_536_U9 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_536_U11 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_536_U13 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_536_U15 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_ADD_536_U17 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_536_U18 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_ADD_536_U21 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_ADD_536_U23 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_ADD_536_U25 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_ADD_536_U27 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P3_ADD_536_U29 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_ADD_536_U31 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_ADD_536_U33 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P3_ADD_536_U35 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P3_ADD_536_U37 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_ADD_536_U39 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_ADD_536_U41 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P3_ADD_536_U43 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P3_ADD_536_U45 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_ADD_536_U47 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_ADD_536_U49 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_ADD_536_U51 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_ADD_536_U53 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P3_ADD_536_U55 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P3_ADD_536_U57 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P3_ADD_536_U59 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P3_ADD_536_U61 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P3_ADD_536_U92 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P2_R2167_U17 = ~P2_STATE2_REG_0__SCAN_IN; 
assign P2_R2027_U5 = ~P2_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P2_R2027_U6 = ~P2_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P2_R2027_U7 = ~(P2_INSTADDRPOINTER_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P2_R2027_U8 = ~P2_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P2_R2027_U10 = ~P2_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P2_R2027_U12 = ~P2_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P2_R2027_U14 = ~P2_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P2_R2027_U16 = ~P2_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P2_R2027_U18 = ~P2_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P2_R2027_U20 = ~P2_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P2_R2027_U21 = ~P2_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P2_R2027_U24 = ~P2_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P2_R2027_U26 = ~P2_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P2_R2027_U28 = ~P2_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P2_R2027_U30 = ~P2_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P2_R2027_U32 = ~P2_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P2_R2027_U34 = ~P2_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P2_R2027_U36 = ~P2_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P2_R2027_U38 = ~P2_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P2_R2027_U40 = ~P2_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P2_R2027_U42 = ~P2_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P2_R2027_U44 = ~P2_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P2_R2027_U46 = ~P2_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P2_R2027_U48 = ~P2_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P2_R2027_U50 = ~P2_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P2_R2027_U52 = ~P2_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P2_R2027_U54 = ~P2_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P2_R2027_U56 = ~P2_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P2_R2027_U58 = ~P2_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P2_R2027_U60 = ~P2_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P2_R2027_U62 = ~P2_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P2_R2027_U64 = ~P2_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P2_R2027_U96 = ~P2_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P2_R2337_U4 = ~P2_PHYADDRPOINTER_REG_1__SCAN_IN; 
assign P2_R2337_U5 = ~P2_PHYADDRPOINTER_REG_3__SCAN_IN; 
assign P2_R2337_U6 = ~P2_PHYADDRPOINTER_REG_2__SCAN_IN; 
assign P2_R2337_U7 = ~(P2_PHYADDRPOINTER_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_2__SCAN_IN & P2_PHYADDRPOINTER_REG_3__SCAN_IN); 
assign P2_R2337_U8 = ~P2_PHYADDRPOINTER_REG_4__SCAN_IN; 
assign P2_R2337_U10 = ~P2_PHYADDRPOINTER_REG_5__SCAN_IN; 
assign P2_R2337_U12 = ~P2_PHYADDRPOINTER_REG_6__SCAN_IN; 
assign P2_R2337_U14 = ~P2_PHYADDRPOINTER_REG_7__SCAN_IN; 
assign P2_R2337_U16 = ~P2_PHYADDRPOINTER_REG_8__SCAN_IN; 
assign P2_R2337_U17 = ~P2_PHYADDRPOINTER_REG_9__SCAN_IN; 
assign P2_R2337_U20 = ~P2_PHYADDRPOINTER_REG_10__SCAN_IN; 
assign P2_R2337_U22 = ~P2_PHYADDRPOINTER_REG_11__SCAN_IN; 
assign P2_R2337_U24 = ~P2_PHYADDRPOINTER_REG_12__SCAN_IN; 
assign P2_R2337_U26 = ~P2_PHYADDRPOINTER_REG_13__SCAN_IN; 
assign P2_R2337_U28 = ~P2_PHYADDRPOINTER_REG_14__SCAN_IN; 
assign P2_R2337_U30 = ~P2_PHYADDRPOINTER_REG_15__SCAN_IN; 
assign P2_R2337_U32 = ~P2_PHYADDRPOINTER_REG_16__SCAN_IN; 
assign P2_R2337_U34 = ~P2_PHYADDRPOINTER_REG_17__SCAN_IN; 
assign P2_R2337_U36 = ~P2_PHYADDRPOINTER_REG_18__SCAN_IN; 
assign P2_R2337_U38 = ~P2_PHYADDRPOINTER_REG_19__SCAN_IN; 
assign P2_R2337_U40 = ~P2_PHYADDRPOINTER_REG_20__SCAN_IN; 
assign P2_R2337_U42 = ~P2_PHYADDRPOINTER_REG_21__SCAN_IN; 
assign P2_R2337_U44 = ~P2_PHYADDRPOINTER_REG_22__SCAN_IN; 
assign P2_R2337_U46 = ~P2_PHYADDRPOINTER_REG_23__SCAN_IN; 
assign P2_R2337_U48 = ~P2_PHYADDRPOINTER_REG_24__SCAN_IN; 
assign P2_R2337_U50 = ~P2_PHYADDRPOINTER_REG_25__SCAN_IN; 
assign P2_R2337_U52 = ~P2_PHYADDRPOINTER_REG_26__SCAN_IN; 
assign P2_R2337_U54 = ~P2_PHYADDRPOINTER_REG_27__SCAN_IN; 
assign P2_R2337_U56 = ~P2_PHYADDRPOINTER_REG_28__SCAN_IN; 
assign P2_R2337_U58 = ~P2_PHYADDRPOINTER_REG_29__SCAN_IN; 
assign P2_R2337_U60 = ~P2_PHYADDRPOINTER_REG_30__SCAN_IN; 
assign P2_R2337_U91 = ~(P2_PHYADDRPOINTER_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_2__SCAN_IN); 
assign P2_R2337_U92 = ~P2_PHYADDRPOINTER_REG_31__SCAN_IN; 
assign P2_R2147_U4 = ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P2_R2147_U5 = ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_R2147_U6 = ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P2_R2147_U11 = ~(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P2_R2147_U12 = ~(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P2_LT_563_U8 = ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign P2_LT_563_U9 = ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P2_LT_563_U12 = ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign P2_LT_563_U13 = ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign P2_R2238_U8 = ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P2_R2238_U10 = ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign P2_R2238_U11 = ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P2_R2238_U12 = ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P2_R2238_U13 = ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_R2238_U14 = ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign P2_R2238_U15 = ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign P2_R2238_U17 = ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P2_R2238_U18 = ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN; 
assign P2_R2238_U29 = ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P2_R2278_U8 = ~P2_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P2_R2278_U10 = ~P2_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P2_R2278_U12 = ~P2_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P2_R2278_U14 = ~P2_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P2_R2278_U17 = ~P2_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P2_R2278_U19 = ~P2_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P2_R2278_U22 = ~P2_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P2_R2278_U25 = ~P2_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P2_R2278_U28 = ~P2_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P2_R2278_U29 = ~P2_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P2_R2278_U32 = ~P2_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P2_R2278_U34 = ~P2_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P2_R2278_U36 = ~P2_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P2_R2278_U38 = ~P2_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P2_R2278_U40 = ~P2_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P2_R2278_U42 = ~P2_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P2_R2278_U44 = ~P2_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P2_R2278_U46 = ~P2_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P2_R2278_U48 = ~P2_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P2_R2278_U51 = ~P2_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P2_R2278_U54 = ~P2_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P2_R2278_U57 = ~P2_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P2_R2278_U60 = ~P2_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P2_R2278_U63 = ~P2_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P2_R2278_U65 = ~P2_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P2_R2278_U67 = ~P2_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P2_R2278_U70 = ~P2_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P2_R2278_U73 = ~P2_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P2_R2278_U75 = ~P2_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P2_R2278_U77 = ~P2_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P2_R2278_U80 = ~P2_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P2_R2278_U159 = ~P2_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P2_SUB_450_U8 = ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign P2_SUB_450_U9 = ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P2_SUB_450_U10 = ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P2_SUB_450_U11 = ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_SUB_450_U12 = ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign P2_SUB_450_U13 = ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign P2_SUB_450_U15 = ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P2_SUB_450_U16 = ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN; 
assign P2_SUB_450_U27 = ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P2_ADD_394_U4 = ~P2_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P2_ADD_394_U6 = ~P2_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P2_ADD_394_U7 = ~P2_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P2_ADD_394_U9 = ~P2_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P2_ADD_394_U11 = ~P2_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P2_ADD_394_U12 = ~P2_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P2_ADD_394_U15 = ~P2_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P2_ADD_394_U17 = ~P2_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P2_ADD_394_U19 = ~P2_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P2_ADD_394_U21 = ~P2_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P2_ADD_394_U23 = ~P2_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P2_ADD_394_U25 = ~P2_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P2_ADD_394_U27 = ~P2_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P2_ADD_394_U29 = ~P2_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P2_ADD_394_U31 = ~P2_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P2_ADD_394_U33 = ~P2_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P2_ADD_394_U35 = ~P2_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P2_ADD_394_U37 = ~P2_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P2_ADD_394_U39 = ~P2_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P2_ADD_394_U41 = ~P2_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P2_ADD_394_U43 = ~P2_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P2_ADD_394_U45 = ~P2_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P2_ADD_394_U47 = ~P2_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P2_ADD_394_U49 = ~P2_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P2_ADD_394_U51 = ~P2_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P2_ADD_394_U53 = ~P2_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P2_ADD_394_U55 = ~P2_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P2_ADD_394_U57 = ~P2_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P2_ADD_394_U59 = ~P2_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P2_ADD_394_U60 = ~P2_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P2_ADD_394_U62 = ~P2_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P2_ADD_394_U92 = ~P2_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P2_ADD_394_U96 = ~(P2_INSTADDRPOINTER_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P2_ADD_394_U125 = ~(P2_INSTADDRPOINTER_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_1__SCAN_IN & P2_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P2_ADD_371_1212_U5 = P2_INSTADDRPOINTER_REG_9__SCAN_IN & P2_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P2_ADD_371_1212_U10 = P2_INSTADDRPOINTER_REG_9__SCAN_IN & P2_INSTADDRPOINTER_REG_10__SCAN_IN & P2_INSTADDRPOINTER_REG_11__SCAN_IN & P2_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P2_ADD_371_1212_U26 = ~P2_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P2_ADD_371_1212_U28 = ~P2_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P2_ADD_371_1212_U32 = ~P2_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P2_ADD_371_1212_U34 = ~P2_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P2_ADD_371_1212_U36 = ~P2_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P2_ADD_371_1212_U38 = ~P2_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P2_ADD_371_1212_U39 = ~P2_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P2_ADD_371_1212_U42 = ~P2_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P2_ADD_371_1212_U44 = ~P2_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P2_ADD_371_1212_U45 = ~P2_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P2_ADD_371_1212_U46 = ~P2_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P2_ADD_371_1212_U47 = ~P2_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P2_ADD_371_1212_U48 = ~P2_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P2_ADD_371_1212_U49 = ~P2_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P2_ADD_371_1212_U50 = ~P2_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P2_ADD_371_1212_U51 = ~P2_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P2_ADD_371_1212_U52 = ~P2_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P2_ADD_371_1212_U53 = ~P2_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P2_ADD_371_1212_U54 = ~P2_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P2_ADD_371_1212_U55 = ~P2_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P2_ADD_371_1212_U56 = ~P2_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P2_ADD_371_1212_U57 = ~P2_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P2_ADD_371_1212_U58 = ~P2_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P2_ADD_371_1212_U59 = ~P2_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P2_ADD_371_1212_U60 = ~P2_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P2_ADD_371_1212_U61 = ~P2_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P2_ADD_371_1212_U62 = ~P2_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P2_ADD_371_1212_U63 = ~P2_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P2_ADD_371_1212_U64 = ~P2_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P2_ADD_371_1212_U65 = ~P2_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P2_ADD_371_1212_U66 = ~P2_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P2_ADD_371_1212_U87 = P2_INSTADDRPOINTER_REG_13__SCAN_IN & P2_INSTADDRPOINTER_REG_14__SCAN_IN & P2_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P2_ADD_371_1212_U88 = P2_INSTADDRPOINTER_REG_16__SCAN_IN & P2_INSTADDRPOINTER_REG_17__SCAN_IN & P2_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P2_ADD_371_1212_U89 = P2_INSTADDRPOINTER_REG_19__SCAN_IN & P2_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P2_ADD_371_1212_U90 = P2_INSTADDRPOINTER_REG_21__SCAN_IN & P2_INSTADDRPOINTER_REG_22__SCAN_IN & P2_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P2_ADD_371_1212_U91 = P2_INSTADDRPOINTER_REG_24__SCAN_IN & P2_INSTADDRPOINTER_REG_25__SCAN_IN & P2_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P2_ADD_371_1212_U92 = P2_INSTADDRPOINTER_REG_27__SCAN_IN & P2_INSTADDRPOINTER_REG_28__SCAN_IN & P2_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P2_ADD_371_1212_U94 = P2_INSTADDRPOINTER_REG_27__SCAN_IN & P2_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P2_ADD_371_1212_U98 = P2_INSTADDRPOINTER_REG_21__SCAN_IN & P2_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P2_ADD_371_1212_U101 = P2_INSTADDRPOINTER_REG_16__SCAN_IN & P2_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P2_ADD_371_1212_U104 = P2_INSTADDRPOINTER_REG_24__SCAN_IN & P2_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P2_ADD_371_1212_U128 = ~P2_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P1_R2027_U5 = ~P1_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P1_R2027_U6 = ~P1_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P1_R2027_U7 = ~P1_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P1_R2027_U8 = ~P1_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P1_R2027_U9 = ~P1_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P1_R2027_U10 = ~(P1_INSTADDRPOINTER_REG_0__SCAN_IN & P1_INSTADDRPOINTER_REG_1__SCAN_IN & P1_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P1_R2027_U11 = ~P1_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P1_R2027_U12 = ~P1_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P1_R2027_U14 = ~P1_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P1_R2027_U15 = ~P1_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P1_R2027_U18 = ~P1_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P1_R2027_U19 = ~P1_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P1_R2027_U20 = ~P1_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P1_R2027_U21 = ~P1_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P1_R2027_U23 = ~P1_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P1_R2027_U24 = ~P1_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P1_R2027_U26 = ~P1_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P1_R2027_U28 = ~P1_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P1_R2027_U29 = ~P1_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P1_R2027_U30 = ~P1_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P1_R2027_U32 = ~P1_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P1_R2027_U33 = ~P1_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P1_R2027_U35 = ~P1_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P1_R2027_U37 = ~P1_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P1_R2027_U38 = ~P1_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P1_R2027_U39 = ~P1_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P1_R2027_U41 = ~P1_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P1_R2027_U42 = ~P1_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P1_R2027_U44 = ~P1_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P1_R2027_U45 = ~P1_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P1_R2027_U47 = ~P1_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P1_R2027_U50 = ~P1_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P1_R2027_U82 = P1_INSTADDRPOINTER_REG_3__SCAN_IN & P1_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P1_R2027_U83 = P1_INSTADDRPOINTER_REG_5__SCAN_IN & P1_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P1_R2027_U84 = P1_INSTADDRPOINTER_REG_7__SCAN_IN & P1_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P1_R2027_U85 = P1_INSTADDRPOINTER_REG_9__SCAN_IN & P1_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P1_R2027_U86 = P1_INSTADDRPOINTER_REG_11__SCAN_IN & P1_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P1_R2027_U87 = P1_INSTADDRPOINTER_REG_13__SCAN_IN & P1_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P1_R2027_U88 = P1_INSTADDRPOINTER_REG_15__SCAN_IN & P1_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P1_R2027_U89 = P1_INSTADDRPOINTER_REG_17__SCAN_IN & P1_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P1_R2027_U90 = P1_INSTADDRPOINTER_REG_19__SCAN_IN & P1_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P1_R2027_U91 = P1_INSTADDRPOINTER_REG_21__SCAN_IN & P1_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P1_R2027_U92 = P1_INSTADDRPOINTER_REG_23__SCAN_IN & P1_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P1_R2027_U93 = P1_INSTADDRPOINTER_REG_25__SCAN_IN & P1_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P1_R2027_U94 = P1_INSTADDRPOINTER_REG_27__SCAN_IN & P1_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P1_R2027_U98 = ~P1_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P1_R2027_U100 = ~(P1_INSTADDRPOINTER_REG_0__SCAN_IN & P1_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P1_R2278_U21 = ~P1_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P1_R2278_U23 = ~P1_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P1_R2278_U25 = ~P1_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P1_R2278_U27 = ~P1_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P1_R2278_U30 = ~P1_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P1_R2278_U31 = ~P1_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P1_R2278_U34 = ~P1_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P1_R2278_U36 = ~P1_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P1_R2278_U38 = ~P1_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P1_R2278_U44 = ~P1_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P1_R2278_U46 = ~P1_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P1_R2278_U48 = ~P1_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P1_R2278_U50 = ~P1_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P1_R2278_U52 = ~P1_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P1_R2278_U54 = ~P1_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P1_R2278_U56 = ~P1_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P1_R2278_U58 = ~P1_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P1_R2278_U60 = ~P1_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P1_R2278_U62 = ~P1_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P1_R2278_U64 = ~P1_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P1_R2278_U66 = ~P1_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P1_R2278_U69 = ~P1_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P1_R2278_U71 = ~P1_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P1_R2278_U74 = ~P1_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P1_R2278_U77 = ~P1_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P1_R2278_U82 = ~P1_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P1_R2278_U83 = ~P1_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P1_R2278_U89 = ~P1_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P1_R2278_U91 = ~P1_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P1_R2278_U185 = ~P1_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P1_R2167_U16 = ~P1_STATE2_REG_0__SCAN_IN; 
assign P1_R2337_U4 = ~P1_PHYADDRPOINTER_REG_1__SCAN_IN; 
assign P1_R2337_U5 = ~P1_PHYADDRPOINTER_REG_2__SCAN_IN; 
assign P1_R2337_U6 = ~(P1_PHYADDRPOINTER_REG_1__SCAN_IN & P1_PHYADDRPOINTER_REG_2__SCAN_IN); 
assign P1_R2337_U7 = ~P1_PHYADDRPOINTER_REG_3__SCAN_IN; 
assign P1_R2337_U9 = ~P1_PHYADDRPOINTER_REG_4__SCAN_IN; 
assign P1_R2337_U11 = ~P1_PHYADDRPOINTER_REG_5__SCAN_IN; 
assign P1_R2337_U13 = ~P1_PHYADDRPOINTER_REG_6__SCAN_IN; 
assign P1_R2337_U15 = ~P1_PHYADDRPOINTER_REG_7__SCAN_IN; 
assign P1_R2337_U17 = ~P1_PHYADDRPOINTER_REG_8__SCAN_IN; 
assign P1_R2337_U18 = ~P1_PHYADDRPOINTER_REG_9__SCAN_IN; 
assign P1_R2337_U21 = ~P1_PHYADDRPOINTER_REG_10__SCAN_IN; 
assign P1_R2337_U23 = ~P1_PHYADDRPOINTER_REG_11__SCAN_IN; 
assign P1_R2337_U25 = ~P1_PHYADDRPOINTER_REG_12__SCAN_IN; 
assign P1_R2337_U27 = ~P1_PHYADDRPOINTER_REG_13__SCAN_IN; 
assign P1_R2337_U29 = ~P1_PHYADDRPOINTER_REG_14__SCAN_IN; 
assign P1_R2337_U31 = ~P1_PHYADDRPOINTER_REG_15__SCAN_IN; 
assign P1_R2337_U33 = ~P1_PHYADDRPOINTER_REG_16__SCAN_IN; 
assign P1_R2337_U35 = ~P1_PHYADDRPOINTER_REG_17__SCAN_IN; 
assign P1_R2337_U37 = ~P1_PHYADDRPOINTER_REG_18__SCAN_IN; 
assign P1_R2337_U39 = ~P1_PHYADDRPOINTER_REG_19__SCAN_IN; 
assign P1_R2337_U41 = ~P1_PHYADDRPOINTER_REG_20__SCAN_IN; 
assign P1_R2337_U43 = ~P1_PHYADDRPOINTER_REG_21__SCAN_IN; 
assign P1_R2337_U45 = ~P1_PHYADDRPOINTER_REG_22__SCAN_IN; 
assign P1_R2337_U47 = ~P1_PHYADDRPOINTER_REG_23__SCAN_IN; 
assign P1_R2337_U49 = ~P1_PHYADDRPOINTER_REG_24__SCAN_IN; 
assign P1_R2337_U51 = ~P1_PHYADDRPOINTER_REG_25__SCAN_IN; 
assign P1_R2337_U53 = ~P1_PHYADDRPOINTER_REG_26__SCAN_IN; 
assign P1_R2337_U55 = ~P1_PHYADDRPOINTER_REG_27__SCAN_IN; 
assign P1_R2337_U57 = ~P1_PHYADDRPOINTER_REG_28__SCAN_IN; 
assign P1_R2337_U59 = ~P1_PHYADDRPOINTER_REG_29__SCAN_IN; 
assign P1_R2337_U61 = ~P1_PHYADDRPOINTER_REG_30__SCAN_IN; 
assign P1_R2337_U92 = ~P1_PHYADDRPOINTER_REG_31__SCAN_IN; 
assign P1_SUB_580_U7 = ~P1_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P1_SUB_580_U8 = ~P1_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P1_R2096_U4 = ~P1_REIP_REG_1__SCAN_IN; 
assign P1_R2096_U5 = ~P1_REIP_REG_2__SCAN_IN; 
assign P1_R2096_U6 = ~(P1_REIP_REG_1__SCAN_IN & P1_REIP_REG_2__SCAN_IN); 
assign P1_R2096_U7 = ~P1_REIP_REG_3__SCAN_IN; 
assign P1_R2096_U9 = ~P1_REIP_REG_4__SCAN_IN; 
assign P1_R2096_U11 = ~P1_REIP_REG_5__SCAN_IN; 
assign P1_R2096_U13 = ~P1_REIP_REG_6__SCAN_IN; 
assign P1_R2096_U15 = ~P1_REIP_REG_7__SCAN_IN; 
assign P1_R2096_U17 = ~P1_REIP_REG_8__SCAN_IN; 
assign P1_R2096_U18 = ~P1_REIP_REG_9__SCAN_IN; 
assign P1_R2096_U21 = ~P1_REIP_REG_10__SCAN_IN; 
assign P1_R2096_U23 = ~P1_REIP_REG_11__SCAN_IN; 
assign P1_R2096_U25 = ~P1_REIP_REG_12__SCAN_IN; 
assign P1_R2096_U27 = ~P1_REIP_REG_13__SCAN_IN; 
assign P1_R2096_U29 = ~P1_REIP_REG_14__SCAN_IN; 
assign P1_R2096_U31 = ~P1_REIP_REG_15__SCAN_IN; 
assign P1_R2096_U33 = ~P1_REIP_REG_16__SCAN_IN; 
assign P1_R2096_U35 = ~P1_REIP_REG_17__SCAN_IN; 
assign P1_R2096_U37 = ~P1_REIP_REG_18__SCAN_IN; 
assign P1_R2096_U39 = ~P1_REIP_REG_19__SCAN_IN; 
assign P1_R2096_U41 = ~P1_REIP_REG_20__SCAN_IN; 
assign P1_R2096_U43 = ~P1_REIP_REG_21__SCAN_IN; 
assign P1_R2096_U45 = ~P1_REIP_REG_22__SCAN_IN; 
assign P1_R2096_U47 = ~P1_REIP_REG_23__SCAN_IN; 
assign P1_R2096_U49 = ~P1_REIP_REG_24__SCAN_IN; 
assign P1_R2096_U51 = ~P1_REIP_REG_25__SCAN_IN; 
assign P1_R2096_U53 = ~P1_REIP_REG_26__SCAN_IN; 
assign P1_R2096_U55 = ~P1_REIP_REG_27__SCAN_IN; 
assign P1_R2096_U57 = ~P1_REIP_REG_28__SCAN_IN; 
assign P1_R2096_U59 = ~P1_REIP_REG_29__SCAN_IN; 
assign P1_R2096_U61 = ~P1_REIP_REG_30__SCAN_IN; 
assign P1_R2096_U92 = ~P1_REIP_REG_31__SCAN_IN; 
assign P1_LT_563_U7 = ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P1_LT_563_U10 = ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign P1_LT_563_U11 = ~P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign P1_R2238_U8 = ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_R2238_U10 = ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign P1_R2238_U11 = ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P1_R2238_U12 = ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P1_R2238_U13 = ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P1_R2238_U14 = ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign P1_R2238_U15 = ~P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign P1_R2238_U17 = ~P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P1_R2238_U18 = ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN; 
assign P1_R2238_U29 = ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P1_SUB_450_U8 = ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_SUB_450_U10 = ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign P1_SUB_450_U11 = ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P1_SUB_450_U12 = ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P1_SUB_450_U13 = ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P1_SUB_450_U14 = ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign P1_SUB_450_U15 = ~P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign P1_SUB_450_U17 = ~P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P1_SUB_450_U18 = ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN; 
assign P1_SUB_450_U29 = ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P1_ADD_405_U4 = ~P1_INSTADDRPOINTER_REG_0__SCAN_IN; 
assign P1_ADD_405_U6 = ~P1_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P1_ADD_405_U7 = ~P1_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P1_ADD_405_U9 = ~P1_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P1_ADD_405_U11 = ~P1_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P1_ADD_405_U12 = ~P1_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P1_ADD_405_U15 = ~P1_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P1_ADD_405_U17 = ~P1_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P1_ADD_405_U19 = ~P1_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P1_ADD_405_U21 = ~P1_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P1_ADD_405_U23 = ~P1_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P1_ADD_405_U25 = ~P1_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P1_ADD_405_U27 = ~P1_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P1_ADD_405_U29 = ~P1_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P1_ADD_405_U31 = ~P1_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P1_ADD_405_U33 = ~P1_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P1_ADD_405_U35 = ~P1_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P1_ADD_405_U37 = ~P1_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P1_ADD_405_U39 = ~P1_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P1_ADD_405_U41 = ~P1_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P1_ADD_405_U43 = ~P1_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P1_ADD_405_U45 = ~P1_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P1_ADD_405_U47 = ~P1_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P1_ADD_405_U49 = ~P1_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P1_ADD_405_U51 = ~P1_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P1_ADD_405_U53 = ~P1_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P1_ADD_405_U55 = ~P1_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P1_ADD_405_U57 = ~P1_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P1_ADD_405_U59 = ~P1_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P1_ADD_405_U60 = ~P1_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P1_ADD_405_U62 = ~P1_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P1_ADD_405_U92 = ~P1_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P1_ADD_405_U96 = ~(P1_INSTADDRPOINTER_REG_0__SCAN_IN & P1_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P1_ADD_405_U125 = ~(P1_INSTADDRPOINTER_REG_0__SCAN_IN & P1_INSTADDRPOINTER_REG_1__SCAN_IN & P1_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P1_ADD_515_U4 = ~P1_INSTADDRPOINTER_REG_1__SCAN_IN; 
assign P1_ADD_515_U5 = ~P1_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P1_ADD_515_U6 = ~(P1_INSTADDRPOINTER_REG_1__SCAN_IN & P1_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P1_ADD_515_U7 = ~P1_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P1_ADD_515_U9 = ~P1_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P1_ADD_515_U11 = ~P1_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P1_ADD_515_U12 = ~P1_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P1_ADD_515_U15 = ~P1_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P1_ADD_515_U17 = ~P1_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P1_ADD_515_U19 = ~P1_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P1_ADD_515_U21 = ~P1_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P1_ADD_515_U23 = ~P1_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P1_ADD_515_U25 = ~P1_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P1_ADD_515_U27 = ~P1_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P1_ADD_515_U29 = ~P1_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P1_ADD_515_U31 = ~P1_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P1_ADD_515_U33 = ~P1_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P1_ADD_515_U35 = ~P1_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P1_ADD_515_U37 = ~P1_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P1_ADD_515_U39 = ~P1_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P1_ADD_515_U41 = ~P1_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P1_ADD_515_U43 = ~P1_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P1_ADD_515_U45 = ~P1_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P1_ADD_515_U47 = ~P1_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P1_ADD_515_U49 = ~P1_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P1_ADD_515_U51 = ~P1_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P1_ADD_515_U53 = ~P1_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P1_ADD_515_U55 = ~P1_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P1_ADD_515_U57 = ~P1_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P1_ADD_515_U59 = ~P1_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P1_ADD_515_U60 = ~P1_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P1_ADD_515_U92 = ~P1_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign U208 = U378 & U377 & P2_W_R_N_REG_SCAN_IN & P2_M_IO_N_REG_SCAN_IN; 
assign P3_U2352 = ~(U209 | P3_STATEBS16_REG_SCAN_IN); 
assign P3_U2466 = P3_U3093 & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P3_U2468 = P3_U3094 & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P3_U2492 = P3_U3128 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P3_U2629 = P3_U3207 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P3_U2630 = ~U209; 
assign P3_U2632 = P3_U3207 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P3_U3077 = ~(P3_U3085 & P3_STATE_REG_1__SCAN_IN); 
assign P3_U3082 = ~(P3_U3079 & P3_STATE_REG_1__SCAN_IN); 
assign P3_U3087 = ~(P3_U3084 & P3_REQUESTPENDING_REG_SCAN_IN); 
assign P3_U3098 = ~(P3_U3100 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_U3124 = ~(P3_U3089 & P3_STATE2_REG_2__SCAN_IN); 
assign P3_U3126 = ~(P3_LTE_597_U6 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U3153 = ~(P3_U3129 & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P3_U3169 = ~(P3_U3457 & P3_U2501); 
assign P3_U3177 = ~(P3_U3129 & P3_U2501 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_U3199 = ~(P3_U3133 & P3_U2501 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_U3205 = ~(P3_U3634 & P3_U2501); 
assign P3_U3223 = ~(P3_U5503 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_U3227 = ~(P3_U3095 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_U3228 = ~(P3_U3091 & P3_U3095); 
assign P3_U3234 = ~(P3_U3135 & P3_U3123); 
assign P3_U3257 = U209 | P3_STATEBS16_REG_SCAN_IN; 
assign P3_U3279 = P3_U3083 & P3_U4286; 
assign P3_U3422 = P3_U3129 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign P3_U3475 = P3_U3131 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign P3_U3527 = P3_U3133 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign P3_U3545 = P3_U3133 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P3_U3670 = P3_U3093 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P3_U3952 = P3_U3121 & P3_STATE2_REG_2__SCAN_IN; 
assign P3_U4138 = P3_U4137 & P3_U4136; 
assign P3_U4141 = P3_U4140 & P3_U4139; 
assign P3_U4144 = P3_U4143 & P3_U4142; 
assign P3_U4148 = P3_U4147 & P3_U7366 & P3_U4146 & P3_U4145; 
assign P3_U4289 = ~(P3_U3091 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_U4295 = ~P3_U3135; 
assign P3_U4329 = ~(P3_U3121 & P3_U3090 & P3_U2631 & P3_STATE2_REG_1__SCAN_IN); 
assign P3_U4330 = ~(P3_U3653 & P3_U2453); 
assign P3_U4332 = ~P3_U3095; 
assign P3_U4338 = ~(P3_U3090 & U209 & P3_STATE2_REG_0__SCAN_IN); 
assign P3_U4340 = ~P3_U3123; 
assign P3_U4354 = ~P3_U3125; 
assign P3_U4448 = ~P3_U3088; 
assign P3_U4452 = ~P3_U3083; 
assign P3_U4461 = ~(NA & P3_U3085); 
assign P3_U4464 = ~(P3_U4286 & P3_U3083); 
assign P3_U4465 = ~(P3_U3076 & P3_STATE_REG_2__SCAN_IN); 
assign P3_U4467 = ~P3_U3091; 
assign P3_U4628 = ~(U209 & P3_STATE2_REG_1__SCAN_IN); 
assign P3_U4641 = ~(P3_U3128 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_U4648 = ~P3_U3130; 
assign P3_U4665 = ~(P3_U3090 & P3_STATE2_REG_1__SCAN_IN); 
assign P3_U5498 = ~(P3_U3121 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U5500 = ~(P3_U3095 & P3_U3097); 
assign P3_U5502 = ~(P3_U2481 & P3_U3095); 
assign P3_U5596 = ~(P3_U3130 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U5601 = ~(P3_U3129 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U5607 = ~(P3_U3128 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U5613 = ~(P3_U3128 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U6758 = ~(P3_U2453 & P3_U3121); 
assign P3_U7096 = U209 | P3_STATEBS16_REG_SCAN_IN; 
assign P3_U7774 = ~(P3_U3097 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_U7905 = U209 | P3_STATE2_REG_2__SCAN_IN; 
assign P3_U7928 = ~(P3_U3079 & P3_STATE_REG_0__SCAN_IN & P3_REQUESTPENDING_REG_SCAN_IN); 
assign P3_U7960 = ~(P3_U3130 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_U7983 = ~(P3_U4284 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_U7986 = ~(P3_U4284 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_U8005 = ~(P3_U3240 & P3_DATAWIDTH_REG_0__SCAN_IN); 
assign P3_U8032 = ~(P3_U3097 & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P3_U8033 = ~(P3_U3094 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_U8038 = ~(P3_U3207 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_U8040 = ~(P3_U3207 & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P3_U8042 = ~(P3_U3207 & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P2_U2360 = ~(U211 | P2_STATEBS16_REG_SCAN_IN); 
assign P2_U2452 = P2_U3272 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P2_U2453 = P2_U3271 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P2_U2454 = P2_U3271 & P2_U3272 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P2_U2455 = P2_U3276 & P2_U3272 & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P2_U2456 = P2_U3276 & P2_U3271 & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P2_U2465 = P2_U3309 & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P2_U2615 = P2_U3519 & P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P2_U2813 = P2_U3519 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P2_U3259 = ~(P2_U3266 & P2_STATE_REG_1__SCAN_IN); 
assign P2_U3262 = ~(P2_U3244 & P2_STATE_REG_1__SCAN_IN); 
assign P2_U3265 = ~U211; 
assign P2_U3267 = ~(P2_U3264 & P2_REQUESTPENDING_REG_SCAN_IN); 
assign P2_U3274 = ~(P2_U3276 & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P2_U3301 = ~(P2_U3270 & P2_STATE2_REG_0__SCAN_IN); 
assign P2_U3304 = ~(P2_U3269 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U3335 = ~(P2_U3307 & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P2_U3349 = ~(P2_U3308 & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P2_U3365 = ~(P2_U2478 & P2_U2464); 
assign P2_U3376 = ~(P2_U3310 & P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P2_U3508 = ~(P2_U2503 & P2_U2478); 
assign P2_U3531 = ~P2_R2147_U4; 
assign P2_U3540 = ~(P2_U3284 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U3545 = U211 | P2_STATEBS16_REG_SCAN_IN; 
assign P2_U3590 = P2_U3263 & P2_U4401; 
assign P2_U3607 = P2_U4183 & P2_U7898; 
assign P2_U3714 = P2_U3573 & P2_STATE2_REG_2__SCAN_IN; 
assign P2_U3718 = P2_U3269 & P2_STATE2_REG_3__SCAN_IN; 
assign P2_U4171 = P2_U4170 & P2_U4169; 
assign P2_U4174 = P2_U4173 & P2_U4172; 
assign P2_U4177 = P2_U4176 & P2_U4175; 
assign P2_U4181 = P2_U4180 & P2_U6835 & P2_U4179 & P2_U4178; 
assign P2_U4276 = P2_U3300 & P2_STATE2_REG_2__SCAN_IN & P2_STATE2_REG_0__SCAN_IN; 
assign P2_U4405 = ~(P2_U7006 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P2_U4430 = ~P2_U3313; 
assign P2_U4454 = ~(P2_U3302 & P2_U3270 & P2_U3284 & P2_STATE2_REG_1__SCAN_IN); 
assign P2_U4455 = ~(P2_U3867 & P2_U2448); 
assign P2_U4466 = ~P2_U3303; 
assign P2_U4471 = ~P2_U3573; 
assign P2_U4571 = ~P2_U3268; 
assign P2_U4574 = ~P2_U3263; 
assign P2_U4576 = ~(P2_U3268 & U211 & P2_STATE_REG_1__SCAN_IN); 
assign P2_U4586 = ~(NA & P2_U3266); 
assign P2_U4589 = ~(P2_U4401 & P2_U3263); 
assign P2_U4590 = ~P2_U3277; 
assign P2_U4593 = ~P2_U3275; 
assign P2_U4594 = ~(P2_U3258 & P2_STATE_REG_2__SCAN_IN); 
assign P2_U4622 = ~(P2_U3284 & P2_STATEBS16_REG_SCAN_IN); 
assign P2_U4642 = ~P2_U3311; 
assign P2_U4646 = ~(P2_U3311 & P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P2_U4655 = ~(P2_U3270 & P2_STATE2_REG_1__SCAN_IN); 
assign P2_U5583 = ~(P2_U3284 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U5585 = ~(P2_U4591 & P2_U3276); 
assign P2_U5615 = ~(P2_U4591 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P2_U5661 = ~(P2_U3313 & P2_U3303); 
assign P2_U5939 = ~(P2_U3302 & P2_STATE2_REG_1__SCAN_IN); 
assign P2_U6572 = U211 | P2_STATEBS16_REG_SCAN_IN; 
assign P2_U7585 = ~(P2_U3284 & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P2_U7727 = ~(P2_U3284 & P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P2_U7729 = ~(P2_U3284 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7731 = ~(P2_U3284 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P2_U7733 = ~(P2_U3284 & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P2_U7735 = ~(P2_U3284 & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P2_U7892 = ~(P2_U3244 & P2_STATE_REG_0__SCAN_IN & P2_REQUESTPENDING_REG_SCAN_IN); 
assign P2_U7909 = ~(P2_U3266 & P2_STATE_REG_2__SCAN_IN); 
assign P2_U7922 = ~(P2_U3388 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7925 = ~(P2_U3422 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7927 = ~(P2_U3411 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7928 = ~(P2_U3374 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7930 = ~(P2_U3333 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7932 = ~(P2_U3363 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7934 = ~(P2_U3347 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7936 = ~(P2_U3399 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7938 = ~(P2_U3389 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7941 = ~(P2_U3423 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7943 = ~(P2_U3412 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7944 = ~(P2_U3375 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7946 = ~(P2_U3334 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7948 = ~(P2_U3364 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7950 = ~(P2_U3348 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7952 = ~(P2_U3400 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7954 = ~(P2_U3385 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7957 = ~(P2_U3419 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7959 = ~(P2_U3408 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7960 = ~(P2_U3371 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7962 = ~(P2_U3330 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7964 = ~(P2_U3360 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7966 = ~(P2_U3344 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7968 = ~(P2_U3396 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7970 = ~(P2_U3383 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7973 = ~(P2_U3417 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7975 = ~(P2_U3406 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7976 = ~(P2_U3369 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7978 = ~(P2_U3328 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7980 = ~(P2_U3358 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7982 = ~(P2_U3342 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7984 = ~(P2_U3394 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7986 = ~(P2_U3384 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7989 = ~(P2_U3418 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7991 = ~(P2_U3407 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7992 = ~(P2_U3370 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7994 = ~(P2_U3329 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7996 = ~(P2_U3359 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7998 = ~(P2_U3343 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8000 = ~(P2_U3395 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8002 = ~(P2_U3387 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8005 = ~(P2_U3421 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8007 = ~(P2_U3410 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8008 = ~(P2_U3373 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8010 = ~(P2_U3332 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8012 = ~(P2_U3362 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8014 = ~(P2_U3346 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8016 = ~(P2_U3398 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8018 = ~(P2_U3386 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8021 = ~(P2_U3420 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8023 = ~(P2_U3409 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8024 = ~(P2_U3372 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8026 = ~(P2_U3331 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8028 = ~(P2_U3361 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8030 = ~(P2_U3345 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8032 = ~(P2_U3397 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8034 = ~(P2_U3382 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8037 = ~(P2_U3416 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8039 = ~(P2_U3405 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8040 = ~(P2_U3368 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8042 = ~(P2_U3327 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8044 = ~(P2_U3357 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8046 = ~(P2_U3341 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8048 = ~(P2_U3393 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8056 = U211 | P2_STATE2_REG_0__SCAN_IN; 
assign P2_U8065 = ~(P2_U3311 & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P2_U8079 = ~(P2_U4591 & P2_U3276 & P2_U3273); 
assign P2_U8080 = ~(P2_U3277 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8098 = ~(P2_U3271 & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P2_U8099 = ~(P2_U3272 & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P2_U8150 = ~(P2_U3273 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P2_U8151 = ~(P2_U3276 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8281 = ~(P2_U3519 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P2_U8283 = ~(P2_U3519 & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P2_U8285 = ~(P2_U3519 & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P2_U8419 = ~(P2_R2337_U4 & P2_U3284); 
assign P2_U8421 = ~(P2_U3284 & P2_PHYADDRPOINTER_REG_0__SCAN_IN); 
assign P1_U2430 = P1_U3387 & P1_STATE2_REG_1__SCAN_IN; 
assign P1_U2454 = P1_U3266 & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P1_U2455 = P1_U3266 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P1_U2456 = P1_U3265 & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_U2457 = P1_U3265 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_U2459 = P1_U3264 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_U2460 = P1_U3264 & P1_U3266 & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P1_U2461 = P1_U3506 & P1_U3505; 
assign P1_U2462 = P1_U3264 & P1_U3265 & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_U2463 = P1_U3504 & P1_U3503; 
assign P1_U2465 = P1_U3502 & P1_U3501; 
assign P1_U2466 = P1_U3500 & P1_U3499; 
assign P1_U2468 = P1_U3498 & P1_U3497; 
assign P1_U2470 = P1_U3266 & P1_U2469 & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P1_U2471 = P1_U3265 & P1_U2469 & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_U2479 = P1_U3303 & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign P1_U3249 = ~(P1_U3258 & P1_STATE_REG_1__SCAN_IN); 
assign P1_U3254 = ~(P1_U3251 & P1_STATE_REG_1__SCAN_IN); 
assign P1_U3257 = ~U210; 
assign P1_U3260 = ~(P1_U3256 & P1_REQUESTPENDING_REG_SCAN_IN); 
assign P1_U3267 = ~(P1_U3270 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U3274 = ~(P1_U3270 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_U3280 = U210 | P1_STATEBS16_REG_SCAN_IN; 
assign P1_U3297 = ~(P1_U3262 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U3323 = ~(P1_U3301 & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P1_U3329 = ~(P1_U3302 & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P1_U3337 = ~(P1_U2488 & P1_U2478); 
assign P1_U3340 = ~(P1_U3304 & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P1_U3384 = ~(P1_U2510 & P1_U2488); 
assign P1_U3402 = ~(P1_U3269 & P1_U3275); 
assign P1_U3408 = ~(P1_U2427 & P1_U3294); 
assign P1_U3440 = ~(P1_U3263 & P1_STATEBS16_REG_SCAN_IN); 
assign P1_U3444 = ~(P1_U3264 & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U3463 = P1_U3255 & P1_U4179; 
assign P1_U3888 = ~(U210 | P1_STATEBS16_REG_SCAN_IN); 
assign P1_U3952 = P1_U3951 & P1_U3950; 
assign P1_U3955 = P1_U3954 & P1_U3953; 
assign P1_U3958 = P1_U3957 & P1_U3956; 
assign P1_U3962 = P1_U3961 & P1_U6598 & P1_U3960 & P1_U3959; 
assign P1_U3966 = ~(U210 | P1_STATE2_REG_0__SCAN_IN); 
assign P1_U4157 = P1_U2427 & P1_STATE2_REG_0__SCAN_IN; 
assign P1_U4183 = ~(P1_U3269 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_U4209 = ~P1_U3307; 
assign P1_U4242 = ~(P1_U3731 & P1_U2428); 
assign P1_U4244 = ~(P1_U3294 & P1_U2352 & P1_STATE2_REG_1__SCAN_IN); 
assign P1_U4246 = ~(P1_U3263 & U210 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U4261 = ~P1_U3298; 
assign P1_U4360 = ~P1_U3261; 
assign P1_U4364 = ~P1_U3255; 
assign P1_U4366 = ~(P1_U3261 & U210 & P1_STATE_REG_1__SCAN_IN); 
assign P1_U4373 = ~(NA & P1_U3258); 
assign P1_U4376 = ~(P1_U4179 & P1_U3255); 
assign P1_U4378 = ~P1_U3269; 
assign P1_U4380 = ~P1_U3268; 
assign P1_U4398 = ~(P1_U2453 & P1_INSTQUEUE_REG_15__3__SCAN_IN); 
assign P1_U4401 = ~(P1_U3270 & P1_INSTQUEUE_REG_7__5__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U4403 = ~(P1_U2469 & P1_U3265 & P1_INSTQUEUE_REG_1__5__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U4404 = ~(P1_U2469 & P1_U3266 & P1_INSTQUEUE_REG_2__5__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U4406 = ~(P1_U3520 & P1_U3521 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_U4407 = ~(P1_U3522 & P1_U3523 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_U4409 = ~(P1_U3525 & P1_U3526 & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U4410 = ~(P1_U3264 & P1_INSTQUEUE_REG_11__5__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U4412 = ~(P1_U3265 & P1_INSTQUEUE_REG_13__5__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U4413 = ~(P1_U3266 & P1_INSTQUEUE_REG_14__5__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U4431 = ~(P1_U2453 & P1_INSTQUEUE_REG_15__2__SCAN_IN); 
assign P1_U4448 = ~(P1_U2453 & P1_INSTQUEUE_REG_15__7__SCAN_IN); 
assign P1_U4459 = ~(P1_U3507 & P1_U3498 & P1_INSTQUEUE_REG_15__6__SCAN_IN); 
assign P1_U4476 = ~(P1_U2453 & P1_INSTQUEUE_REG_15__1__SCAN_IN); 
assign P1_U4493 = ~(P1_U2453 & P1_INSTQUEUE_REG_15__0__SCAN_IN); 
assign P1_U4495 = ~(P1_U3248 & P1_STATE_REG_2__SCAN_IN); 
assign P1_U4513 = ~(U210 & P1_STATE2_REG_1__SCAN_IN); 
assign P1_U4533 = ~P1_U3305; 
assign P1_U4539 = ~(P1_U3305 & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P1_U4546 = ~(P1_U3263 & P1_STATE2_REG_1__SCAN_IN); 
assign P1_U5475 = ~(P1_U3294 & P1_STATE2_REG_3__SCAN_IN); 
assign P1_U5478 = ~(P1_U5477 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P1_U5481 = ~(P1_U3498 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_U5484 = ~(P1_U3275 & P1_U3264); 
assign P1_U5486 = ~(P1_U2469 & P1_U3275); 
assign P1_U5510 = ~(P1_U3275 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_U5538 = ~(P1_U3296 & P1_STATE2_REG_1__SCAN_IN); 
assign P1_U5796 = ~(P1_U3294 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U5797 = ~(P1_U3308 & P1_STATE2_REG_1__SCAN_IN); 
assign P1_U6054 = ~(P1_U2428 & P1_U3294); 
assign P1_U6367 = U210 | P1_STATEBS16_REG_SCAN_IN; 
assign P1_U6862 = ~(P1_R2337_U4 & P1_U2352); 
assign P1_U6867 = ~(P1_U2352 & P1_PHYADDRPOINTER_REG_0__SCAN_IN); 
assign P1_U7064 = ~(P1_U3264 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P1_U7377 = ~(P1_U3294 & P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P1_U7379 = ~(P1_U3294 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P1_U7383 = ~(P1_U3294 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_U7386 = ~(P1_U3294 & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U7389 = ~(P1_U3294 & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U7469 = U210 | P1_STATE2_REG_2__SCAN_IN; 
assign P1_U7641 = ~(P1_U3251 & P1_STATE_REG_0__SCAN_IN & P1_REQUESTPENDING_REG_SCAN_IN); 
assign P1_U7655 = ~(P1_U3541 & P1_U3540 & P1_U3265); 
assign P1_U7656 = ~(P1_U3270 & P1_INSTQUEUE_REG_7__4__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U7657 = ~(P1_U3270 & P1_U3265 & P1_INSTQUEUE_REG_5__4__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U7658 = ~(P1_U3270 & P1_U3264 & P1_U3266 & P1_INSTQUEUE_REG_2__4__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U7659 = ~(P1_U3543 & P1_U3542 & P1_U3270); 
assign P1_U7660 = ~(P1_U3545 & P1_U3544 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P1_U7661 = ~(P1_U3547 & P1_U3546 & P1_U3265); 
assign P1_U7662 = ~(P1_U3549 & P1_U3548 & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U7663 = ~(P1_U3551 & P1_U3550 & P1_U3266); 
assign P1_U7665 = ~(P1_U3264 & P1_U3265 & P1_U3266 & P1_U3270 & P1_INSTQUEUE_REG_0__4__SCAN_IN); 
assign P1_U7666 = ~(P1_U3264 & P1_U3265 & P1_U3266 & P1_INSTQUEUE_REG_8__4__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P1_U7667 = ~(P1_U3264 & P1_U3266 & P1_INSTQUEUE_REG_10__4__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U7668 = ~(P1_U3553 & P1_U3552 & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U7669 = ~(P1_U3264 & P1_U3270 & P1_INSTQUEUE_REG_3__4__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U7670 = ~(P1_U3264 & P1_INSTQUEUE_REG_11__4__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U7671 = ~(P1_U3264 & P1_U3270 & P1_INSTQUEUE_REG_3__5__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U7672 = ~(P1_U3529 & P1_U3528 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P1_U7673 = ~(P1_U3264 & P1_U3265 & P1_INSTQUEUE_REG_9__6__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U7674 = ~(P1_U3535 & P1_U3534 & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U7675 = ~(P1_U3264 & P1_U3266 & P1_INSTQUEUE_REG_10__6__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U7676 = ~(P1_U3264 & P1_INSTQUEUE_REG_11__6__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U7677 = ~(P1_U3264 & P1_U3265 & P1_U3266 & P1_U3270 & P1_INSTQUEUE_REG_0__6__SCAN_IN); 
assign P1_U7678 = ~(P1_U3264 & P1_U3265 & P1_U3266 & P1_INSTQUEUE_REG_8__6__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P1_U7694 = ~(P1_U3305 & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P1_U7710 = ~(P1_U4174 & P1_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P1_U7713 = ~(P1_U4174 & P1_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P1_U7718 = ~(P1_U3264 & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U7719 = ~(P1_U3265 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_U7749 = ~(P1_U3413 & P1_DATAWIDTH_REG_0__SCAN_IN); 
assign LT_782_120_U6 = ~(LT_782_120_U7 & P3_DATAO_REG_30__SCAN_IN); 
assign LT_782_U6 = ~(LT_782_U7 & P1_DATAO_REG_30__SCAN_IN); 
assign R170_U8 = ~(R170_U7 | P2_ADDRESS_REG_25__SCAN_IN | P2_ADDRESS_REG_24__SCAN_IN | P2_ADDRESS_REG_19__SCAN_IN | P2_ADDRESS_REG_10__SCAN_IN); 
assign R170_U10 = ~(R170_U9 | P2_ADDRESS_REG_23__SCAN_IN | P2_ADDRESS_REG_11__SCAN_IN | P2_ADDRESS_REG_1__SCAN_IN); 
assign R170_U12 = ~(R170_U11 | P2_ADDRESS_REG_14__SCAN_IN | P2_ADDRESS_REG_12__SCAN_IN | P2_ADDRESS_REG_4__SCAN_IN); 
assign R170_U14 = ~(R170_U13 | P2_ADDRESS_REG_15__SCAN_IN | P2_ADDRESS_REG_5__SCAN_IN | P2_ADDRESS_REG_2__SCAN_IN); 
assign R165_U8 = ~(R165_U7 | P1_ADDRESS_REG_25__SCAN_IN | P1_ADDRESS_REG_24__SCAN_IN | P1_ADDRESS_REG_19__SCAN_IN | P1_ADDRESS_REG_10__SCAN_IN); 
assign R165_U10 = ~(R165_U9 | P1_ADDRESS_REG_23__SCAN_IN | P1_ADDRESS_REG_11__SCAN_IN | P1_ADDRESS_REG_1__SCAN_IN); 
assign R165_U12 = ~(R165_U11 | P1_ADDRESS_REG_14__SCAN_IN | P1_ADDRESS_REG_12__SCAN_IN | P1_ADDRESS_REG_4__SCAN_IN); 
assign R165_U14 = ~(R165_U13 | P1_ADDRESS_REG_15__SCAN_IN | P1_ADDRESS_REG_5__SCAN_IN | P1_ADDRESS_REG_2__SCAN_IN); 
assign LT_782_119_U6 = ~(LT_782_119_U7 & P2_DATAO_REG_30__SCAN_IN); 
assign P3_ADD_526_U111 = ~P3_ADD_526_U10; 
assign P3_ADD_526_U130 = ~P3_ADD_526_U100; 
assign P3_ADD_526_U154 = ~(P3_ADD_526_U10 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_526_U159 = ~(P3_ADD_526_U100 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_526_U181 = ~(P3_ADD_526_U7 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_ADD_526_U182 = ~(P3_ADD_526_U5 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_552_U111 = ~P3_ADD_552_U10; 
assign P3_ADD_552_U130 = ~P3_ADD_552_U100; 
assign P3_ADD_552_U154 = ~(P3_ADD_552_U10 & P3_EBX_REG_3__SCAN_IN); 
assign P3_ADD_552_U159 = ~(P3_ADD_552_U100 & P3_EBX_REG_2__SCAN_IN); 
assign P3_ADD_552_U181 = ~(P3_ADD_552_U7 & P3_EBX_REG_0__SCAN_IN); 
assign P3_ADD_552_U182 = ~(P3_ADD_552_U5 & P3_EBX_REG_1__SCAN_IN); 
assign P3_ADD_546_U111 = ~P3_ADD_546_U10; 
assign P3_ADD_546_U130 = ~P3_ADD_546_U100; 
assign P3_ADD_546_U154 = ~(P3_ADD_546_U10 & P3_EAX_REG_3__SCAN_IN); 
assign P3_ADD_546_U159 = ~(P3_ADD_546_U100 & P3_EAX_REG_2__SCAN_IN); 
assign P3_ADD_546_U181 = ~(P3_ADD_546_U7 & P3_EAX_REG_0__SCAN_IN); 
assign P3_ADD_546_U182 = ~(P3_ADD_546_U5 & P3_EAX_REG_1__SCAN_IN); 
assign P3_ADD_476_U94 = ~P3_ADD_476_U6; 
assign P3_ADD_476_U135 = ~(P3_ADD_476_U6 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_476_U141 = ~(P3_ADD_476_U4 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_476_U142 = ~(P3_ADD_476_U5 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_531_U98 = ~P3_ADD_531_U7; 
assign P3_ADD_531_U146 = ~(P3_ADD_531_U7 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_531_U168 = ~(P3_ADD_531_U5 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_531_U169 = ~(P3_ADD_531_U6 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_SUB_320_U71 = ~P3_ADD_318_U4; 
assign P3_SUB_320_U104 = P3_ADD_318_U4 | P3_PHYADDRPOINTER_REG_0__SCAN_IN; 
assign P3_SUB_320_U148 = ~(P3_ADD_318_U4 & P3_SUB_320_U72); 
assign P3_ADD_505_U18 = ~P3_ADD_505_U8; 
assign P3_ADD_505_U25 = ~(P3_ADD_505_U8 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_ADD_505_U27 = ~(P3_ADD_505_U5 & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P3_ADD_505_U28 = ~(P3_ADD_505_U7 & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P3_ADD_318_U94 = ~P3_ADD_318_U6; 
assign P3_ADD_318_U135 = ~(P3_ADD_318_U6 & P3_PHYADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_318_U141 = ~(P3_ADD_318_U4 & P3_PHYADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_318_U142 = ~(P3_ADD_318_U5 & P3_PHYADDRPOINTER_REG_1__SCAN_IN); 
assign P3_SUB_370_U9 = ~(P3_SUB_370_U18 & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P3_SUB_370_U35 = ~(P3_SUB_370_U12 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_370_U37 = ~(P3_SUB_370_U11 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_370_U39 = ~(P3_SUB_370_U14 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_370_U41 = ~(P3_SUB_370_U13 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_370_U43 = ~(P3_SUB_370_U17 & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_370_U45 = ~(P3_SUB_370_U15 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_370_U46 = ~(P3_SUB_370_U8 & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P3_SUB_370_U47 = ~(P3_SUB_370_U15 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_370_U48 = ~(P3_SUB_370_U17 & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_370_U52 = ~(P3_SUB_370_U14 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_370_U53 = ~(P3_SUB_370_U13 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_370_U57 = ~(P3_SUB_370_U12 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_370_U58 = ~(P3_SUB_370_U11 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_370_U62 = ~(P3_SUB_370_U10 & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P3_SUB_370_U63 = ~(P3_SUB_370_U29 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_ADD_315_U91 = ~P3_ADD_315_U6; 
assign P3_ADD_315_U129 = ~(P3_ADD_315_U6 & P3_PHYADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_315_U131 = ~(P3_ADD_315_U4 & P3_PHYADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_315_U132 = ~(P3_ADD_315_U5 & P3_PHYADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_467_U94 = ~P3_ADD_467_U6; 
assign P3_ADD_467_U135 = ~(P3_ADD_467_U6 & P3_REIP_REG_3__SCAN_IN); 
assign P3_ADD_467_U141 = ~(P3_ADD_467_U4 & P3_REIP_REG_2__SCAN_IN); 
assign P3_ADD_467_U142 = ~(P3_ADD_467_U5 & P3_REIP_REG_1__SCAN_IN); 
assign P3_ADD_430_U94 = ~P3_ADD_430_U6; 
assign P3_ADD_430_U135 = ~(P3_ADD_430_U6 & P3_REIP_REG_3__SCAN_IN); 
assign P3_ADD_430_U141 = ~(P3_ADD_430_U4 & P3_REIP_REG_2__SCAN_IN); 
assign P3_ADD_430_U142 = ~(P3_ADD_430_U5 & P3_REIP_REG_1__SCAN_IN); 
assign P3_ADD_380_U98 = ~P3_ADD_380_U7; 
assign P3_ADD_380_U146 = ~(P3_ADD_380_U7 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_380_U168 = ~(P3_ADD_380_U5 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_380_U169 = ~(P3_ADD_380_U6 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_ADD_344_U98 = ~P3_ADD_344_U7; 
assign P3_ADD_344_U146 = ~(P3_ADD_344_U7 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_344_U168 = ~(P3_ADD_344_U5 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_344_U169 = ~(P3_ADD_344_U6 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_ADD_339_U94 = ~P3_ADD_339_U6; 
assign P3_ADD_339_U135 = ~(P3_ADD_339_U6 & P3_PHYADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_339_U141 = ~(P3_ADD_339_U4 & P3_PHYADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_339_U142 = ~(P3_ADD_339_U5 & P3_PHYADDRPOINTER_REG_1__SCAN_IN); 
assign P3_SUB_580_U9 = ~(P3_SUB_580_U8 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_SUB_580_U10 = ~(P3_SUB_580_U7 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_ADD_541_U94 = ~P3_ADD_541_U6; 
assign P3_ADD_541_U135 = ~(P3_ADD_541_U6 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_541_U141 = ~(P3_ADD_541_U4 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_541_U142 = ~(P3_ADD_541_U5 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_SUB_355_U9 = ~(P3_SUB_355_U18 & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P3_SUB_355_U35 = ~(P3_SUB_355_U12 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_355_U37 = ~(P3_SUB_355_U11 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_355_U39 = ~(P3_SUB_355_U14 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_355_U41 = ~(P3_SUB_355_U13 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_355_U43 = ~(P3_SUB_355_U17 & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_355_U45 = ~(P3_SUB_355_U15 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_355_U46 = ~(P3_SUB_355_U8 & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P3_SUB_355_U47 = ~(P3_SUB_355_U15 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_355_U48 = ~(P3_SUB_355_U17 & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_355_U52 = ~(P3_SUB_355_U14 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_355_U53 = ~(P3_SUB_355_U13 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_355_U57 = ~(P3_SUB_355_U12 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_355_U58 = ~(P3_SUB_355_U11 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_355_U62 = ~(P3_SUB_355_U10 & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P3_SUB_355_U63 = ~(P3_SUB_355_U29 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_SUB_450_U7 = ~(P3_SUB_450_U27 & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P3_SUB_450_U33 = ~(P3_SUB_450_U10 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_450_U35 = ~(P3_SUB_450_U9 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_450_U37 = ~(P3_SUB_450_U12 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_450_U39 = ~(P3_SUB_450_U11 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_450_U41 = ~(P3_SUB_450_U15 & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_450_U43 = ~(P3_SUB_450_U13 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_450_U44 = ~(P3_SUB_450_U13 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_450_U45 = ~(P3_SUB_450_U15 & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_450_U49 = ~(P3_SUB_450_U12 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_450_U50 = ~(P3_SUB_450_U11 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_450_U54 = ~(P3_SUB_450_U10 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_450_U55 = ~(P3_SUB_450_U9 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_450_U59 = ~(P3_SUB_450_U8 & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P3_SUB_450_U60 = ~(P3_SUB_450_U26 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_SUB_357_1258_U207 = ~P3_SUB_357_1258_U57; 
assign P3_ADD_486_U18 = ~P3_ADD_486_U8; 
assign P3_ADD_486_U25 = ~(P3_ADD_486_U8 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_ADD_486_U27 = ~(P3_ADD_486_U5 & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P3_ADD_486_U28 = ~(P3_ADD_486_U7 & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P3_SUB_485_U7 = ~(P3_SUB_485_U27 & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P3_SUB_485_U33 = ~(P3_SUB_485_U10 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_485_U35 = ~(P3_SUB_485_U9 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_485_U37 = ~(P3_SUB_485_U12 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_485_U39 = ~(P3_SUB_485_U11 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_485_U41 = ~(P3_SUB_485_U15 & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_485_U43 = ~(P3_SUB_485_U13 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_485_U44 = ~(P3_SUB_485_U13 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_485_U45 = ~(P3_SUB_485_U15 & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_485_U49 = ~(P3_SUB_485_U12 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_485_U50 = ~(P3_SUB_485_U11 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_485_U54 = ~(P3_SUB_485_U10 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_485_U55 = ~(P3_SUB_485_U9 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_485_U59 = ~(P3_SUB_485_U8 & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P3_SUB_485_U60 = ~(P3_SUB_485_U26 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_ADD_515_U94 = ~P3_ADD_515_U6; 
assign P3_ADD_515_U135 = ~(P3_ADD_515_U6 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_515_U141 = ~(P3_ADD_515_U4 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_515_U142 = ~(P3_ADD_515_U5 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_394_U92 = ~(P3_ADD_394_U62 & P3_ADD_394_U96); 
assign P3_ADD_394_U165 = ~(P3_ADD_394_U4 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_394_U166 = ~(P3_ADD_394_U6 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_SUB_414_U83 = ~P3_SUB_414_U21; 
assign P3_SUB_414_U105 = ~(P3_SUB_414_U104 & P3_EBX_REG_2__SCAN_IN); 
assign P3_SUB_414_U134 = ~(P3_SUB_414_U21 & P3_EBX_REG_3__SCAN_IN); 
assign P3_SUB_414_U148 = ~(P3_SUB_414_U72 & P3_EBX_REG_1__SCAN_IN); 
assign P3_SUB_414_U149 = ~(P3_SUB_414_U71 & P3_EBX_REG_0__SCAN_IN); 
assign P3_ADD_441_U94 = ~P3_ADD_441_U6; 
assign P3_ADD_441_U135 = ~(P3_ADD_441_U6 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_441_U141 = ~(P3_ADD_441_U4 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_441_U142 = ~(P3_ADD_441_U5 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_349_U98 = ~P3_ADD_349_U7; 
assign P3_ADD_349_U146 = ~(P3_ADD_349_U7 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_349_U168 = ~(P3_ADD_349_U5 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_349_U169 = ~(P3_ADD_349_U6 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_ADD_405_U92 = ~(P3_ADD_405_U62 & P3_ADD_405_U96); 
assign P3_ADD_405_U165 = ~(P3_ADD_405_U4 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_405_U166 = ~(P3_ADD_405_U6 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_ADD_553_U98 = ~P3_ADD_553_U7; 
assign P3_ADD_553_U146 = ~(P3_ADD_553_U7 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_553_U168 = ~(P3_ADD_553_U5 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_553_U169 = ~(P3_ADD_553_U6 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_ADD_558_U98 = ~P3_ADD_558_U7; 
assign P3_ADD_558_U146 = ~(P3_ADD_558_U7 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_558_U168 = ~(P3_ADD_558_U5 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_558_U169 = ~(P3_ADD_558_U6 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_ADD_385_U98 = ~P3_ADD_385_U7; 
assign P3_ADD_385_U146 = ~(P3_ADD_385_U7 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_385_U168 = ~(P3_ADD_385_U5 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_385_U169 = ~(P3_ADD_385_U6 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_ADD_547_U98 = ~P3_ADD_547_U7; 
assign P3_ADD_547_U146 = ~(P3_ADD_547_U7 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_547_U168 = ~(P3_ADD_547_U5 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_547_U169 = ~(P3_ADD_547_U6 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_SUB_412_U7 = ~(P3_SUB_412_U27 & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P3_SUB_412_U33 = ~(P3_SUB_412_U10 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_412_U35 = ~(P3_SUB_412_U9 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_412_U37 = ~(P3_SUB_412_U12 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_412_U39 = ~(P3_SUB_412_U11 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_412_U41 = ~(P3_SUB_412_U15 & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_412_U43 = ~(P3_SUB_412_U13 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_412_U44 = ~(P3_SUB_412_U13 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_412_U45 = ~(P3_SUB_412_U15 & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_412_U49 = ~(P3_SUB_412_U12 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_412_U50 = ~(P3_SUB_412_U11 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_412_U54 = ~(P3_SUB_412_U10 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_412_U55 = ~(P3_SUB_412_U9 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_412_U59 = ~(P3_SUB_412_U8 & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P3_SUB_412_U60 = ~(P3_SUB_412_U26 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_SUB_504_U7 = ~(P3_SUB_504_U27 & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P3_SUB_504_U33 = ~(P3_SUB_504_U10 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_504_U35 = ~(P3_SUB_504_U9 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_504_U37 = ~(P3_SUB_504_U12 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_504_U39 = ~(P3_SUB_504_U11 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_504_U41 = ~(P3_SUB_504_U15 & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_504_U43 = ~(P3_SUB_504_U13 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_504_U44 = ~(P3_SUB_504_U13 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_504_U45 = ~(P3_SUB_504_U15 & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_504_U49 = ~(P3_SUB_504_U12 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_504_U50 = ~(P3_SUB_504_U11 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_504_U54 = ~(P3_SUB_504_U10 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_504_U55 = ~(P3_SUB_504_U9 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_504_U59 = ~(P3_SUB_504_U8 & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P3_SUB_504_U60 = ~(P3_SUB_504_U26 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_SUB_401_U9 = ~(P3_SUB_401_U18 & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P3_SUB_401_U35 = ~(P3_SUB_401_U12 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_401_U37 = ~(P3_SUB_401_U11 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_401_U39 = ~(P3_SUB_401_U14 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_401_U41 = ~(P3_SUB_401_U13 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_401_U43 = ~(P3_SUB_401_U17 & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_401_U45 = ~(P3_SUB_401_U15 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_401_U46 = ~(P3_SUB_401_U8 & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P3_SUB_401_U47 = ~(P3_SUB_401_U15 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_401_U48 = ~(P3_SUB_401_U17 & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_401_U52 = ~(P3_SUB_401_U14 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_401_U53 = ~(P3_SUB_401_U13 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_401_U57 = ~(P3_SUB_401_U12 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_401_U58 = ~(P3_SUB_401_U11 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_401_U62 = ~(P3_SUB_401_U10 & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P3_SUB_401_U63 = ~(P3_SUB_401_U29 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_SUB_390_U9 = ~(P3_SUB_390_U18 & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P3_SUB_390_U35 = ~(P3_SUB_390_U12 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_390_U37 = ~(P3_SUB_390_U11 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_390_U39 = ~(P3_SUB_390_U14 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_390_U41 = ~(P3_SUB_390_U13 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_390_U43 = ~(P3_SUB_390_U17 & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_390_U45 = ~(P3_SUB_390_U15 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_390_U46 = ~(P3_SUB_390_U8 & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P3_SUB_390_U47 = ~(P3_SUB_390_U15 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_390_U48 = ~(P3_SUB_390_U17 & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_390_U52 = ~(P3_SUB_390_U14 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_390_U53 = ~(P3_SUB_390_U13 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_390_U57 = ~(P3_SUB_390_U12 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_390_U58 = ~(P3_SUB_390_U11 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_SUB_390_U62 = ~(P3_SUB_390_U10 & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P3_SUB_390_U63 = ~(P3_SUB_390_U29 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_ADD_495_U13 = ~P3_ADD_495_U6; 
assign P3_ADD_495_U17 = ~(P3_ADD_495_U6 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_ADD_495_U19 = ~(P3_ADD_495_U4 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_ADD_495_U20 = ~(P3_ADD_495_U5 & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P3_ADD_494_U94 = ~P3_ADD_494_U6; 
assign P3_ADD_494_U135 = ~(P3_ADD_494_U6 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_494_U141 = ~(P3_ADD_494_U4 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_494_U142 = ~(P3_ADD_494_U5 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_536_U94 = ~P3_ADD_536_U6; 
assign P3_ADD_536_U135 = ~(P3_ADD_536_U6 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_536_U141 = ~(P3_ADD_536_U4 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_536_U142 = ~(P3_ADD_536_U5 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P2_R2027_U98 = ~P2_R2027_U7; 
assign P2_R2027_U146 = ~(P2_R2027_U7 & P2_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P2_R2027_U168 = ~(P2_R2027_U5 & P2_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P2_R2027_U169 = ~(P2_R2027_U6 & P2_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P2_R2337_U94 = ~P2_R2337_U91; 
assign P2_R2337_U95 = ~P2_R2337_U7; 
assign P2_R2337_U133 = ~(P2_R2337_U7 & P2_PHYADDRPOINTER_REG_4__SCAN_IN); 
assign P2_R2337_U135 = ~(P2_R2337_U91 & P2_PHYADDRPOINTER_REG_3__SCAN_IN); 
assign P2_R2337_U141 = ~(P2_R2337_U4 & P2_PHYADDRPOINTER_REG_2__SCAN_IN); 
assign P2_R2337_U142 = ~(P2_R2337_U6 & P2_PHYADDRPOINTER_REG_1__SCAN_IN); 
assign P2_R2147_U13 = ~P2_R2147_U11; 
assign P2_R2147_U14 = ~P2_R2147_U12; 
assign P2_R2147_U17 = ~(P2_R2147_U12 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_R2147_U19 = ~(P2_R2147_U4 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P2_R2147_U20 = ~(P2_R2147_U6 & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P2_R2238_U9 = ~(P2_R2238_U18 & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P2_R2238_U35 = ~(P2_R2238_U12 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P2_R2238_U37 = ~(P2_R2238_U11 & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P2_R2238_U39 = ~(P2_R2238_U14 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_R2238_U41 = ~(P2_R2238_U13 & P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P2_R2238_U43 = ~(P2_R2238_U17 & P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P2_R2238_U45 = ~(P2_R2238_U15 & P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P2_R2238_U46 = ~(P2_R2238_U8 & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P2_R2238_U47 = ~(P2_R2238_U15 & P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P2_R2238_U48 = ~(P2_R2238_U17 & P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P2_R2238_U52 = ~(P2_R2238_U14 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_R2238_U53 = ~(P2_R2238_U13 & P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P2_R2238_U57 = ~(P2_R2238_U12 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P2_R2238_U58 = ~(P2_R2238_U11 & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P2_R2238_U62 = ~(P2_R2238_U10 & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P2_R2238_U63 = ~(P2_R2238_U29 & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P2_SUB_450_U7 = ~(P2_SUB_450_U16 & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P2_SUB_450_U33 = ~(P2_SUB_450_U10 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P2_SUB_450_U35 = ~(P2_SUB_450_U9 & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P2_SUB_450_U37 = ~(P2_SUB_450_U12 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_SUB_450_U39 = ~(P2_SUB_450_U11 & P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P2_SUB_450_U41 = ~(P2_SUB_450_U15 & P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P2_SUB_450_U43 = ~(P2_SUB_450_U13 & P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P2_SUB_450_U44 = ~(P2_SUB_450_U13 & P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P2_SUB_450_U45 = ~(P2_SUB_450_U15 & P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P2_SUB_450_U49 = ~(P2_SUB_450_U12 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_SUB_450_U50 = ~(P2_SUB_450_U11 & P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P2_SUB_450_U54 = ~(P2_SUB_450_U10 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P2_SUB_450_U55 = ~(P2_SUB_450_U9 & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P2_SUB_450_U59 = ~(P2_SUB_450_U8 & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P2_SUB_450_U60 = ~(P2_SUB_450_U27 & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P2_ADD_394_U94 = ~(P2_ADD_394_U62 & P2_ADD_394_U96); 
assign P2_ADD_394_U173 = ~(P2_ADD_394_U4 & P2_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P2_ADD_394_U174 = ~(P2_ADD_394_U6 & P2_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P2_ADD_371_1212_U4 = P2_ADD_371_1212_U10 & P2_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P2_ADD_371_1212_U7 = P2_ADD_371_1212_U10 & P2_ADD_371_1212_U87; 
assign P2_ADD_371_1212_U102 = P2_ADD_371_1212_U5 & P2_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P1_R2027_U111 = ~P1_R2027_U10; 
assign P1_R2027_U130 = ~P1_R2027_U100; 
assign P1_R2027_U154 = ~(P1_R2027_U10 & P1_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P1_R2027_U159 = ~(P1_R2027_U100 & P1_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P1_R2027_U181 = ~(P1_R2027_U7 & P1_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P1_R2027_U182 = ~(P1_R2027_U5 & P1_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P1_R2358_U23 = ~P1_U2352; 
assign P1_R2337_U94 = ~P1_R2337_U6; 
assign P1_R2337_U135 = ~(P1_R2337_U6 & P1_PHYADDRPOINTER_REG_3__SCAN_IN); 
assign P1_R2337_U141 = ~(P1_R2337_U4 & P1_PHYADDRPOINTER_REG_2__SCAN_IN); 
assign P1_R2337_U142 = ~(P1_R2337_U5 & P1_PHYADDRPOINTER_REG_1__SCAN_IN); 
assign P1_SUB_580_U9 = ~(P1_SUB_580_U8 & P1_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P1_SUB_580_U10 = ~(P1_SUB_580_U7 & P1_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P1_R2096_U94 = ~P1_R2096_U6; 
assign P1_R2096_U135 = ~(P1_R2096_U6 & P1_REIP_REG_3__SCAN_IN); 
assign P1_R2096_U141 = ~(P1_R2096_U4 & P1_REIP_REG_2__SCAN_IN); 
assign P1_R2096_U142 = ~(P1_R2096_U5 & P1_REIP_REG_1__SCAN_IN); 
assign P1_R2238_U9 = ~(P1_R2238_U18 & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_R2238_U35 = ~(P1_R2238_U12 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_R2238_U37 = ~(P1_R2238_U11 & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P1_R2238_U39 = ~(P1_R2238_U14 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P1_R2238_U41 = ~(P1_R2238_U13 & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P1_R2238_U43 = ~(P1_R2238_U17 & P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P1_R2238_U45 = ~(P1_R2238_U15 & P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P1_R2238_U46 = ~(P1_R2238_U8 & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P1_R2238_U47 = ~(P1_R2238_U15 & P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P1_R2238_U48 = ~(P1_R2238_U17 & P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P1_R2238_U52 = ~(P1_R2238_U14 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P1_R2238_U53 = ~(P1_R2238_U13 & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P1_R2238_U57 = ~(P1_R2238_U12 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_R2238_U58 = ~(P1_R2238_U11 & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P1_R2238_U62 = ~(P1_R2238_U10 & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_R2238_U63 = ~(P1_R2238_U29 & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P1_SUB_450_U9 = ~(P1_SUB_450_U18 & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_SUB_450_U35 = ~(P1_SUB_450_U12 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_SUB_450_U37 = ~(P1_SUB_450_U11 & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P1_SUB_450_U39 = ~(P1_SUB_450_U14 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P1_SUB_450_U41 = ~(P1_SUB_450_U13 & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P1_SUB_450_U43 = ~(P1_SUB_450_U17 & P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P1_SUB_450_U45 = ~(P1_SUB_450_U15 & P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P1_SUB_450_U46 = ~(P1_SUB_450_U8 & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P1_SUB_450_U47 = ~(P1_SUB_450_U15 & P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P1_SUB_450_U48 = ~(P1_SUB_450_U17 & P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P1_SUB_450_U52 = ~(P1_SUB_450_U14 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P1_SUB_450_U53 = ~(P1_SUB_450_U13 & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P1_SUB_450_U57 = ~(P1_SUB_450_U12 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_SUB_450_U58 = ~(P1_SUB_450_U11 & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P1_SUB_450_U62 = ~(P1_SUB_450_U10 & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_SUB_450_U63 = ~(P1_SUB_450_U29 & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P1_ADD_405_U94 = ~(P1_ADD_405_U62 & P1_ADD_405_U96); 
assign P1_ADD_405_U173 = ~(P1_ADD_405_U4 & P1_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P1_ADD_405_U174 = ~(P1_ADD_405_U6 & P1_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P1_ADD_515_U94 = ~P1_ADD_515_U6; 
assign P1_ADD_515_U133 = ~(P1_ADD_515_U4 & P1_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P1_ADD_515_U134 = ~(P1_ADD_515_U5 & P1_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P1_ADD_515_U169 = ~(P1_ADD_515_U6 & P1_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign U215 = ~(LT_748_U6 & U208); 
assign U382 = ~(LT_782_120_U6 & LT_782_U6 & LT_782_119_U6); 
assign P3_U2465 = P3_U2464 & P3_U4332; 
assign P3_U2467 = P3_U2464 & P3_U2466; 
assign P3_U2469 = P3_U2464 & P3_U2468; 
assign P3_U2470 = P3_U2464 & P3_U4467; 
assign P3_U2472 = P3_U2466 & P3_U3097; 
assign P3_U2474 = P3_U2468 & P3_U3097; 
assign P3_U2482 = P3_U2466 & P3_U2481; 
assign P3_U2483 = P3_U2468 & P3_U2481; 
assign P3_U2519 = P3_U3228 & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P3_U2522 = P3_U3093 & P3_U3228; 
assign P3_U3086 = ~(P3_U3087 & P3_STATE_REG_0__SCAN_IN); 
assign P3_U3092 = ~(P3_U4467 & P3_U3097); 
assign P3_U3096 = ~(P3_U4332 & P3_U3097); 
assign P3_U3132 = ~(P3_U4648 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_U3136 = ~(P3_U4295 & P3_STATEBS16_REG_SCAN_IN); 
assign P3_U3137 = ~(P3_U3153 & P3_U4641); 
assign P3_U3147 = ~(P3_U3386 & P3_U2492); 
assign P3_U3161 = ~(P3_U3422 & P3_U2492); 
assign P3_U3164 = ~(P3_U3131 & P3_U4648 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_U3186 = ~(P3_U3527 & P3_U2492); 
assign P3_U3194 = ~(P3_U3563 & P3_U2492); 
assign P3_U3196 = ~(P3_U3581 & P3_U4648); 
assign P3_U3239 = ~(P3_U4295 & P3_U3089); 
assign P3_U3261 = ~(P3_U4148 & P3_U4144 & P3_U4141 & P3_U4138); 
assign P3_U3268 = ~(P3_U3098 & P3_U7774); 
assign P3_U3272 = ~(P3_U8033 & P3_U8032); 
assign P3_U3286 = ~(P3_U7987 & P3_U7986); 
assign P3_U3364 = P3_U4340 & P3_U2630; 
assign P3_U3658 = P3_U5498 & P3_U4330; 
assign P3_U4292 = ~(HOLD & P3_U2630); 
assign P3_U4308 = ~P3_U3077; 
assign P3_U4315 = ~(P3_U4295 & P3_U2631); 
assign P3_U4328 = ~(P3_U3365 & P3_U4354); 
assign P3_U4335 = ~(P3_U4452 & P3_U3085); 
assign P3_U4345 = ~P3_U3126; 
assign P3_U4346 = ~P3_U3082; 
assign P3_U4353 = ~P3_U3124; 
assign P3_U4357 = ~(P3_U3077 & P3_ADDRESS_REG_29__SCAN_IN); 
assign P3_U4360 = ~(P3_U3077 & P3_ADDRESS_REG_28__SCAN_IN); 
assign P3_U4363 = ~(P3_U3077 & P3_ADDRESS_REG_27__SCAN_IN); 
assign P3_U4366 = ~(P3_U3077 & P3_ADDRESS_REG_26__SCAN_IN); 
assign P3_U4369 = ~(P3_U3077 & P3_ADDRESS_REG_25__SCAN_IN); 
assign P3_U4372 = ~(P3_U3077 & P3_ADDRESS_REG_24__SCAN_IN); 
assign P3_U4375 = ~(P3_U3077 & P3_ADDRESS_REG_23__SCAN_IN); 
assign P3_U4378 = ~(P3_U3077 & P3_ADDRESS_REG_22__SCAN_IN); 
assign P3_U4381 = ~(P3_U3077 & P3_ADDRESS_REG_21__SCAN_IN); 
assign P3_U4384 = ~(P3_U3077 & P3_ADDRESS_REG_20__SCAN_IN); 
assign P3_U4387 = ~(P3_U3077 & P3_ADDRESS_REG_19__SCAN_IN); 
assign P3_U4390 = ~(P3_U3077 & P3_ADDRESS_REG_18__SCAN_IN); 
assign P3_U4393 = ~(P3_U3077 & P3_ADDRESS_REG_17__SCAN_IN); 
assign P3_U4396 = ~(P3_U3077 & P3_ADDRESS_REG_16__SCAN_IN); 
assign P3_U4399 = ~(P3_U3077 & P3_ADDRESS_REG_15__SCAN_IN); 
assign P3_U4402 = ~(P3_U3077 & P3_ADDRESS_REG_14__SCAN_IN); 
assign P3_U4405 = ~(P3_U3077 & P3_ADDRESS_REG_13__SCAN_IN); 
assign P3_U4408 = ~(P3_U3077 & P3_ADDRESS_REG_12__SCAN_IN); 
assign P3_U4411 = ~(P3_U3077 & P3_ADDRESS_REG_11__SCAN_IN); 
assign P3_U4414 = ~(P3_U3077 & P3_ADDRESS_REG_10__SCAN_IN); 
assign P3_U4417 = ~(P3_U3077 & P3_ADDRESS_REG_9__SCAN_IN); 
assign P3_U4420 = ~(P3_U3077 & P3_ADDRESS_REG_8__SCAN_IN); 
assign P3_U4423 = ~(P3_U3077 & P3_ADDRESS_REG_7__SCAN_IN); 
assign P3_U4426 = ~(P3_U3077 & P3_ADDRESS_REG_6__SCAN_IN); 
assign P3_U4429 = ~(P3_U3077 & P3_ADDRESS_REG_5__SCAN_IN); 
assign P3_U4432 = ~(P3_U3077 & P3_ADDRESS_REG_4__SCAN_IN); 
assign P3_U4435 = ~(P3_U3077 & P3_ADDRESS_REG_3__SCAN_IN); 
assign P3_U4438 = ~(P3_U3077 & P3_ADDRESS_REG_2__SCAN_IN); 
assign P3_U4441 = ~(P3_U3077 & P3_ADDRESS_REG_1__SCAN_IN); 
assign P3_U4444 = ~(P3_U3077 & P3_ADDRESS_REG_0__SCAN_IN); 
assign P3_U4445 = ~P3_U3087; 
assign P3_U4449 = ~(P3_U4448 & P3_U2630); 
assign P3_U4454 = ~(HOLD & P3_U3075 & P3_U4452); 
assign P3_U4460 = ~(P3_U3087 & P3_STATE_REG_2__SCAN_IN); 
assign P3_U4466 = ~(P3_U3082 & P3_U4465); 
assign P3_U4470 = ~P3_U3098; 
assign P3_U4640 = ~P3_U3153; 
assign P3_U4666 = ~(P3_U3124 & P3_U4665 & P3_U3126); 
assign P3_U4923 = ~P3_U3169; 
assign P3_U4930 = ~(P3_U3169 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U5027 = ~P3_U3177; 
assign P3_U5033 = ~(P3_U3177 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U5332 = ~P3_U3199; 
assign P3_U5339 = ~(P3_U3199 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U5434 = ~P3_U3205; 
assign P3_U5440 = ~(P3_U3205 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U5501 = ~(P3_U5500 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_U5504 = ~P3_U3223; 
assign P3_U5505 = ~(P3_U4332 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_U5547 = ~P3_U3227; 
assign P3_U5558 = ~P3_U3228; 
assign P3_U5592 = ~(P3_U3131 & P3_U4648 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U5611 = ~P3_U3234; 
assign P3_U6403 = ~(P3_U3234 & P3_U3121); 
assign P3_U7095 = ~P3_U3257; 
assign P3_U7371 = ~(P3_U2453 & P3_U2630); 
assign P3_U7645 = ~P3_U4289; 
assign P3_U7920 = ~(P3_U3077 & P3_BE_N_REG_3__SCAN_IN); 
assign P3_U7922 = ~(P3_U3077 & P3_BE_N_REG_2__SCAN_IN); 
assign P3_U7924 = ~(P3_U3077 & P3_BE_N_REG_1__SCAN_IN); 
assign P3_U7926 = ~(P3_U3077 & P3_BE_N_REG_0__SCAN_IN); 
assign P3_U7933 = ~(P3_U3087 & P3_STATE_REG_2__SCAN_IN & P3_STATE_REG_0__SCAN_IN); 
assign P3_U7953 = ~(P3_U4628 & P3_U3121); 
assign P3_U7957 = ~(P3_U7905 & P3_STATE2_REG_0__SCAN_IN); 
assign P3_U7961 = ~(P3_U4648 & P3_U3131); 
assign P3_U8006 = ~(P3_U8005 & P3_U8004); 
assign P3_U8017 = ~(P3_U3077 & P3_W_R_N_REG_SCAN_IN); 
assign P3_U8025 = ~(P3_U3077 & P3_D_C_N_REG_SCAN_IN); 
assign P3_U8026 = ~(P3_U3077 & P3_M_IO_N_REG_SCAN_IN); 
assign P3_U8035 = ~(P3_U4289 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U2398 = P2_U4430 & P2_STATEBS16_REG_SCAN_IN; 
assign P2_U3243 = ~(P2_U3349 & P2_U3335); 
assign P2_U3312 = ~(P2_U4642 & P2_U2464); 
assign P2_U3424 = ~(P2_U2465 & P2_U4642); 
assign P2_U3462 = ~(P2_U2478 & P2_U2465); 
assign P2_U3473 = ~(P2_U2503 & P2_U4642); 
assign P2_U3530 = ~(P2_U3274 & P2_U5615); 
assign P2_U3534 = ~(P2_U4430 & P2_U3269); 
assign P2_U3547 = ~(P2_U4181 & P2_U4177 & P2_U4174 & P2_U4171); 
assign P2_U3553 = ~(P2_U4405 & P2_U3275); 
assign P2_U3582 = ~(P2_U8099 & P2_U8098); 
assign P2_U3584 = ~(P2_U8151 & P2_U8150); 
assign P2_U3682 = ~(P2_U8420 & P2_U8419); 
assign P2_U3683 = ~(P2_U8422 & P2_U8421); 
assign P2_U3711 = P2_U2360 & P2_U3266; 
assign P2_U3717 = P2_U4466 & P2_U3265; 
assign P2_U3872 = P2_U5583 & P2_U4455; 
assign P2_U4187 = P2_U3265 & P2_STATE2_REG_1__SCAN_IN; 
assign P2_U4380 = P2_U7585 & P2_U3269; 
assign P2_U4410 = ~(HOLD & P2_U3265); 
assign P2_U4439 = ~P2_U3259; 
assign P2_U4445 = ~(P2_U4430 & P2_U3302); 
assign P2_U4463 = ~(P2_U4574 & P2_U3266); 
assign P2_U4467 = ~P2_U3540; 
assign P2_U4468 = ~P2_U3304; 
assign P2_U4473 = ~P2_U3262; 
assign P2_U4474 = ~P2_U3301; 
assign P2_U4480 = ~(P2_U3259 & P2_ADDRESS_REG_29__SCAN_IN); 
assign P2_U4483 = ~(P2_U3259 & P2_ADDRESS_REG_28__SCAN_IN); 
assign P2_U4486 = ~(P2_U3259 & P2_ADDRESS_REG_27__SCAN_IN); 
assign P2_U4489 = ~(P2_U3259 & P2_ADDRESS_REG_26__SCAN_IN); 
assign P2_U4492 = ~(P2_U3259 & P2_ADDRESS_REG_25__SCAN_IN); 
assign P2_U4495 = ~(P2_U3259 & P2_ADDRESS_REG_24__SCAN_IN); 
assign P2_U4498 = ~(P2_U3259 & P2_ADDRESS_REG_23__SCAN_IN); 
assign P2_U4501 = ~(P2_U3259 & P2_ADDRESS_REG_22__SCAN_IN); 
assign P2_U4504 = ~(P2_U3259 & P2_ADDRESS_REG_21__SCAN_IN); 
assign P2_U4507 = ~(P2_U3259 & P2_ADDRESS_REG_20__SCAN_IN); 
assign P2_U4510 = ~(P2_U3259 & P2_ADDRESS_REG_19__SCAN_IN); 
assign P2_U4513 = ~(P2_U3259 & P2_ADDRESS_REG_18__SCAN_IN); 
assign P2_U4516 = ~(P2_U3259 & P2_ADDRESS_REG_17__SCAN_IN); 
assign P2_U4519 = ~(P2_U3259 & P2_ADDRESS_REG_16__SCAN_IN); 
assign P2_U4522 = ~(P2_U3259 & P2_ADDRESS_REG_15__SCAN_IN); 
assign P2_U4525 = ~(P2_U3259 & P2_ADDRESS_REG_14__SCAN_IN); 
assign P2_U4528 = ~(P2_U3259 & P2_ADDRESS_REG_13__SCAN_IN); 
assign P2_U4531 = ~(P2_U3259 & P2_ADDRESS_REG_12__SCAN_IN); 
assign P2_U4534 = ~(P2_U3259 & P2_ADDRESS_REG_11__SCAN_IN); 
assign P2_U4537 = ~(P2_U3259 & P2_ADDRESS_REG_10__SCAN_IN); 
assign P2_U4540 = ~(P2_U3259 & P2_ADDRESS_REG_9__SCAN_IN); 
assign P2_U4543 = ~(P2_U3259 & P2_ADDRESS_REG_8__SCAN_IN); 
assign P2_U4546 = ~(P2_U3259 & P2_ADDRESS_REG_7__SCAN_IN); 
assign P2_U4549 = ~(P2_U3259 & P2_ADDRESS_REG_6__SCAN_IN); 
assign P2_U4552 = ~(P2_U3259 & P2_ADDRESS_REG_5__SCAN_IN); 
assign P2_U4555 = ~(P2_U3259 & P2_ADDRESS_REG_4__SCAN_IN); 
assign P2_U4558 = ~(P2_U3259 & P2_ADDRESS_REG_3__SCAN_IN); 
assign P2_U4561 = ~(P2_U3259 & P2_ADDRESS_REG_2__SCAN_IN); 
assign P2_U4564 = ~(P2_U3259 & P2_ADDRESS_REG_1__SCAN_IN); 
assign P2_U4567 = ~(P2_U3259 & P2_ADDRESS_REG_0__SCAN_IN); 
assign P2_U4568 = ~P2_U3267; 
assign P2_U4572 = ~(P2_U4571 & P2_U3265); 
assign P2_U4575 = ~(HOLD & P2_U3256 & P2_U4574); 
assign P2_U4585 = ~(P2_U3267 & P2_STATE_REG_2__SCAN_IN); 
assign P2_U4592 = ~P2_U3274; 
assign P2_U4595 = ~(P2_U3262 & P2_U4594); 
assign P2_U4645 = ~P2_U3376; 
assign P2_U4648 = ~P2_U3349; 
assign P2_U4649 = ~P2_U3335; 
assign P2_U4827 = ~P2_U3365; 
assign P2_U4836 = ~(P2_U3365 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U5515 = ~P2_U3508; 
assign P2_U5524 = ~(P2_U3508 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U5937 = ~(P2_U5661 & P2_U3284); 
assign P2_U5940 = ~(P2_U3540 & P2_U5939); 
assign P2_U6571 = ~P2_U3545; 
assign P2_U6842 = ~(P2_U4466 & P2_U3284); 
assign P2_U7007 = ~P2_U4405; 
assign P2_U7165 = ~(P2_U4430 & P2_U3307); 
assign P2_U7582 = ~(P2_U4471 & P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P2_U7587 = ~(P2_U4471 & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P2_U7590 = ~(P2_U4471 & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P2_U7762 = ~(P2_U8005 & P2_U8004 & P2_U4593); 
assign P2_U7763 = ~(P2_U7973 & P2_U7972 & P2_U4593); 
assign P2_U7764 = ~(P2_U7957 & P2_U7956 & P2_U4593); 
assign P2_U7765 = ~(P2_U8037 & P2_U8036 & P2_U4593); 
assign P2_U7766 = ~(P2_U8021 & P2_U8020 & P2_U4593); 
assign P2_U7767 = ~(P2_U7989 & P2_U7988 & P2_U4593); 
assign P2_U7768 = ~(P2_U7941 & P2_U7940 & P2_U4593); 
assign P2_U7769 = ~(P2_U7925 & P2_U7924 & P2_U4593); 
assign P2_U7778 = ~(P2_U8007 & P2_U8006 & P2_U2456); 
assign P2_U7779 = ~(P2_U7975 & P2_U7974 & P2_U2456); 
assign P2_U7780 = ~(P2_U7959 & P2_U7958 & P2_U2456); 
assign P2_U7781 = ~(P2_U8039 & P2_U8038 & P2_U2456); 
assign P2_U7782 = ~(P2_U8023 & P2_U8022 & P2_U2456); 
assign P2_U7783 = ~(P2_U7991 & P2_U7990 & P2_U2456); 
assign P2_U7784 = ~(P2_U7943 & P2_U7942 & P2_U2456); 
assign P2_U7785 = ~(P2_U7927 & P2_U7926 & P2_U2456); 
assign P2_U7794 = ~(P2_U8009 & P2_U8008 & P2_U2454); 
assign P2_U7795 = ~(P2_U7977 & P2_U7976 & P2_U2454); 
assign P2_U7796 = ~(P2_U7961 & P2_U7960 & P2_U2454); 
assign P2_U7797 = ~(P2_U8041 & P2_U8040 & P2_U2454); 
assign P2_U7798 = ~(P2_U8025 & P2_U8024 & P2_U2454); 
assign P2_U7799 = ~(P2_U7993 & P2_U7992 & P2_U2454); 
assign P2_U7800 = ~(P2_U7945 & P2_U7944 & P2_U2454); 
assign P2_U7801 = ~(P2_U7929 & P2_U7928 & P2_U2454); 
assign P2_U7810 = ~(P2_U8011 & P2_U8010 & P2_U4590); 
assign P2_U7811 = ~(P2_U7979 & P2_U7978 & P2_U4590); 
assign P2_U7812 = ~(P2_U7963 & P2_U7962 & P2_U4590); 
assign P2_U7813 = ~(P2_U8043 & P2_U8042 & P2_U4590); 
assign P2_U7814 = ~(P2_U8027 & P2_U8026 & P2_U4590); 
assign P2_U7815 = ~(P2_U7995 & P2_U7994 & P2_U4590); 
assign P2_U7816 = ~(P2_U7947 & P2_U7946 & P2_U4590); 
assign P2_U7817 = ~(P2_U7931 & P2_U7930 & P2_U4590); 
assign P2_U7826 = ~(P2_U8013 & P2_U8012 & P2_U2453); 
assign P2_U7827 = ~(P2_U7981 & P2_U7980 & P2_U2453); 
assign P2_U7828 = ~(P2_U7965 & P2_U7964 & P2_U2453); 
assign P2_U7829 = ~(P2_U8045 & P2_U8044 & P2_U2453); 
assign P2_U7830 = ~(P2_U8029 & P2_U8028 & P2_U2453); 
assign P2_U7831 = ~(P2_U7997 & P2_U7996 & P2_U2453); 
assign P2_U7832 = ~(P2_U7949 & P2_U7948 & P2_U2453); 
assign P2_U7833 = ~(P2_U7933 & P2_U7932 & P2_U2453); 
assign P2_U7842 = ~(P2_U8015 & P2_U8014 & P2_U2452); 
assign P2_U7843 = ~(P2_U7983 & P2_U7982 & P2_U2452); 
assign P2_U7844 = ~(P2_U7967 & P2_U7966 & P2_U2452); 
assign P2_U7845 = ~(P2_U8047 & P2_U8046 & P2_U2452); 
assign P2_U7846 = ~(P2_U8031 & P2_U8030 & P2_U2452); 
assign P2_U7847 = ~(P2_U7999 & P2_U7998 & P2_U2452); 
assign P2_U7848 = ~(P2_U7951 & P2_U7950 & P2_U2452); 
assign P2_U7849 = ~(P2_U7935 & P2_U7934 & P2_U2452); 
assign P2_U7858 = ~(P2_U8017 & P2_U8016 & P2_U2455); 
assign P2_U7860 = ~(P2_U7985 & P2_U7984 & P2_U2455); 
assign P2_U7862 = ~(P2_U7969 & P2_U7968 & P2_U2455); 
assign P2_U7864 = ~(P2_U8049 & P2_U8048 & P2_U2455); 
assign P2_U7866 = ~(P2_U8033 & P2_U8032 & P2_U2455); 
assign P2_U7868 = ~(P2_U8001 & P2_U8000 & P2_U2455); 
assign P2_U7870 = ~(P2_U7953 & P2_U7952 & P2_U2455); 
assign P2_U7872 = ~(P2_U7937 & P2_U7936 & P2_U2455); 
assign P2_U7899 = ~(P2_U3259 & P2_BE_N_REG_3__SCAN_IN); 
assign P2_U7901 = ~(P2_U3259 & P2_BE_N_REG_2__SCAN_IN); 
assign P2_U7903 = ~(P2_U3259 & P2_BE_N_REG_1__SCAN_IN); 
assign P2_U7905 = ~(P2_U3259 & P2_BE_N_REG_0__SCAN_IN); 
assign P2_U7907 = ~(P2_U3268 & P2_U3267 & P2_STATE_REG_0__SCAN_IN); 
assign P2_U7913 = ~(P2_U3267 & P2_STATE_REG_2__SCAN_IN & P2_STATE_REG_0__SCAN_IN); 
assign P2_U8066 = ~(P2_U4642 & P2_U3310); 
assign P2_U8078 = ~(P2_U5585 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8081 = ~(P2_U4590 & P2_U3273); 
assign P2_U8130 = ~(P2_U3259 & P2_W_R_N_REG_SCAN_IN); 
assign P2_U8140 = ~(P2_U3259 & P2_D_C_N_REG_SCAN_IN); 
assign P2_U8141 = ~(P2_U3259 & P2_M_IO_N_REG_SCAN_IN); 
assign P2_U8147 = ~(P2_U4405 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8424 = ~(P2_U2615 & P2_STATE2_REG_1__SCAN_IN); 
assign P2_U8426 = ~(P2_U2615 & P2_STATE2_REG_1__SCAN_IN); 
assign P1_U2388 = P1_U4209 & P1_STATEBS16_REG_SCAN_IN; 
assign P1_U2458 = P1_U3507 & P1_U4378; 
assign P1_U2464 = P1_U4380 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P1_U2467 = P1_U3270 & P1_U4378 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P1_U2472 = P1_U4380 & P1_U3270; 
assign P1_U2521 = P1_U3402 & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_U2524 = P1_U3266 & P1_U3402; 
assign P1_U2607 = P1_U7672 & P1_U7671; 
assign P1_U3235 = ~(P1_U3329 & P1_U3323); 
assign P1_U3259 = ~(P1_U3260 & P1_STATE_REG_0__SCAN_IN); 
assign P1_U3306 = ~(P1_U4533 & P1_U2478); 
assign P1_U3320 = ~(P1_U4209 & P1_U3308); 
assign P1_U3356 = ~(P1_U2479 & P1_U4533); 
assign P1_U3370 = ~(P1_U2488 & P1_U2479); 
assign P1_U3373 = ~(P1_U2510 & P1_U4533); 
assign P1_U3401 = ~(P1_U3444 & P1_U5510); 
assign P1_U3432 = ~(P1_U4209 & P1_U3262); 
assign P1_U3433 = ~(P1_U3962 & P1_U3958 & P1_U3955 & P1_U3952); 
assign P1_U3445 = ~(P1_U3274 & P1_U7064); 
assign P1_U3452 = ~(P1_U4183 & P1_U3268); 
assign P1_U3456 = ~(P1_U7719 & P1_U7718); 
assign P1_U3471 = ~(P1_U7714 & P1_U7713); 
assign P1_U3533 = P1_U4414 & P1_U4413; 
assign P1_U3539 = P1_U7678 & P1_U7677 & P1_U7676 & P1_U7675; 
assign P1_U3554 = P1_U7658 & P1_U7657 & P1_U7656 & P1_U7655; 
assign P1_U3555 = P1_U7662 & P1_U7661 & P1_U7660 & P1_U7659; 
assign P1_U3556 = P1_U7666 & P1_U7665 & P1_U7664 & P1_U7663; 
assign P1_U3557 = P1_U7670 & P1_U7669 & P1_U7668 & P1_U7667; 
assign P1_U3576 = P1_U4414 & P1_U4413; 
assign P1_U3583 = P1_U2427 & P1_U3257; 
assign P1_U3739 = P1_U5475 & P1_U4242; 
assign P1_U3964 = P1_U3257 & P1_STATE2_REG_2__SCAN_IN; 
assign P1_U4071 = P1_U4414 & P1_U4413; 
assign P1_U4170 = P1_U7674 & P1_U7673; 
assign P1_U4185 = ~(HOLD & P1_U3257); 
assign P1_U4187 = ~P1_U3440; 
assign P1_U4203 = ~P1_U3408; 
assign P1_U4221 = ~P1_U3249; 
assign P1_U4235 = ~P1_U3297; 
assign P1_U4241 = ~(P1_U3584 & P1_U4261); 
assign P1_U4243 = ~(P1_U4364 & P1_U3258); 
assign P1_U4258 = ~P1_U3254; 
assign P1_U4269 = ~(P1_U3249 & P1_ADDRESS_REG_29__SCAN_IN); 
assign P1_U4272 = ~(P1_U3249 & P1_ADDRESS_REG_28__SCAN_IN); 
assign P1_U4275 = ~(P1_U3249 & P1_ADDRESS_REG_27__SCAN_IN); 
assign P1_U4278 = ~(P1_U3249 & P1_ADDRESS_REG_26__SCAN_IN); 
assign P1_U4281 = ~(P1_U3249 & P1_ADDRESS_REG_25__SCAN_IN); 
assign P1_U4284 = ~(P1_U3249 & P1_ADDRESS_REG_24__SCAN_IN); 
assign P1_U4287 = ~(P1_U3249 & P1_ADDRESS_REG_23__SCAN_IN); 
assign P1_U4290 = ~(P1_U3249 & P1_ADDRESS_REG_22__SCAN_IN); 
assign P1_U4293 = ~(P1_U3249 & P1_ADDRESS_REG_21__SCAN_IN); 
assign P1_U4296 = ~(P1_U3249 & P1_ADDRESS_REG_20__SCAN_IN); 
assign P1_U4299 = ~(P1_U3249 & P1_ADDRESS_REG_19__SCAN_IN); 
assign P1_U4302 = ~(P1_U3249 & P1_ADDRESS_REG_18__SCAN_IN); 
assign P1_U4305 = ~(P1_U3249 & P1_ADDRESS_REG_17__SCAN_IN); 
assign P1_U4308 = ~(P1_U3249 & P1_ADDRESS_REG_16__SCAN_IN); 
assign P1_U4311 = ~(P1_U3249 & P1_ADDRESS_REG_15__SCAN_IN); 
assign P1_U4314 = ~(P1_U3249 & P1_ADDRESS_REG_14__SCAN_IN); 
assign P1_U4317 = ~(P1_U3249 & P1_ADDRESS_REG_13__SCAN_IN); 
assign P1_U4320 = ~(P1_U3249 & P1_ADDRESS_REG_12__SCAN_IN); 
assign P1_U4323 = ~(P1_U3249 & P1_ADDRESS_REG_11__SCAN_IN); 
assign P1_U4326 = ~(P1_U3249 & P1_ADDRESS_REG_10__SCAN_IN); 
assign P1_U4329 = ~(P1_U3249 & P1_ADDRESS_REG_9__SCAN_IN); 
assign P1_U4332 = ~(P1_U3249 & P1_ADDRESS_REG_8__SCAN_IN); 
assign P1_U4335 = ~(P1_U3249 & P1_ADDRESS_REG_7__SCAN_IN); 
assign P1_U4338 = ~(P1_U3249 & P1_ADDRESS_REG_6__SCAN_IN); 
assign P1_U4341 = ~(P1_U3249 & P1_ADDRESS_REG_5__SCAN_IN); 
assign P1_U4344 = ~(P1_U3249 & P1_ADDRESS_REG_4__SCAN_IN); 
assign P1_U4347 = ~(P1_U3249 & P1_ADDRESS_REG_3__SCAN_IN); 
assign P1_U4350 = ~(P1_U3249 & P1_ADDRESS_REG_2__SCAN_IN); 
assign P1_U4353 = ~(P1_U3249 & P1_ADDRESS_REG_1__SCAN_IN); 
assign P1_U4356 = ~(P1_U3249 & P1_ADDRESS_REG_0__SCAN_IN); 
assign P1_U4357 = ~P1_U3260; 
assign P1_U4361 = ~(P1_U4360 & P1_U3257); 
assign P1_U4365 = ~(HOLD & P1_U3247 & P1_U4364); 
assign P1_U4372 = ~(P1_U3260 & P1_STATE_REG_2__SCAN_IN); 
assign P1_U4377 = ~P1_U3280; 
assign P1_U4379 = ~P1_U3444; 
assign P1_U4381 = ~P1_U3274; 
assign P1_U4382 = ~P1_U3267; 
assign P1_U4385 = ~(P1_U2471 & P1_INSTQUEUE_REG_1__3__SCAN_IN); 
assign P1_U4386 = ~(P1_U2470 & P1_INSTQUEUE_REG_2__3__SCAN_IN); 
assign P1_U4387 = ~(P1_U2468 & P1_INSTQUEUE_REG_3__3__SCAN_IN); 
assign P1_U4389 = ~(P1_U2466 & P1_INSTQUEUE_REG_5__3__SCAN_IN); 
assign P1_U4390 = ~(P1_U2465 & P1_INSTQUEUE_REG_6__3__SCAN_IN); 
assign P1_U4392 = ~(P1_U2463 & P1_INSTQUEUE_REG_9__3__SCAN_IN); 
assign P1_U4393 = ~(P1_U2461 & P1_INSTQUEUE_REG_10__3__SCAN_IN); 
assign P1_U4394 = ~(P1_U2459 & P1_INSTQUEUE_REG_11__3__SCAN_IN); 
assign P1_U4396 = ~(P1_U2457 & P1_INSTQUEUE_REG_13__3__SCAN_IN); 
assign P1_U4397 = ~(P1_U2455 & P1_INSTQUEUE_REG_14__3__SCAN_IN); 
assign P1_U4402 = ~(P1_U3270 & P1_U4380 & P1_INSTQUEUE_REG_0__5__SCAN_IN); 
assign P1_U4405 = ~(P1_U4378 & P1_U3270 & P1_INSTQUEUE_REG_4__5__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_U4408 = ~(P1_U3524 & P1_U4380); 
assign P1_U4411 = ~(P1_U4378 & P1_U3527 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_U4418 = ~(P1_U2471 & P1_INSTQUEUE_REG_1__2__SCAN_IN); 
assign P1_U4419 = ~(P1_U2470 & P1_INSTQUEUE_REG_2__2__SCAN_IN); 
assign P1_U4420 = ~(P1_U2468 & P1_INSTQUEUE_REG_3__2__SCAN_IN); 
assign P1_U4422 = ~(P1_U2466 & P1_INSTQUEUE_REG_5__2__SCAN_IN); 
assign P1_U4423 = ~(P1_U2465 & P1_INSTQUEUE_REG_6__2__SCAN_IN); 
assign P1_U4425 = ~(P1_U2463 & P1_INSTQUEUE_REG_9__2__SCAN_IN); 
assign P1_U4426 = ~(P1_U2461 & P1_INSTQUEUE_REG_10__2__SCAN_IN); 
assign P1_U4427 = ~(P1_U2459 & P1_INSTQUEUE_REG_11__2__SCAN_IN); 
assign P1_U4429 = ~(P1_U2457 & P1_INSTQUEUE_REG_13__2__SCAN_IN); 
assign P1_U4430 = ~(P1_U2455 & P1_INSTQUEUE_REG_14__2__SCAN_IN); 
assign P1_U4435 = ~(P1_U2471 & P1_INSTQUEUE_REG_1__7__SCAN_IN); 
assign P1_U4436 = ~(P1_U2470 & P1_INSTQUEUE_REG_2__7__SCAN_IN); 
assign P1_U4437 = ~(P1_U2468 & P1_INSTQUEUE_REG_3__7__SCAN_IN); 
assign P1_U4439 = ~(P1_U2466 & P1_INSTQUEUE_REG_5__7__SCAN_IN); 
assign P1_U4440 = ~(P1_U2465 & P1_INSTQUEUE_REG_6__7__SCAN_IN); 
assign P1_U4442 = ~(P1_U2463 & P1_INSTQUEUE_REG_9__7__SCAN_IN); 
assign P1_U4443 = ~(P1_U2461 & P1_INSTQUEUE_REG_10__7__SCAN_IN); 
assign P1_U4444 = ~(P1_U2459 & P1_INSTQUEUE_REG_11__7__SCAN_IN); 
assign P1_U4446 = ~(P1_U2457 & P1_INSTQUEUE_REG_13__7__SCAN_IN); 
assign P1_U4447 = ~(P1_U2455 & P1_INSTQUEUE_REG_14__7__SCAN_IN); 
assign P1_U4451 = ~(P1_U2469 & P1_U2456 & P1_INSTQUEUE_REG_1__6__SCAN_IN); 
assign P1_U4452 = ~(P1_U2469 & P1_U2454 & P1_INSTQUEUE_REG_2__6__SCAN_IN); 
assign P1_U4456 = ~(P1_U4378 & P1_U3507 & P1_INSTQUEUE_REG_12__6__SCAN_IN); 
assign P1_U4457 = ~(P1_U3507 & P1_U2456 & P1_INSTQUEUE_REG_13__6__SCAN_IN); 
assign P1_U4458 = ~(P1_U3507 & P1_U2454 & P1_INSTQUEUE_REG_14__6__SCAN_IN); 
assign P1_U4463 = ~(P1_U2471 & P1_INSTQUEUE_REG_1__1__SCAN_IN); 
assign P1_U4464 = ~(P1_U2470 & P1_INSTQUEUE_REG_2__1__SCAN_IN); 
assign P1_U4465 = ~(P1_U2468 & P1_INSTQUEUE_REG_3__1__SCAN_IN); 
assign P1_U4467 = ~(P1_U2466 & P1_INSTQUEUE_REG_5__1__SCAN_IN); 
assign P1_U4468 = ~(P1_U2465 & P1_INSTQUEUE_REG_6__1__SCAN_IN); 
assign P1_U4470 = ~(P1_U2463 & P1_INSTQUEUE_REG_9__1__SCAN_IN); 
assign P1_U4471 = ~(P1_U2461 & P1_INSTQUEUE_REG_10__1__SCAN_IN); 
assign P1_U4472 = ~(P1_U2459 & P1_INSTQUEUE_REG_11__1__SCAN_IN); 
assign P1_U4474 = ~(P1_U2457 & P1_INSTQUEUE_REG_13__1__SCAN_IN); 
assign P1_U4475 = ~(P1_U2455 & P1_INSTQUEUE_REG_14__1__SCAN_IN); 
assign P1_U4480 = ~(P1_U2471 & P1_INSTQUEUE_REG_1__0__SCAN_IN); 
assign P1_U4481 = ~(P1_U2470 & P1_INSTQUEUE_REG_2__0__SCAN_IN); 
assign P1_U4482 = ~(P1_U2468 & P1_INSTQUEUE_REG_3__0__SCAN_IN); 
assign P1_U4484 = ~(P1_U2466 & P1_INSTQUEUE_REG_5__0__SCAN_IN); 
assign P1_U4485 = ~(P1_U2465 & P1_INSTQUEUE_REG_6__0__SCAN_IN); 
assign P1_U4487 = ~(P1_U2463 & P1_INSTQUEUE_REG_9__0__SCAN_IN); 
assign P1_U4488 = ~(P1_U2461 & P1_INSTQUEUE_REG_10__0__SCAN_IN); 
assign P1_U4489 = ~(P1_U2459 & P1_INSTQUEUE_REG_11__0__SCAN_IN); 
assign P1_U4491 = ~(P1_U2457 & P1_INSTQUEUE_REG_13__0__SCAN_IN); 
assign P1_U4492 = ~(P1_U2455 & P1_INSTQUEUE_REG_14__0__SCAN_IN); 
assign P1_U4496 = ~(P1_U3254 & P1_U4495); 
assign P1_U4538 = ~P1_U3340; 
assign P1_U4541 = ~P1_U3329; 
assign P1_U4542 = ~P1_U3323; 
assign P1_U4718 = ~P1_U3337; 
assign P1_U4726 = ~(P1_U3337 & P1_STATE2_REG_3__SCAN_IN); 
assign P1_U5406 = ~P1_U3384; 
assign P1_U5414 = ~(P1_U3384 & P1_STATE2_REG_3__SCAN_IN); 
assign P1_U5482 = ~(P1_U5481 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P1_U5485 = ~(P1_U5484 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P1_U5519 = ~P1_U3402; 
assign P1_U5794 = ~(P1_U4209 & P1_U3294); 
assign P1_U5798 = ~(P1_U5797 & P1_U5796); 
assign P1_U6602 = ~(P1_U3966 & P1_U2428); 
assign P1_U7095 = ~(P1_U3297 & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P1_U7215 = ~(P1_U3297 & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P1_U7217 = ~(P1_U3297 & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P1_U7219 = ~P1_U4183; 
assign P1_U7457 = ~(P1_U2430 & P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P1_U7459 = ~(P1_U2430 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P1_U7462 = ~(P1_U2430 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_U7465 = ~(P1_U2430 & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U7467 = ~(P1_U2430 & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U7633 = ~(P1_U3249 & P1_BE_N_REG_3__SCAN_IN); 
assign P1_U7635 = ~(P1_U3249 & P1_BE_N_REG_2__SCAN_IN); 
assign P1_U7637 = ~(P1_U3249 & P1_BE_N_REG_1__SCAN_IN); 
assign P1_U7639 = ~(P1_U3249 & P1_BE_N_REG_0__SCAN_IN); 
assign P1_U7646 = ~(P1_U3260 & P1_STATE_REG_2__SCAN_IN & P1_STATE_REG_0__SCAN_IN); 
assign P1_U7684 = ~(P1_U4513 & P1_U3294); 
assign P1_U7688 = ~(P1_U7469 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U7695 = ~(P1_U4533 & P1_U3304); 
assign P1_U7750 = ~(P1_U7749 & P1_U7748); 
assign P1_U7761 = ~(P1_U3249 & P1_W_R_N_REG_SCAN_IN); 
assign P1_U7769 = ~(P1_U3249 & P1_D_C_N_REG_SCAN_IN); 
assign P1_U7770 = ~(P1_U3249 & P1_M_IO_N_REG_SCAN_IN); 
assign P1_U7787 = ~(P1_U3297 & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P1_U7788 = ~(P1_U4183 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign R170_U15 = ~(R170_U14 & R170_U12 & R170_U10 & R170_U8); 
assign R165_U15 = ~(R165_U14 & R165_U12 & R165_U10 & R165_U8); 
assign P3_ADD_526_U13 = ~(P3_ADD_526_U82 & P3_ADD_526_U111); 
assign P3_ADD_526_U71 = ~(P3_ADD_526_U182 & P3_ADD_526_U181); 
assign P3_ADD_526_U97 = ~(P3_ADD_526_U111 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_526_U153 = ~(P3_ADD_526_U111 & P3_ADD_526_U9); 
assign P3_ADD_526_U160 = ~(P3_ADD_526_U130 & P3_ADD_526_U6); 
assign P3_ADD_552_U13 = ~(P3_ADD_552_U82 & P3_ADD_552_U111); 
assign P3_ADD_552_U71 = ~(P3_ADD_552_U182 & P3_ADD_552_U181); 
assign P3_ADD_552_U97 = ~(P3_ADD_552_U111 & P3_EBX_REG_3__SCAN_IN); 
assign P3_ADD_552_U153 = ~(P3_ADD_552_U111 & P3_ADD_552_U9); 
assign P3_ADD_552_U160 = ~(P3_ADD_552_U130 & P3_ADD_552_U6); 
assign P3_ADD_546_U13 = ~(P3_ADD_546_U82 & P3_ADD_546_U111); 
assign P3_ADD_546_U71 = ~(P3_ADD_546_U182 & P3_ADD_546_U181); 
assign P3_ADD_546_U97 = ~(P3_ADD_546_U111 & P3_EAX_REG_3__SCAN_IN); 
assign P3_ADD_546_U153 = ~(P3_ADD_546_U111 & P3_ADD_546_U9); 
assign P3_ADD_546_U160 = ~(P3_ADD_546_U130 & P3_ADD_546_U6); 
assign P3_ADD_476_U8 = ~(P3_ADD_476_U94 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_476_U71 = ~(P3_ADD_476_U142 & P3_ADD_476_U141); 
assign P3_ADD_476_U136 = ~(P3_ADD_476_U94 & P3_ADD_476_U7); 
assign P3_ADD_531_U9 = ~(P3_ADD_531_U98 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_531_U85 = ~(P3_ADD_531_U169 & P3_ADD_531_U168); 
assign P3_ADD_531_U147 = ~(P3_ADD_531_U98 & P3_ADD_531_U8); 
assign P3_SUB_320_U149 = ~(P3_SUB_320_U71 & P3_PHYADDRPOINTER_REG_0__SCAN_IN); 
assign P3_ADD_505_U10 = ~(P3_ADD_505_U18 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_ADD_505_U17 = ~(P3_ADD_505_U28 & P3_ADD_505_U27); 
assign P3_ADD_505_U26 = ~(P3_ADD_505_U18 & P3_ADD_505_U9); 
assign P3_ADD_318_U8 = ~(P3_ADD_318_U94 & P3_PHYADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_318_U71 = ~(P3_ADD_318_U142 & P3_ADD_318_U141); 
assign P3_ADD_318_U136 = ~(P3_ADD_318_U94 & P3_ADD_318_U7); 
assign P3_SUB_370_U7 = ~(P3_SUB_370_U9 & P3_SUB_370_U46); 
assign P3_SUB_370_U23 = ~(P3_SUB_370_U48 & P3_SUB_370_U47); 
assign P3_SUB_370_U24 = ~(P3_SUB_370_U53 & P3_SUB_370_U52); 
assign P3_SUB_370_U25 = ~(P3_SUB_370_U58 & P3_SUB_370_U57); 
assign P3_SUB_370_U26 = ~(P3_SUB_370_U63 & P3_SUB_370_U62); 
assign P3_SUB_370_U30 = ~P3_SUB_370_U9; 
assign P3_SUB_370_U33 = ~(P3_SUB_370_U9 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_ADD_315_U8 = ~(P3_ADD_315_U91 & P3_PHYADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_315_U66 = ~(P3_ADD_315_U132 & P3_ADD_315_U131); 
assign P3_ADD_315_U130 = ~(P3_ADD_315_U91 & P3_ADD_315_U7); 
assign P3_SUB_589_U8 = ~P3_U2632; 
assign P3_ADD_467_U8 = ~(P3_ADD_467_U94 & P3_REIP_REG_3__SCAN_IN); 
assign P3_ADD_467_U71 = ~(P3_ADD_467_U142 & P3_ADD_467_U141); 
assign P3_ADD_467_U136 = ~(P3_ADD_467_U94 & P3_ADD_467_U7); 
assign P3_ADD_430_U8 = ~(P3_ADD_430_U94 & P3_REIP_REG_3__SCAN_IN); 
assign P3_ADD_430_U71 = ~(P3_ADD_430_U142 & P3_ADD_430_U141); 
assign P3_ADD_430_U136 = ~(P3_ADD_430_U94 & P3_ADD_430_U7); 
assign P3_ADD_380_U9 = ~(P3_ADD_380_U98 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_380_U85 = ~(P3_ADD_380_U169 & P3_ADD_380_U168); 
assign P3_ADD_380_U147 = ~(P3_ADD_380_U98 & P3_ADD_380_U8); 
assign P3_ADD_344_U9 = ~(P3_ADD_344_U98 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_344_U85 = ~(P3_ADD_344_U169 & P3_ADD_344_U168); 
assign P3_ADD_344_U147 = ~(P3_ADD_344_U98 & P3_ADD_344_U8); 
assign P3_ADD_339_U8 = ~(P3_ADD_339_U94 & P3_PHYADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_339_U71 = ~(P3_ADD_339_U142 & P3_ADD_339_U141); 
assign P3_ADD_339_U136 = ~(P3_ADD_339_U94 & P3_ADD_339_U7); 
assign P3_SUB_580_U6 = ~(P3_SUB_580_U10 & P3_SUB_580_U9); 
assign P3_ADD_541_U8 = ~(P3_ADD_541_U94 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_541_U71 = ~(P3_ADD_541_U142 & P3_ADD_541_U141); 
assign P3_ADD_541_U136 = ~(P3_ADD_541_U94 & P3_ADD_541_U7); 
assign P3_SUB_355_U7 = ~(P3_SUB_355_U9 & P3_SUB_355_U46); 
assign P3_SUB_355_U23 = ~(P3_SUB_355_U48 & P3_SUB_355_U47); 
assign P3_SUB_355_U24 = ~(P3_SUB_355_U53 & P3_SUB_355_U52); 
assign P3_SUB_355_U25 = ~(P3_SUB_355_U58 & P3_SUB_355_U57); 
assign P3_SUB_355_U26 = ~(P3_SUB_355_U63 & P3_SUB_355_U62); 
assign P3_SUB_355_U30 = ~P3_SUB_355_U9; 
assign P3_SUB_355_U33 = ~(P3_SUB_355_U9 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_SUB_450_U20 = ~(P3_SUB_450_U45 & P3_SUB_450_U44); 
assign P3_SUB_450_U21 = ~(P3_SUB_450_U50 & P3_SUB_450_U49); 
assign P3_SUB_450_U22 = ~(P3_SUB_450_U55 & P3_SUB_450_U54); 
assign P3_SUB_450_U23 = ~(P3_SUB_450_U60 & P3_SUB_450_U59); 
assign P3_SUB_450_U28 = ~P3_SUB_450_U7; 
assign P3_SUB_450_U31 = ~(P3_SUB_450_U7 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_SUB_357_1258_U208 = ~(P3_SUB_357_1258_U207 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_486_U10 = ~(P3_ADD_486_U18 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_ADD_486_U17 = ~(P3_ADD_486_U28 & P3_ADD_486_U27); 
assign P3_ADD_486_U26 = ~(P3_ADD_486_U18 & P3_ADD_486_U9); 
assign P3_SUB_485_U20 = ~(P3_SUB_485_U45 & P3_SUB_485_U44); 
assign P3_SUB_485_U21 = ~(P3_SUB_485_U50 & P3_SUB_485_U49); 
assign P3_SUB_485_U22 = ~(P3_SUB_485_U55 & P3_SUB_485_U54); 
assign P3_SUB_485_U23 = ~(P3_SUB_485_U60 & P3_SUB_485_U59); 
assign P3_SUB_485_U28 = ~P3_SUB_485_U7; 
assign P3_SUB_485_U31 = ~(P3_SUB_485_U7 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_ADD_515_U8 = ~(P3_ADD_515_U94 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_515_U71 = ~(P3_ADD_515_U142 & P3_ADD_515_U141); 
assign P3_ADD_515_U136 = ~(P3_ADD_515_U94 & P3_ADD_515_U7); 
assign P3_ADD_394_U5 = ~(P3_ADD_394_U92 & P3_ADD_394_U126); 
assign P3_ADD_394_U8 = ~(P3_ADD_394_U92 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_394_U81 = ~(P3_ADD_394_U166 & P3_ADD_394_U165); 
assign P3_ADD_394_U97 = ~P3_ADD_394_U92; 
assign P3_ADD_394_U139 = ~(P3_ADD_394_U92 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_SUB_414_U17 = P3_SUB_414_U105 & P3_SUB_414_U21; 
assign P3_SUB_414_U22 = ~(P3_SUB_414_U27 & P3_SUB_414_U58 & P3_SUB_414_U83); 
assign P3_SUB_414_U50 = ~(P3_SUB_414_U149 & P3_SUB_414_U148); 
assign P3_SUB_414_U91 = ~(P3_SUB_414_U83 & P3_SUB_414_U58); 
assign P3_SUB_414_U135 = ~(P3_SUB_414_U83 & P3_SUB_414_U58); 
assign P3_ADD_441_U8 = ~(P3_ADD_441_U94 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_441_U71 = ~(P3_ADD_441_U142 & P3_ADD_441_U141); 
assign P3_ADD_441_U136 = ~(P3_ADD_441_U94 & P3_ADD_441_U7); 
assign P3_ADD_349_U9 = ~(P3_ADD_349_U98 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_349_U85 = ~(P3_ADD_349_U169 & P3_ADD_349_U168); 
assign P3_ADD_349_U147 = ~(P3_ADD_349_U98 & P3_ADD_349_U8); 
assign P3_ADD_405_U5 = ~(P3_ADD_405_U92 & P3_ADD_405_U126); 
assign P3_ADD_405_U8 = ~(P3_ADD_405_U92 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_405_U81 = ~(P3_ADD_405_U166 & P3_ADD_405_U165); 
assign P3_ADD_405_U97 = ~P3_ADD_405_U92; 
assign P3_ADD_405_U139 = ~(P3_ADD_405_U92 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_553_U9 = ~(P3_ADD_553_U98 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_553_U85 = ~(P3_ADD_553_U169 & P3_ADD_553_U168); 
assign P3_ADD_553_U147 = ~(P3_ADD_553_U98 & P3_ADD_553_U8); 
assign P3_ADD_558_U9 = ~(P3_ADD_558_U98 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_558_U85 = ~(P3_ADD_558_U169 & P3_ADD_558_U168); 
assign P3_ADD_558_U147 = ~(P3_ADD_558_U98 & P3_ADD_558_U8); 
assign P3_ADD_385_U9 = ~(P3_ADD_385_U98 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_385_U85 = ~(P3_ADD_385_U169 & P3_ADD_385_U168); 
assign P3_ADD_385_U147 = ~(P3_ADD_385_U98 & P3_ADD_385_U8); 
assign P3_ADD_547_U9 = ~(P3_ADD_547_U98 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_547_U85 = ~(P3_ADD_547_U169 & P3_ADD_547_U168); 
assign P3_ADD_547_U147 = ~(P3_ADD_547_U98 & P3_ADD_547_U8); 
assign P3_SUB_412_U20 = ~(P3_SUB_412_U45 & P3_SUB_412_U44); 
assign P3_SUB_412_U21 = ~(P3_SUB_412_U50 & P3_SUB_412_U49); 
assign P3_SUB_412_U22 = ~(P3_SUB_412_U55 & P3_SUB_412_U54); 
assign P3_SUB_412_U23 = ~(P3_SUB_412_U60 & P3_SUB_412_U59); 
assign P3_SUB_412_U28 = ~P3_SUB_412_U7; 
assign P3_SUB_412_U31 = ~(P3_SUB_412_U7 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_SUB_504_U20 = ~(P3_SUB_504_U45 & P3_SUB_504_U44); 
assign P3_SUB_504_U21 = ~(P3_SUB_504_U50 & P3_SUB_504_U49); 
assign P3_SUB_504_U22 = ~(P3_SUB_504_U55 & P3_SUB_504_U54); 
assign P3_SUB_504_U23 = ~(P3_SUB_504_U60 & P3_SUB_504_U59); 
assign P3_SUB_504_U28 = ~P3_SUB_504_U7; 
assign P3_SUB_504_U31 = ~(P3_SUB_504_U7 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_SUB_401_U7 = ~(P3_SUB_401_U9 & P3_SUB_401_U46); 
assign P3_SUB_401_U23 = ~(P3_SUB_401_U48 & P3_SUB_401_U47); 
assign P3_SUB_401_U24 = ~(P3_SUB_401_U53 & P3_SUB_401_U52); 
assign P3_SUB_401_U25 = ~(P3_SUB_401_U58 & P3_SUB_401_U57); 
assign P3_SUB_401_U26 = ~(P3_SUB_401_U63 & P3_SUB_401_U62); 
assign P3_SUB_401_U30 = ~P3_SUB_401_U9; 
assign P3_SUB_401_U33 = ~(P3_SUB_401_U9 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_SUB_390_U7 = ~(P3_SUB_390_U9 & P3_SUB_390_U46); 
assign P3_SUB_390_U23 = ~(P3_SUB_390_U48 & P3_SUB_390_U47); 
assign P3_SUB_390_U24 = ~(P3_SUB_390_U53 & P3_SUB_390_U52); 
assign P3_SUB_390_U25 = ~(P3_SUB_390_U58 & P3_SUB_390_U57); 
assign P3_SUB_390_U26 = ~(P3_SUB_390_U63 & P3_SUB_390_U62); 
assign P3_SUB_390_U30 = ~P3_SUB_390_U9; 
assign P3_SUB_390_U33 = ~(P3_SUB_390_U9 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_ADD_495_U10 = ~(P3_ADD_495_U20 & P3_ADD_495_U19); 
assign P3_ADD_495_U12 = ~(P3_ADD_495_U13 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_ADD_495_U18 = ~(P3_ADD_495_U13 & P3_ADD_495_U7); 
assign P3_ADD_494_U8 = ~(P3_ADD_494_U94 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_494_U71 = ~(P3_ADD_494_U142 & P3_ADD_494_U141); 
assign P3_ADD_494_U136 = ~(P3_ADD_494_U94 & P3_ADD_494_U7); 
assign P3_ADD_536_U8 = ~(P3_ADD_536_U94 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_536_U71 = ~(P3_ADD_536_U142 & P3_ADD_536_U141); 
assign P3_ADD_536_U136 = ~(P3_ADD_536_U94 & P3_ADD_536_U7); 
assign P2_R2027_U9 = ~(P2_R2027_U98 & P2_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P2_R2027_U85 = ~(P2_R2027_U169 & P2_R2027_U168); 
assign P2_R2027_U147 = ~(P2_R2027_U98 & P2_R2027_U8); 
assign P2_R2337_U9 = ~(P2_R2337_U95 & P2_PHYADDRPOINTER_REG_4__SCAN_IN); 
assign P2_R2337_U70 = ~(P2_R2337_U142 & P2_R2337_U141); 
assign P2_R2337_U134 = ~(P2_R2337_U95 & P2_R2337_U8); 
assign P2_R2337_U136 = ~(P2_R2337_U94 & P2_R2337_U5); 
assign P2_R2147_U9 = ~(P2_R2147_U20 & P2_R2147_U19); 
assign P2_R2147_U18 = ~(P2_R2147_U14 & P2_R2147_U5); 
assign P2_SUB_589_U8 = ~P2_U2813; 
assign P2_R2238_U7 = ~(P2_R2238_U9 & P2_R2238_U46); 
assign P2_R2238_U23 = ~(P2_R2238_U48 & P2_R2238_U47); 
assign P2_R2238_U24 = ~(P2_R2238_U53 & P2_R2238_U52); 
assign P2_R2238_U25 = ~(P2_R2238_U58 & P2_R2238_U57); 
assign P2_R2238_U26 = ~(P2_R2238_U63 & P2_R2238_U62); 
assign P2_R2238_U30 = ~P2_R2238_U9; 
assign P2_R2238_U33 = ~(P2_R2238_U9 & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P2_SUB_450_U21 = ~(P2_SUB_450_U45 & P2_SUB_450_U44); 
assign P2_SUB_450_U22 = ~(P2_SUB_450_U50 & P2_SUB_450_U49); 
assign P2_SUB_450_U23 = ~(P2_SUB_450_U55 & P2_SUB_450_U54); 
assign P2_SUB_450_U24 = ~(P2_SUB_450_U60 & P2_SUB_450_U59); 
assign P2_SUB_450_U28 = ~P2_SUB_450_U7; 
assign P2_SUB_450_U31 = ~(P2_SUB_450_U7 & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P2_ADD_394_U5 = ~(P2_ADD_394_U94 & P2_ADD_394_U125); 
assign P2_ADD_394_U8 = ~(P2_ADD_394_U94 & P2_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P2_ADD_394_U85 = ~(P2_ADD_394_U174 & P2_ADD_394_U173); 
assign P2_ADD_394_U97 = ~P2_ADD_394_U94; 
assign P2_ADD_394_U171 = ~(P2_ADD_394_U94 & P2_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P2_ADD_371_1212_U11 = P2_ADD_371_1212_U7 & P2_ADD_371_1212_U88; 
assign P2_ADD_371_1212_U95 = P2_ADD_371_1212_U7 & P2_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P2_ADD_371_1212_U100 = P2_ADD_371_1212_U7 & P2_ADD_371_1212_U101; 
assign P2_ADD_371_1212_U105 = P2_ADD_371_1212_U4 & P2_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P1_R2027_U13 = ~(P1_R2027_U82 & P1_R2027_U111); 
assign P1_R2027_U71 = ~(P1_R2027_U182 & P1_R2027_U181); 
assign P1_R2027_U97 = ~(P1_R2027_U111 & P1_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P1_R2027_U153 = ~(P1_R2027_U111 & P1_R2027_U9); 
assign P1_R2027_U160 = ~(P1_R2027_U130 & P1_R2027_U6); 
assign P1_R2337_U8 = ~(P1_R2337_U94 & P1_PHYADDRPOINTER_REG_3__SCAN_IN); 
assign P1_R2337_U71 = ~(P1_R2337_U142 & P1_R2337_U141); 
assign P1_R2337_U136 = ~(P1_R2337_U94 & P1_R2337_U7); 
assign P1_SUB_580_U6 = ~(P1_SUB_580_U10 & P1_SUB_580_U9); 
assign P1_R2096_U8 = ~(P1_R2096_U94 & P1_REIP_REG_3__SCAN_IN); 
assign P1_R2096_U71 = ~(P1_R2096_U142 & P1_R2096_U141); 
assign P1_R2096_U136 = ~(P1_R2096_U94 & P1_R2096_U7); 
assign P1_R2238_U7 = ~(P1_R2238_U9 & P1_R2238_U46); 
assign P1_R2238_U23 = ~(P1_R2238_U48 & P1_R2238_U47); 
assign P1_R2238_U24 = ~(P1_R2238_U53 & P1_R2238_U52); 
assign P1_R2238_U25 = ~(P1_R2238_U58 & P1_R2238_U57); 
assign P1_R2238_U26 = ~(P1_R2238_U63 & P1_R2238_U62); 
assign P1_R2238_U30 = ~P1_R2238_U9; 
assign P1_R2238_U33 = ~(P1_R2238_U9 & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P1_SUB_450_U7 = ~(P1_SUB_450_U9 & P1_SUB_450_U46); 
assign P1_SUB_450_U23 = ~(P1_SUB_450_U48 & P1_SUB_450_U47); 
assign P1_SUB_450_U24 = ~(P1_SUB_450_U53 & P1_SUB_450_U52); 
assign P1_SUB_450_U25 = ~(P1_SUB_450_U58 & P1_SUB_450_U57); 
assign P1_SUB_450_U26 = ~(P1_SUB_450_U63 & P1_SUB_450_U62); 
assign P1_SUB_450_U30 = ~P1_SUB_450_U9; 
assign P1_SUB_450_U33 = ~(P1_SUB_450_U9 & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P1_ADD_405_U5 = ~(P1_ADD_405_U94 & P1_ADD_405_U125); 
assign P1_ADD_405_U8 = ~(P1_ADD_405_U94 & P1_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P1_ADD_405_U85 = ~(P1_ADD_405_U174 & P1_ADD_405_U173); 
assign P1_ADD_405_U97 = ~P1_ADD_405_U94; 
assign P1_ADD_405_U171 = ~(P1_ADD_405_U94 & P1_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P1_ADD_515_U8 = ~(P1_ADD_515_U94 & P1_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P1_ADD_515_U67 = ~(P1_ADD_515_U134 & P1_ADD_515_U133); 
assign P1_ADD_515_U170 = ~(P1_ADD_515_U94 & P1_ADD_515_U7); 
assign U213 = ~(U380 & U379 & U215 & P3_M_IO_N_REG_SCAN_IN); 
assign U384 = ~U382; 
assign U386 = ~U215; 
assign U485 = ~(U215 & BUF2_REG_0__SCAN_IN); 
assign U487 = ~(U215 & BUF2_REG_1__SCAN_IN); 
assign U489 = ~(U215 & BUF2_REG_2__SCAN_IN); 
assign U491 = ~(U215 & BUF2_REG_3__SCAN_IN); 
assign U493 = ~(U215 & BUF2_REG_4__SCAN_IN); 
assign U495 = ~(U215 & BUF2_REG_5__SCAN_IN); 
assign U497 = ~(U215 & BUF2_REG_6__SCAN_IN); 
assign U499 = ~(U215 & BUF2_REG_7__SCAN_IN); 
assign U501 = ~(U215 & BUF2_REG_8__SCAN_IN); 
assign U503 = ~(U215 & BUF2_REG_9__SCAN_IN); 
assign U505 = ~(U215 & BUF2_REG_10__SCAN_IN); 
assign U507 = ~(U215 & BUF2_REG_11__SCAN_IN); 
assign U509 = ~(U215 & BUF2_REG_12__SCAN_IN); 
assign U511 = ~(U215 & BUF2_REG_13__SCAN_IN); 
assign U513 = ~(U215 & BUF2_REG_14__SCAN_IN); 
assign U515 = ~(U215 & BUF2_REG_15__SCAN_IN); 
assign U517 = ~(U215 & BUF2_REG_16__SCAN_IN); 
assign U519 = ~(U215 & BUF2_REG_17__SCAN_IN); 
assign U521 = ~(U215 & BUF2_REG_18__SCAN_IN); 
assign U523 = ~(U215 & BUF2_REG_19__SCAN_IN); 
assign U525 = ~(U215 & BUF2_REG_20__SCAN_IN); 
assign U527 = ~(U215 & BUF2_REG_21__SCAN_IN); 
assign U529 = ~(U215 & BUF2_REG_22__SCAN_IN); 
assign U531 = ~(U215 & BUF2_REG_23__SCAN_IN); 
assign U533 = ~(U215 & BUF2_REG_24__SCAN_IN); 
assign U535 = ~(U215 & BUF2_REG_25__SCAN_IN); 
assign U537 = ~(U215 & BUF2_REG_26__SCAN_IN); 
assign U539 = ~(U215 & BUF2_REG_27__SCAN_IN); 
assign U541 = ~(U215 & BUF2_REG_28__SCAN_IN); 
assign U543 = ~(U215 & BUF2_REG_29__SCAN_IN); 
assign U545 = ~(U215 & BUF2_REG_30__SCAN_IN); 
assign U547 = ~(U215 & BUF2_REG_31__SCAN_IN); 
assign U677 = ~(U382 & P2_ADDRESS_REG_9__SCAN_IN); 
assign U679 = ~(U382 & P2_ADDRESS_REG_8__SCAN_IN); 
assign U681 = ~(U382 & P2_ADDRESS_REG_7__SCAN_IN); 
assign U683 = ~(U382 & P2_ADDRESS_REG_6__SCAN_IN); 
assign U685 = ~(U382 & P2_ADDRESS_REG_5__SCAN_IN); 
assign U687 = ~(U382 & P2_ADDRESS_REG_4__SCAN_IN); 
assign U689 = ~(U382 & P2_ADDRESS_REG_3__SCAN_IN); 
assign U691 = ~(U382 & P2_ADDRESS_REG_2__SCAN_IN); 
assign U693 = ~(U382 & P2_ADDRESS_REG_29__SCAN_IN); 
assign U695 = ~(U382 & P2_ADDRESS_REG_28__SCAN_IN); 
assign U697 = ~(U382 & P2_ADDRESS_REG_27__SCAN_IN); 
assign U699 = ~(U382 & P2_ADDRESS_REG_26__SCAN_IN); 
assign U701 = ~(U382 & P2_ADDRESS_REG_25__SCAN_IN); 
assign U703 = ~(U382 & P2_ADDRESS_REG_24__SCAN_IN); 
assign U705 = ~(U382 & P2_ADDRESS_REG_23__SCAN_IN); 
assign U707 = ~(U382 & P2_ADDRESS_REG_22__SCAN_IN); 
assign U709 = ~(U382 & P2_ADDRESS_REG_21__SCAN_IN); 
assign U711 = ~(U382 & P2_ADDRESS_REG_20__SCAN_IN); 
assign U713 = ~(U382 & P2_ADDRESS_REG_1__SCAN_IN); 
assign U715 = ~(U382 & P2_ADDRESS_REG_19__SCAN_IN); 
assign U717 = ~(U382 & P2_ADDRESS_REG_18__SCAN_IN); 
assign U719 = ~(U382 & P2_ADDRESS_REG_17__SCAN_IN); 
assign U721 = ~(U382 & P2_ADDRESS_REG_16__SCAN_IN); 
assign U723 = ~(U382 & P2_ADDRESS_REG_15__SCAN_IN); 
assign U725 = ~(U382 & P2_ADDRESS_REG_14__SCAN_IN); 
assign U727 = ~(U382 & P2_ADDRESS_REG_13__SCAN_IN); 
assign U729 = ~(U382 & P2_ADDRESS_REG_12__SCAN_IN); 
assign U731 = ~(U382 & P2_ADDRESS_REG_11__SCAN_IN); 
assign U733 = ~(U382 & P2_ADDRESS_REG_10__SCAN_IN); 
assign U735 = ~(U382 & P2_ADDRESS_REG_0__SCAN_IN); 
assign P3_U2390 = P3_U4353 & P3_STATE2_REG_0__SCAN_IN; 
assign P3_U2473 = P3_U2472 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P3_U2475 = P3_U2474 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P3_U2477 = P3_U4470 & P3_U2466; 
assign P3_U2478 = P3_U4470 & P3_U2468; 
assign P3_U2479 = P3_U4470 & P3_U4467; 
assign P3_U2489 = P3_U3090 & P3_U4315; 
assign P3_U2524 = P3_U5558 & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P3_U2526 = P3_U5558 & P3_U3093; 
assign P3_U2593 = P3_U2472 & P3_U3268; 
assign P3_U2594 = P3_U2474 & P3_U3268; 
assign P3_U2596 = P3_U3268 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P3_U3078 = ~(P3_U4308 & P3_U3079); 
assign P3_U3080 = ~(P3_U4308 & P3_STATE_REG_2__SCAN_IN); 
assign P3_U3099 = ~(P3_U4470 & P3_U4332); 
assign P3_U3105 = ~(P3_U4466 & P3_U3085); 
assign P3_U3127 = ~(P3_U4666 & P3_U3121); 
assign P3_U3138 = ~(P3_U3137 & P3_U3128); 
assign P3_U3150 = ~(P3_U3137 & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P3_U3154 = ~(P3_U3404 & P3_U4640); 
assign P3_U3173 = ~(P3_U3475 & P3_U4640); 
assign P3_U3190 = ~(P3_U3545 & P3_U4640); 
assign P3_U3202 = ~(P3_U3616 & P3_U4640); 
assign P3_U3224 = ~(P3_U5505 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_U3225 = ~(P3_U3096 & P3_U3227); 
assign P3_U3267 = ~(P3_U4289 & P3_U3092); 
assign P3_U3269 = ~(P3_U7961 & P3_U7960); 
assign P3_U3366 = P3_U4338 & P3_U4328; 
assign P3_U3659 = P3_U5502 & P3_U5501; 
assign P3_U3669 = P3_U4470 & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign P3_U4307 = ~P3_U3261; 
assign P3_U4322 = ~P3_U3136; 
assign P3_U4347 = ~P3_U3239; 
assign P3_U4446 = ~(P3_U4445 & P3_U2630); 
assign P3_U4447 = ~(NA & P3_U4346); 
assign P3_U4453 = ~(P3_U3088 & U209 & P3_U4346); 
assign P3_U4458 = ~(P3_U4308 & U209); 
assign P3_U4462 = ~(P3_U4461 & P3_U4460); 
assign P3_U4468 = ~P3_U3096; 
assign P3_U4469 = ~P3_U3092; 
assign P3_U4473 = ~(P3_U2483 & P3_INSTQUEUE_REG_1__0__SCAN_IN); 
assign P3_U4474 = ~(P3_U2482 & P3_INSTQUEUE_REG_2__0__SCAN_IN); 
assign P3_U4484 = ~(P3_U2470 & P3_INSTQUEUE_REG_12__0__SCAN_IN); 
assign P3_U4485 = ~(P3_U2469 & P3_INSTQUEUE_REG_13__0__SCAN_IN); 
assign P3_U4486 = ~(P3_U2467 & P3_INSTQUEUE_REG_14__0__SCAN_IN); 
assign P3_U4487 = ~(P3_U2465 & P3_INSTQUEUE_REG_15__0__SCAN_IN); 
assign P3_U4490 = ~(P3_U2483 & P3_INSTQUEUE_REG_1__1__SCAN_IN); 
assign P3_U4491 = ~(P3_U2482 & P3_INSTQUEUE_REG_2__1__SCAN_IN); 
assign P3_U4501 = ~(P3_U2470 & P3_INSTQUEUE_REG_12__1__SCAN_IN); 
assign P3_U4502 = ~(P3_U2469 & P3_INSTQUEUE_REG_13__1__SCAN_IN); 
assign P3_U4503 = ~(P3_U2467 & P3_INSTQUEUE_REG_14__1__SCAN_IN); 
assign P3_U4504 = ~(P3_U2465 & P3_INSTQUEUE_REG_15__1__SCAN_IN); 
assign P3_U4507 = ~(P3_U2483 & P3_INSTQUEUE_REG_1__4__SCAN_IN); 
assign P3_U4508 = ~(P3_U2482 & P3_INSTQUEUE_REG_2__4__SCAN_IN); 
assign P3_U4518 = ~(P3_U2470 & P3_INSTQUEUE_REG_12__4__SCAN_IN); 
assign P3_U4519 = ~(P3_U2469 & P3_INSTQUEUE_REG_13__4__SCAN_IN); 
assign P3_U4520 = ~(P3_U2467 & P3_INSTQUEUE_REG_14__4__SCAN_IN); 
assign P3_U4521 = ~(P3_U2465 & P3_INSTQUEUE_REG_15__4__SCAN_IN); 
assign P3_U4524 = ~(P3_U2483 & P3_INSTQUEUE_REG_1__2__SCAN_IN); 
assign P3_U4525 = ~(P3_U2482 & P3_INSTQUEUE_REG_2__2__SCAN_IN); 
assign P3_U4535 = ~(P3_U2470 & P3_INSTQUEUE_REG_12__2__SCAN_IN); 
assign P3_U4536 = ~(P3_U2469 & P3_INSTQUEUE_REG_13__2__SCAN_IN); 
assign P3_U4537 = ~(P3_U2467 & P3_INSTQUEUE_REG_14__2__SCAN_IN); 
assign P3_U4538 = ~(P3_U2465 & P3_INSTQUEUE_REG_15__2__SCAN_IN); 
assign P3_U4541 = ~(P3_U2483 & P3_INSTQUEUE_REG_1__3__SCAN_IN); 
assign P3_U4542 = ~(P3_U2482 & P3_INSTQUEUE_REG_2__3__SCAN_IN); 
assign P3_U4552 = ~(P3_U2470 & P3_INSTQUEUE_REG_12__3__SCAN_IN); 
assign P3_U4553 = ~(P3_U2469 & P3_INSTQUEUE_REG_13__3__SCAN_IN); 
assign P3_U4554 = ~(P3_U2467 & P3_INSTQUEUE_REG_14__3__SCAN_IN); 
assign P3_U4555 = ~(P3_U2465 & P3_INSTQUEUE_REG_15__3__SCAN_IN); 
assign P3_U4558 = ~(P3_U2483 & P3_INSTQUEUE_REG_1__7__SCAN_IN); 
assign P3_U4559 = ~(P3_U2482 & P3_INSTQUEUE_REG_2__7__SCAN_IN); 
assign P3_U4569 = ~(P3_U2470 & P3_INSTQUEUE_REG_12__7__SCAN_IN); 
assign P3_U4570 = ~(P3_U2469 & P3_INSTQUEUE_REG_13__7__SCAN_IN); 
assign P3_U4571 = ~(P3_U2467 & P3_INSTQUEUE_REG_14__7__SCAN_IN); 
assign P3_U4572 = ~(P3_U2465 & P3_INSTQUEUE_REG_15__7__SCAN_IN); 
assign P3_U4575 = ~(P3_U2483 & P3_INSTQUEUE_REG_1__5__SCAN_IN); 
assign P3_U4576 = ~(P3_U2482 & P3_INSTQUEUE_REG_2__5__SCAN_IN); 
assign P3_U4586 = ~(P3_U2470 & P3_INSTQUEUE_REG_12__5__SCAN_IN); 
assign P3_U4587 = ~(P3_U2469 & P3_INSTQUEUE_REG_13__5__SCAN_IN); 
assign P3_U4588 = ~(P3_U2467 & P3_INSTQUEUE_REG_14__5__SCAN_IN); 
assign P3_U4589 = ~(P3_U2465 & P3_INSTQUEUE_REG_15__5__SCAN_IN); 
assign P3_U4592 = ~(P3_U2483 & P3_INSTQUEUE_REG_1__6__SCAN_IN); 
assign P3_U4593 = ~(P3_U2482 & P3_INSTQUEUE_REG_2__6__SCAN_IN); 
assign P3_U4603 = ~(P3_U2470 & P3_INSTQUEUE_REG_12__6__SCAN_IN); 
assign P3_U4604 = ~(P3_U2469 & P3_INSTQUEUE_REG_13__6__SCAN_IN); 
assign P3_U4605 = ~(P3_U2467 & P3_INSTQUEUE_REG_14__6__SCAN_IN); 
assign P3_U4606 = ~(P3_U2465 & P3_INSTQUEUE_REG_15__6__SCAN_IN); 
assign P3_U4631 = ~(P3_U7957 & P3_U7956 & P3_STATE2_REG_1__SCAN_IN); 
assign P3_U4637 = ~(P3_U4345 & P3_U4354); 
assign P3_U4642 = ~P3_U3137; 
assign P3_U4649 = ~P3_U3132; 
assign P3_U4651 = ~(P3_U3132 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_U4716 = ~P3_U3147; 
assign P3_U4723 = ~(P3_U3147 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U4820 = ~P3_U3161; 
assign P3_U4826 = ~(P3_U3161 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U4871 = ~P3_U3164; 
assign P3_U4878 = ~(P3_U3164 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U5127 = ~P3_U3186; 
assign P3_U5134 = ~(P3_U3186 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U5231 = ~P3_U3194; 
assign P3_U5237 = ~(P3_U3194 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U5281 = ~P3_U3196; 
assign P3_U5288 = ~(P3_U3196 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U5568 = ~(P3_U5558 & P3_U4345); 
assign P3_U5574 = ~(P3_U4345 & P3_U3093); 
assign P3_U5580 = ~(P3_U3132 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U5582 = ~(P3_U4315 & P3_U3123); 
assign P3_U7372 = ~(P3_U3123 & P3_U7371); 
assign P3_U7515 = ~(P3_U4470 & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P3_U7775 = ~P3_U3268; 
assign P3_U7904 = ~(P3_U4292 & P3_STATE_REG_0__SCAN_IN); 
assign P3_U7911 = ~P3_U3086; 
assign P3_U7921 = ~(P3_U4308 & P3_BYTEENABLE_REG_3__SCAN_IN); 
assign P3_U7923 = ~(P3_U4308 & P3_BYTEENABLE_REG_2__SCAN_IN); 
assign P3_U7925 = ~(P3_U4308 & P3_BYTEENABLE_REG_1__SCAN_IN); 
assign P3_U7927 = ~(P3_U4308 & P3_BYTEENABLE_REG_0__SCAN_IN); 
assign P3_U7929 = ~(P3_U3086 & P3_STATE_REG_2__SCAN_IN); 
assign P3_U7936 = ~(P3_U4346 & P3_STATE_REG_0__SCAN_IN); 
assign P3_U7984 = ~(P3_SUB_580_U6 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_U7988 = ~P3_U3286; 
assign P3_U8002 = ~(P3_U3261 & P3_BYTEENABLE_REG_3__SCAN_IN); 
assign P3_U8007 = ~(P3_U8006 & P3_U3081); 
assign P3_U8010 = ~(P3_U3261 & P3_BYTEENABLE_REG_2__SCAN_IN); 
assign P3_U8012 = ~(P3_U3261 & P3_BYTEENABLE_REG_1__SCAN_IN); 
assign P3_U8014 = ~(P3_U3261 & P3_BYTEENABLE_REG_0__SCAN_IN); 
assign P3_U8016 = ~(P3_U4308 & P3_U3264); 
assign P3_U8024 = ~(P3_U4308 & P3_U3263); 
assign P3_U8027 = ~(P3_U4308 & P3_MEMORYFETCH_REG_SCAN_IN); 
assign P3_U8034 = ~P3_U3272; 
assign P3_U8036 = ~(P3_U7645 & P3_U3100); 
assign P2_U2374 = P2_U4468 & P2_STATE2_REG_0__SCAN_IN; 
assign P2_U2444 = P2_U3243 & P2_U3307; 
assign P2_U2523 = P2_U3530 & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P2_U2525 = P2_U3272 & P2_U3530; 
assign P2_U2540 = ~(P2_R2147_U9 | P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P2_U2547 = P2_R2147_U9 & P2_U3532; 
assign P2_U2549 = P2_R2147_U9 & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P2_U2568 = P2_U3582 & P2_U3272; 
assign P2_U2570 = P2_U3582 & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P2_U3260 = ~(P2_U4439 & P2_U3244); 
assign P2_U3261 = ~(P2_U4439 & P2_STATE_REG_2__SCAN_IN); 
assign P2_U3290 = ~(P2_U4595 & P2_U3266); 
assign P2_U3336 = ~(P2_U4649 & P2_U2464); 
assign P2_U3350 = ~(P2_U4648 & P2_U2464); 
assign P2_U3377 = ~(P2_U4645 & P2_U4642); 
assign P2_U3390 = ~(P2_U4645 & P2_U4649); 
assign P2_U3401 = ~(P2_U4645 & P2_U4648); 
assign P2_U3413 = ~(P2_U4645 & P2_U2478); 
assign P2_U3428 = ~(P2_U3376 & P2_U4646 & P2_U3424); 
assign P2_U3439 = ~(P2_U4649 & P2_U2465); 
assign P2_U3450 = ~(P2_U4648 & P2_U2465); 
assign P2_U3485 = ~(P2_U2503 & P2_U4649); 
assign P2_U3496 = ~(P2_U2503 & P2_U4648); 
assign P2_U3529 = ~P2_R2147_U9; 
assign P2_U3580 = ~(P2_U8066 & P2_U8065); 
assign P2_U3581 = ~(P2_U8081 & P2_U8080); 
assign P2_U3694 = P2_U7868 & P2_U7847 & P2_U7831 & P2_U7815; 
assign P2_U3696 = P2_U7866 & P2_U7846 & P2_U7830 & P2_U7814; 
assign P2_U3698 = P2_U7864 & P2_U7845 & P2_U7829 & P2_U7813; 
assign P2_U3700 = P2_U7862 & P2_U7844 & P2_U7828 & P2_U7812; 
assign P2_U3702 = P2_U7860 & P2_U7843 & P2_U7827 & P2_U7811; 
assign P2_U3704 = P2_U7858 & P2_U7842 & P2_U7826 & P2_U7810; 
assign P2_U3706 = P2_U7872 & P2_U7849 & P2_U7833 & P2_U7817; 
assign P2_U3708 = P2_U7870 & P2_U7848 & P2_U7832 & P2_U7816; 
assign P2_U3710 = P2_U4595 & P2_STATE2_REG_0__SCAN_IN; 
assign P2_U4339 = P2_U4595 & P2_U3300; 
assign P2_U4392 = P2_U7908 & P2_U7907; 
assign P2_U4395 = P2_U8079 & P2_U8078; 
assign P2_U4409 = ~P2_U3553; 
assign P2_U4438 = ~P2_U3547; 
assign P2_U4453 = ~(P2_U3718 & P2_U4474); 
assign P2_U4461 = ~P2_U3534; 
assign P2_U4465 = ~(P2_U4474 & U211); 
assign P2_U4569 = ~(P2_U4568 & P2_U3265); 
assign P2_U4570 = ~(NA & P2_U4473); 
assign P2_U4577 = ~(P2_U4576 & P2_U4575); 
assign P2_U4580 = ~(P2_U4410 & P2_STATE_REG_0__SCAN_IN); 
assign P2_U4583 = ~(U211 & P2_U4439); 
assign P2_U4587 = ~(P2_U4586 & P2_U4585); 
assign P2_U4621 = ~(P2_U4474 & P2_U3265); 
assign P2_U4643 = ~P2_U3312; 
assign P2_U4644 = ~P2_U3424; 
assign P2_U4650 = ~P2_U3243; 
assign P2_U4662 = ~(P2_U3312 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U5122 = ~(P2_U3424 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U5285 = ~P2_U3462; 
assign P2_U5294 = ~(P2_U3462 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U5342 = ~P2_U3473; 
assign P2_U5352 = ~(P2_U3473 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U5616 = ~P2_U3530; 
assign P2_U5644 = ~(P2_U4445 & P2_U3303); 
assign P2_U6231 = ~(P2_U4467 & P2_STATE2_REG_1__SCAN_IN); 
assign P2_U6837 = ~(P2_U3547 & P2_BYTEENABLE_REG_1__SCAN_IN); 
assign P2_U6841 = ~(P2_U4187 & P2_U4467); 
assign P2_U7162 = ~(P2_U4430 & P2_U3243); 
assign P2_U7746 = ~(P2_U8003 & P2_U8002 & P2_U4592); 
assign P2_U7747 = ~(P2_U7971 & P2_U7970 & P2_U4592); 
assign P2_U7748 = ~(P2_U7955 & P2_U7954 & P2_U4592); 
assign P2_U7749 = ~(P2_U8035 & P2_U8034 & P2_U4592); 
assign P2_U7750 = ~(P2_U8019 & P2_U8018 & P2_U4592); 
assign P2_U7751 = ~(P2_U7987 & P2_U7986 & P2_U4592); 
assign P2_U7752 = ~(P2_U7939 & P2_U7938 & P2_U4592); 
assign P2_U7753 = ~(P2_U7923 & P2_U7922 & P2_U4592); 
assign P2_U7900 = ~(P2_U4439 & P2_BYTEENABLE_REG_3__SCAN_IN); 
assign P2_U7902 = ~(P2_U4439 & P2_BYTEENABLE_REG_2__SCAN_IN); 
assign P2_U7904 = ~(P2_U4439 & P2_BYTEENABLE_REG_1__SCAN_IN); 
assign P2_U7906 = ~(P2_U4439 & P2_BYTEENABLE_REG_0__SCAN_IN); 
assign P2_U7910 = ~(P2_U4568 & P2_STATE_REG_0__SCAN_IN); 
assign P2_U7916 = ~(P2_U4473 & P2_STATE_REG_0__SCAN_IN); 
assign P2_U8100 = ~P2_U3582; 
assign P2_U8123 = ~(P2_U3547 & P2_BYTEENABLE_REG_3__SCAN_IN); 
assign P2_U8125 = ~(P2_U3547 & P2_BYTEENABLE_REG_2__SCAN_IN); 
assign P2_U8127 = ~(P2_U3547 & P2_BYTEENABLE_REG_0__SCAN_IN); 
assign P2_U8129 = ~(P2_U4439 & P2_U3552); 
assign P2_U8139 = ~(P2_U4439 & P2_U3551); 
assign P2_U8142 = ~(P2_U4439 & P2_MEMORYFETCH_REG_SCAN_IN); 
assign P2_U8148 = ~(P2_U7007 & P2_U3273); 
assign P2_U8152 = ~P2_U3584; 
assign P2_U8153 = ~(P2_U3584 & P2_U3327); 
assign P2_U8155 = ~(P2_U3584 & P2_U3368); 
assign P2_U8157 = ~(P2_U3584 & P2_U3357); 
assign P2_U8159 = ~(P2_U3584 & P2_U3416); 
assign P2_U8161 = ~(P2_U3584 & P2_U3382); 
assign P2_U8163 = ~(P2_U3584 & P2_U3405); 
assign P2_U8165 = ~(P2_U3584 & P2_U3393); 
assign P2_U8167 = ~(P2_U3584 & P2_U3341); 
assign P2_U8169 = ~(P2_U3584 & P2_U3328); 
assign P2_U8171 = ~(P2_U3584 & P2_U3369); 
assign P2_U8173 = ~(P2_U3584 & P2_U3358); 
assign P2_U8175 = ~(P2_U3584 & P2_U3417); 
assign P2_U8177 = ~(P2_U3584 & P2_U3383); 
assign P2_U8179 = ~(P2_U3584 & P2_U3406); 
assign P2_U8181 = ~(P2_U3584 & P2_U3394); 
assign P2_U8183 = ~(P2_U3584 & P2_U3342); 
assign P2_U8185 = ~(P2_U3584 & P2_U3329); 
assign P2_U8187 = ~(P2_U3584 & P2_U3370); 
assign P2_U8189 = ~(P2_U3584 & P2_U3359); 
assign P2_U8191 = ~(P2_U3584 & P2_U3418); 
assign P2_U8193 = ~(P2_U3584 & P2_U3384); 
assign P2_U8195 = ~(P2_U3584 & P2_U3407); 
assign P2_U8197 = ~(P2_U3584 & P2_U3395); 
assign P2_U8199 = ~(P2_U3584 & P2_U3343); 
assign P2_U8201 = ~(P2_U3584 & P2_U3330); 
assign P2_U8203 = ~(P2_U3584 & P2_U3371); 
assign P2_U8205 = ~(P2_U3584 & P2_U3360); 
assign P2_U8207 = ~(P2_U3584 & P2_U3419); 
assign P2_U8209 = ~(P2_U3584 & P2_U3385); 
assign P2_U8211 = ~(P2_U3584 & P2_U3408); 
assign P2_U8213 = ~(P2_U3584 & P2_U3396); 
assign P2_U8215 = ~(P2_U3584 & P2_U3344); 
assign P2_U8217 = ~(P2_U3584 & P2_U3331); 
assign P2_U8219 = ~(P2_U3584 & P2_U3372); 
assign P2_U8221 = ~(P2_U3584 & P2_U3361); 
assign P2_U8223 = ~(P2_U3584 & P2_U3420); 
assign P2_U8225 = ~(P2_U3584 & P2_U3386); 
assign P2_U8227 = ~(P2_U3584 & P2_U3409); 
assign P2_U8229 = ~(P2_U3584 & P2_U3397); 
assign P2_U8231 = ~(P2_U3584 & P2_U3345); 
assign P2_U8233 = ~(P2_U3584 & P2_U3332); 
assign P2_U8235 = ~(P2_U3584 & P2_U3373); 
assign P2_U8237 = ~(P2_U3584 & P2_U3362); 
assign P2_U8239 = ~(P2_U3584 & P2_U3421); 
assign P2_U8241 = ~(P2_U3584 & P2_U3387); 
assign P2_U8243 = ~(P2_U3584 & P2_U3410); 
assign P2_U8245 = ~(P2_U3584 & P2_U3398); 
assign P2_U8247 = ~(P2_U3584 & P2_U3346); 
assign P2_U8249 = ~(P2_U3584 & P2_U3333); 
assign P2_U8251 = ~(P2_U3584 & P2_U3374); 
assign P2_U8253 = ~(P2_U3584 & P2_U3363); 
assign P2_U8255 = ~(P2_U3584 & P2_U3422); 
assign P2_U8257 = ~(P2_U3584 & P2_U3388); 
assign P2_U8259 = ~(P2_U3584 & P2_U3411); 
assign P2_U8261 = ~(P2_U3584 & P2_U3399); 
assign P2_U8263 = ~(P2_U3584 & P2_U3347); 
assign P2_U8265 = ~(P2_U3584 & P2_U3334); 
assign P2_U8267 = ~(P2_U3584 & P2_U3375); 
assign P2_U8269 = ~(P2_U3584 & P2_U3364); 
assign P2_U8271 = ~(P2_U3584 & P2_U3423); 
assign P2_U8273 = ~(P2_U3584 & P2_U3389); 
assign P2_U8275 = ~(P2_U3584 & P2_U3412); 
assign P2_U8277 = ~(P2_U3584 & P2_U3400); 
assign P2_U8279 = ~(P2_U3584 & P2_U3348); 
assign P2_U8397 = ~(P2_R2337_U70 & P2_U3284); 
assign P2_U8428 = ~(P2_SUB_589_U8 & P2_STATE2_REG_1__SCAN_IN); 
assign P2_U8433 = ~(P2_R2238_U7 & P2_U3269); 
assign P1_U2368 = P1_U4235 & P1_STATE2_REG_0__SCAN_IN; 
assign P1_U2436 = P1_U3235 & P1_U3301; 
assign P1_U2446 = P1_U3471 & P1_STATE2_REG_1__SCAN_IN; 
assign P1_U2526 = P1_U5519 & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P1_U2528 = P1_U5519 & P1_U3266; 
assign P1_U2574 = P1_U4379 & P1_U3445; 
assign P1_U2575 = P1_U2460 & P1_U3445; 
assign P1_U2576 = P1_U2462 & P1_U3445; 
assign P1_U2577 = P1_U4380 & P1_U3445; 
assign P1_U2578 = P1_U3445 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P1_U3250 = ~(P1_U4221 & P1_U3251); 
assign P1_U3252 = ~(P1_U4221 & P1_STATE_REG_2__SCAN_IN); 
assign P1_U3272 = ~(P1_U4496 & P1_U3258); 
assign P1_U3278 = ~(P1_U3557 & P1_U3556 & P1_U3555 & P1_U3554); 
assign P1_U3324 = ~(P1_U4542 & P1_U2478); 
assign P1_U3330 = ~(P1_U4541 & P1_U2478); 
assign P1_U3341 = ~(P1_U4538 & P1_U4533); 
assign P1_U3346 = ~(P1_U4538 & P1_U4542); 
assign P1_U3349 = ~(P1_U4538 & P1_U4541); 
assign P1_U3353 = ~(P1_U4538 & P1_U2488); 
assign P1_U3360 = ~(P1_U3340 & P1_U4539 & P1_U3356); 
assign P1_U3363 = ~(P1_U4542 & P1_U2479); 
assign P1_U3366 = ~(P1_U4541 & P1_U2479); 
assign P1_U3377 = ~(P1_U2510 & P1_U4542); 
assign P1_U3380 = ~(P1_U2510 & P1_U4541); 
assign P1_U3438 = ~(P1_U3267 & P1_U5482); 
assign P1_U3455 = ~(P1_U7695 & P1_U7694); 
assign P1_U3530 = P1_U4404 & P1_U4403 & P1_U4402 & P1_U4401; 
assign P1_U3531 = P1_U4408 & P1_U4407 & P1_U4406 & P1_U4405; 
assign P1_U3532 = P1_U4412 & P1_U4411 & P1_U4410 & P1_U4409; 
assign P1_U3538 = P1_U4458 & P1_U4457 & P1_U4459; 
assign P1_U3573 = P1_U4404 & P1_U4403 & P1_U4402 & P1_U4401; 
assign P1_U3574 = P1_U4408 & P1_U4407 & P1_U4406 & P1_U4405; 
assign P1_U3575 = P1_U4412 & P1_U4411 & P1_U4410 & P1_U4409; 
assign P1_U3585 = P1_U4246 & P1_U4241; 
assign P1_U3740 = P1_U5486 & P1_U5485; 
assign P1_U3863 = P1_U5794 & P1_U3408; 
assign P1_U3967 = P1_U3307 & P1_U3408 & P1_U6602; 
assign P1_U4068 = P1_U4405 & P1_U4404 & P1_U4403 & P1_U4401; 
assign P1_U4069 = P1_U4407 & P1_U4406 & P1_U4408; 
assign P1_U4070 = P1_U4412 & P1_U4411 & P1_U4410 & P1_U4409; 
assign P1_U4108 = P1_U7215 & P1_U3264; 
assign P1_U4110 = P1_U7217 & P1_U3265; 
assign P1_U4184 = ~P1_U3452; 
assign P1_U4220 = ~P1_U3433; 
assign P1_U4226 = ~P1_U3320; 
assign P1_U4255 = ~P1_U3432; 
assign P1_U4358 = ~(P1_U4357 & P1_U3257); 
assign P1_U4359 = ~(NA & P1_U4258); 
assign P1_U4367 = ~(P1_U4366 & P1_U4365); 
assign P1_U4370 = ~(U210 & P1_U4221); 
assign P1_U4374 = ~(P1_U4373 & P1_U4372); 
assign P1_U4383 = ~(P1_U4382 & P1_INSTQUEUE_REG_7__3__SCAN_IN); 
assign P1_U4384 = ~(P1_U2472 & P1_INSTQUEUE_REG_0__3__SCAN_IN); 
assign P1_U4388 = ~(P1_U2467 & P1_INSTQUEUE_REG_4__3__SCAN_IN); 
assign P1_U4391 = ~(P1_U2464 & P1_INSTQUEUE_REG_8__3__SCAN_IN); 
assign P1_U4395 = ~(P1_U2458 & P1_INSTQUEUE_REG_12__3__SCAN_IN); 
assign P1_U4416 = ~(P1_U4382 & P1_INSTQUEUE_REG_7__2__SCAN_IN); 
assign P1_U4417 = ~(P1_U2472 & P1_INSTQUEUE_REG_0__2__SCAN_IN); 
assign P1_U4421 = ~(P1_U2467 & P1_INSTQUEUE_REG_4__2__SCAN_IN); 
assign P1_U4424 = ~(P1_U2464 & P1_INSTQUEUE_REG_8__2__SCAN_IN); 
assign P1_U4428 = ~(P1_U2458 & P1_INSTQUEUE_REG_12__2__SCAN_IN); 
assign P1_U4433 = ~(P1_U4382 & P1_INSTQUEUE_REG_7__7__SCAN_IN); 
assign P1_U4434 = ~(P1_U2472 & P1_INSTQUEUE_REG_0__7__SCAN_IN); 
assign P1_U4438 = ~(P1_U2467 & P1_INSTQUEUE_REG_4__7__SCAN_IN); 
assign P1_U4441 = ~(P1_U2464 & P1_INSTQUEUE_REG_8__7__SCAN_IN); 
assign P1_U4445 = ~(P1_U2458 & P1_INSTQUEUE_REG_12__7__SCAN_IN); 
assign P1_U4450 = ~(P1_U3498 & P1_U4381 & P1_INSTQUEUE_REG_7__6__SCAN_IN); 
assign P1_U4453 = ~(P1_U4378 & P1_U4381 & P1_INSTQUEUE_REG_4__6__SCAN_IN); 
assign P1_U4454 = ~(P1_U2456 & P1_U4381 & P1_INSTQUEUE_REG_5__6__SCAN_IN); 
assign P1_U4455 = ~(P1_U2454 & P1_U4381 & P1_INSTQUEUE_REG_6__6__SCAN_IN); 
assign P1_U4461 = ~(P1_U4382 & P1_INSTQUEUE_REG_7__1__SCAN_IN); 
assign P1_U4462 = ~(P1_U2472 & P1_INSTQUEUE_REG_0__1__SCAN_IN); 
assign P1_U4466 = ~(P1_U2467 & P1_INSTQUEUE_REG_4__1__SCAN_IN); 
assign P1_U4469 = ~(P1_U2464 & P1_INSTQUEUE_REG_8__1__SCAN_IN); 
assign P1_U4473 = ~(P1_U2458 & P1_INSTQUEUE_REG_12__1__SCAN_IN); 
assign P1_U4478 = ~(P1_U4382 & P1_INSTQUEUE_REG_7__0__SCAN_IN); 
assign P1_U4479 = ~(P1_U2472 & P1_INSTQUEUE_REG_0__0__SCAN_IN); 
assign P1_U4483 = ~(P1_U2467 & P1_INSTQUEUE_REG_4__0__SCAN_IN); 
assign P1_U4486 = ~(P1_U2464 & P1_INSTQUEUE_REG_8__0__SCAN_IN); 
assign P1_U4490 = ~(P1_U2458 & P1_INSTQUEUE_REG_12__0__SCAN_IN); 
assign P1_U4515 = ~(P1_U7688 & P1_U7687 & P1_STATE2_REG_1__SCAN_IN); 
assign P1_U4534 = ~P1_U3306; 
assign P1_U4537 = ~P1_U3356; 
assign P1_U4543 = ~P1_U3235; 
assign P1_U4552 = ~(P1_U3306 & P1_STATE2_REG_3__SCAN_IN); 
assign P1_U5012 = ~(P1_U3356 & P1_STATE2_REG_3__SCAN_IN); 
assign P1_U5176 = ~P1_U3370; 
assign P1_U5184 = ~(P1_U3370 & P1_STATE2_REG_3__SCAN_IN); 
assign P1_U5233 = ~P1_U3373; 
assign P1_U5242 = ~(P1_U3373 & P1_STATE2_REG_3__SCAN_IN); 
assign P1_U5479 = ~(P1_U4381 & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U5511 = ~P1_U3401; 
assign P1_U5563 = ~(P1_U4203 & P1_U3263); 
assign P1_U6362 = ~(P1_U4203 & P1_U3263); 
assign P1_U6748 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_9__SCAN_IN); 
assign P1_U6751 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_8__SCAN_IN); 
assign P1_U6754 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_7__SCAN_IN); 
assign P1_U6757 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_6__SCAN_IN); 
assign P1_U6761 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_5__SCAN_IN); 
assign P1_U6765 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_4__SCAN_IN); 
assign P1_U6769 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_31__SCAN_IN); 
assign P1_U6773 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_30__SCAN_IN); 
assign P1_U6777 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_3__SCAN_IN); 
assign P1_U6782 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_29__SCAN_IN); 
assign P1_U6786 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_28__SCAN_IN); 
assign P1_U6790 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_27__SCAN_IN); 
assign P1_U6794 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_26__SCAN_IN); 
assign P1_U6798 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_25__SCAN_IN); 
assign P1_U6802 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_24__SCAN_IN); 
assign P1_U6806 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_23__SCAN_IN); 
assign P1_U6810 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_22__SCAN_IN); 
assign P1_U6814 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_21__SCAN_IN); 
assign P1_U6818 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_20__SCAN_IN); 
assign P1_U6822 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_2__SCAN_IN); 
assign P1_U6823 = ~(P1_R2337_U71 & P1_U2352); 
assign P1_U6827 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_19__SCAN_IN); 
assign P1_U6831 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_18__SCAN_IN); 
assign P1_U6835 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_17__SCAN_IN); 
assign P1_U6839 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_16__SCAN_IN); 
assign P1_U6842 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_15__SCAN_IN); 
assign P1_U6845 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_14__SCAN_IN); 
assign P1_U6848 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_13__SCAN_IN); 
assign P1_U6851 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_12__SCAN_IN); 
assign P1_U6854 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_11__SCAN_IN); 
assign P1_U6857 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_10__SCAN_IN); 
assign P1_U6861 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_1__SCAN_IN); 
assign P1_U6866 = ~(P1_U4187 & P1_PHYADDRPOINTER_REG_0__SCAN_IN); 
assign P1_U7065 = ~P1_U3445; 
assign P1_U7218 = ~(P1_U4203 & P1_U3235); 
assign P1_U7468 = ~(P1_U4185 & P1_STATE_REG_0__SCAN_IN); 
assign P1_U7621 = ~P1_U3259; 
assign P1_U7634 = ~(P1_U4221 & P1_BYTEENABLE_REG_3__SCAN_IN); 
assign P1_U7636 = ~(P1_U4221 & P1_BYTEENABLE_REG_2__SCAN_IN); 
assign P1_U7638 = ~(P1_U4221 & P1_BYTEENABLE_REG_1__SCAN_IN); 
assign P1_U7640 = ~(P1_U4221 & P1_BYTEENABLE_REG_0__SCAN_IN); 
assign P1_U7642 = ~(P1_U3259 & P1_STATE_REG_2__SCAN_IN); 
assign P1_U7649 = ~(P1_U4258 & P1_STATE_REG_0__SCAN_IN); 
assign P1_U7711 = ~(P1_SUB_580_U6 & P1_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P1_U7715 = ~P1_U3471; 
assign P1_U7720 = ~P1_U3456; 
assign P1_U7746 = ~(P1_U3433 & P1_BYTEENABLE_REG_3__SCAN_IN); 
assign P1_U7751 = ~(P1_U7750 & P1_U3253); 
assign P1_U7754 = ~(P1_U3433 & P1_BYTEENABLE_REG_2__SCAN_IN); 
assign P1_U7756 = ~(P1_U3433 & P1_BYTEENABLE_REG_1__SCAN_IN); 
assign P1_U7758 = ~(P1_U3433 & P1_BYTEENABLE_REG_0__SCAN_IN); 
assign P1_U7760 = ~(P1_U4221 & P1_U3436); 
assign P1_U7768 = ~(P1_U4221 & P1_U3435); 
assign P1_U7771 = ~(P1_U4221 & P1_MEMORYFETCH_REG_SCAN_IN); 
assign P1_U7786 = ~(P1_U4203 & P1_U3301); 
assign P1_U7789 = ~(P1_U7219 & P1_U3270); 
assign R170_U6 = R170_U15 & P2_ADDRESS_REG_29__SCAN_IN; 
assign R165_U6 = R165_U15 & P1_ADDRESS_REG_29__SCAN_IN; 
assign P3_ADD_526_U57 = ~(P3_ADD_526_U154 & P3_ADD_526_U153); 
assign P3_ADD_526_U60 = ~(P3_ADD_526_U160 & P3_ADD_526_U159); 
assign P3_ADD_526_U112 = ~P3_ADD_526_U13; 
assign P3_ADD_526_U127 = ~P3_ADD_526_U97; 
assign P3_ADD_526_U150 = ~(P3_ADD_526_U13 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_526_U151 = ~(P3_ADD_526_U97 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_552_U57 = ~(P3_ADD_552_U154 & P3_ADD_552_U153); 
assign P3_ADD_552_U60 = ~(P3_ADD_552_U160 & P3_ADD_552_U159); 
assign P3_ADD_552_U112 = ~P3_ADD_552_U13; 
assign P3_ADD_552_U127 = ~P3_ADD_552_U97; 
assign P3_ADD_552_U150 = ~(P3_ADD_552_U13 & P3_EBX_REG_5__SCAN_IN); 
assign P3_ADD_552_U151 = ~(P3_ADD_552_U97 & P3_EBX_REG_4__SCAN_IN); 
assign P3_ADD_546_U57 = ~(P3_ADD_546_U154 & P3_ADD_546_U153); 
assign P3_ADD_546_U60 = ~(P3_ADD_546_U160 & P3_ADD_546_U159); 
assign P3_ADD_546_U112 = ~P3_ADD_546_U13; 
assign P3_ADD_546_U127 = ~P3_ADD_546_U97; 
assign P3_ADD_546_U150 = ~(P3_ADD_546_U13 & P3_EAX_REG_5__SCAN_IN); 
assign P3_ADD_546_U151 = ~(P3_ADD_546_U97 & P3_EAX_REG_4__SCAN_IN); 
assign P3_ADD_476_U68 = ~(P3_ADD_476_U136 & P3_ADD_476_U135); 
assign P3_ADD_476_U95 = ~P3_ADD_476_U8; 
assign P3_ADD_476_U133 = ~(P3_ADD_476_U8 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_531_U74 = ~(P3_ADD_531_U147 & P3_ADD_531_U146); 
assign P3_ADD_531_U99 = ~P3_ADD_531_U9; 
assign P3_ADD_531_U140 = ~(P3_ADD_531_U9 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_SUB_320_U21 = P3_ADD_318_U4 | P3_ADD_318_U71 | P3_PHYADDRPOINTER_REG_0__SCAN_IN; 
assign P3_SUB_320_U50 = ~(P3_SUB_320_U149 & P3_SUB_320_U148); 
assign P3_SUB_320_U105 = ~(P3_ADD_318_U71 & P3_SUB_320_U104); 
assign P3_ADD_505_U16 = ~(P3_ADD_505_U26 & P3_ADD_505_U25); 
assign P3_ADD_505_U19 = ~P3_ADD_505_U10; 
assign P3_ADD_505_U23 = ~(P3_ADD_505_U10 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_ADD_318_U68 = ~(P3_ADD_318_U136 & P3_ADD_318_U135); 
assign P3_ADD_318_U95 = ~P3_ADD_318_U8; 
assign P3_ADD_318_U133 = ~(P3_ADD_318_U8 & P3_PHYADDRPOINTER_REG_4__SCAN_IN); 
assign P3_SUB_370_U31 = ~(P3_SUB_370_U30 & P3_SUB_370_U10); 
assign P3_SUB_370_U49 = ~P3_SUB_370_U23; 
assign P3_SUB_370_U54 = ~P3_SUB_370_U24; 
assign P3_SUB_370_U59 = ~P3_SUB_370_U25; 
assign P3_SUB_370_U64 = ~P3_SUB_370_U26; 
assign P3_SUB_370_U66 = ~(P3_SUB_370_U26 & P3_SUB_370_U9); 
assign P3_ADD_315_U65 = ~(P3_ADD_315_U130 & P3_ADD_315_U129); 
assign P3_ADD_315_U92 = ~P3_ADD_315_U8; 
assign P3_ADD_315_U127 = ~(P3_ADD_315_U8 & P3_PHYADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_467_U68 = ~(P3_ADD_467_U136 & P3_ADD_467_U135); 
assign P3_ADD_467_U95 = ~P3_ADD_467_U8; 
assign P3_ADD_467_U133 = ~(P3_ADD_467_U8 & P3_REIP_REG_4__SCAN_IN); 
assign P3_ADD_430_U68 = ~(P3_ADD_430_U136 & P3_ADD_430_U135); 
assign P3_ADD_430_U95 = ~P3_ADD_430_U8; 
assign P3_ADD_430_U133 = ~(P3_ADD_430_U8 & P3_REIP_REG_4__SCAN_IN); 
assign P3_ADD_380_U74 = ~(P3_ADD_380_U147 & P3_ADD_380_U146); 
assign P3_ADD_380_U99 = ~P3_ADD_380_U9; 
assign P3_ADD_380_U140 = ~(P3_ADD_380_U9 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_344_U74 = ~(P3_ADD_344_U147 & P3_ADD_344_U146); 
assign P3_ADD_344_U99 = ~P3_ADD_344_U9; 
assign P3_ADD_344_U140 = ~(P3_ADD_344_U9 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_339_U68 = ~(P3_ADD_339_U136 & P3_ADD_339_U135); 
assign P3_ADD_339_U95 = ~P3_ADD_339_U8; 
assign P3_ADD_339_U133 = ~(P3_ADD_339_U8 & P3_PHYADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_541_U68 = ~(P3_ADD_541_U136 & P3_ADD_541_U135); 
assign P3_ADD_541_U95 = ~P3_ADD_541_U8; 
assign P3_ADD_541_U133 = ~(P3_ADD_541_U8 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_SUB_355_U31 = ~(P3_SUB_355_U30 & P3_SUB_355_U10); 
assign P3_SUB_355_U49 = ~P3_SUB_355_U23; 
assign P3_SUB_355_U54 = ~P3_SUB_355_U24; 
assign P3_SUB_355_U59 = ~P3_SUB_355_U25; 
assign P3_SUB_355_U64 = ~P3_SUB_355_U26; 
assign P3_SUB_355_U66 = ~(P3_SUB_355_U26 & P3_SUB_355_U9); 
assign P3_SUB_450_U29 = ~(P3_SUB_450_U28 & P3_SUB_450_U8); 
assign P3_SUB_450_U46 = ~P3_SUB_450_U20; 
assign P3_SUB_450_U51 = ~P3_SUB_450_U21; 
assign P3_SUB_450_U56 = ~P3_SUB_450_U22; 
assign P3_SUB_450_U61 = ~P3_SUB_450_U23; 
assign P3_SUB_450_U63 = ~(P3_SUB_450_U23 & P3_SUB_450_U7); 
assign P3_ADD_486_U16 = ~(P3_ADD_486_U26 & P3_ADD_486_U25); 
assign P3_ADD_486_U19 = ~P3_ADD_486_U10; 
assign P3_ADD_486_U23 = ~(P3_ADD_486_U10 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_SUB_485_U29 = ~(P3_SUB_485_U28 & P3_SUB_485_U8); 
assign P3_SUB_485_U46 = ~P3_SUB_485_U20; 
assign P3_SUB_485_U51 = ~P3_SUB_485_U21; 
assign P3_SUB_485_U56 = ~P3_SUB_485_U22; 
assign P3_SUB_485_U61 = ~P3_SUB_485_U23; 
assign P3_SUB_485_U63 = ~(P3_SUB_485_U23 & P3_SUB_485_U7); 
assign P3_ADD_515_U68 = ~(P3_ADD_515_U136 & P3_ADD_515_U135); 
assign P3_ADD_515_U95 = ~P3_ADD_515_U8; 
assign P3_ADD_515_U133 = ~(P3_ADD_515_U8 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_394_U98 = ~P3_ADD_394_U8; 
assign P3_ADD_394_U137 = ~(P3_ADD_394_U8 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_394_U140 = ~(P3_ADD_394_U97 & P3_ADD_394_U7); 
assign P3_SUB_414_U59 = P3_SUB_414_U135 & P3_SUB_414_U134; 
assign P3_SUB_414_U84 = ~P3_SUB_414_U22; 
assign P3_SUB_414_U92 = ~(P3_SUB_414_U91 & P3_EBX_REG_4__SCAN_IN); 
assign P3_SUB_414_U132 = ~(P3_SUB_414_U22 & P3_EBX_REG_5__SCAN_IN); 
assign P3_ADD_441_U68 = ~(P3_ADD_441_U136 & P3_ADD_441_U135); 
assign P3_ADD_441_U95 = ~P3_ADD_441_U8; 
assign P3_ADD_441_U133 = ~(P3_ADD_441_U8 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_349_U74 = ~(P3_ADD_349_U147 & P3_ADD_349_U146); 
assign P3_ADD_349_U99 = ~P3_ADD_349_U9; 
assign P3_ADD_349_U140 = ~(P3_ADD_349_U9 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_405_U98 = ~P3_ADD_405_U8; 
assign P3_ADD_405_U137 = ~(P3_ADD_405_U8 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_405_U140 = ~(P3_ADD_405_U97 & P3_ADD_405_U7); 
assign P3_ADD_553_U74 = ~(P3_ADD_553_U147 & P3_ADD_553_U146); 
assign P3_ADD_553_U99 = ~P3_ADD_553_U9; 
assign P3_ADD_553_U140 = ~(P3_ADD_553_U9 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_558_U74 = ~(P3_ADD_558_U147 & P3_ADD_558_U146); 
assign P3_ADD_558_U99 = ~P3_ADD_558_U9; 
assign P3_ADD_558_U140 = ~(P3_ADD_558_U9 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_385_U74 = ~(P3_ADD_385_U147 & P3_ADD_385_U146); 
assign P3_ADD_385_U99 = ~P3_ADD_385_U9; 
assign P3_ADD_385_U140 = ~(P3_ADD_385_U9 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_547_U74 = ~(P3_ADD_547_U147 & P3_ADD_547_U146); 
assign P3_ADD_547_U99 = ~P3_ADD_547_U9; 
assign P3_ADD_547_U140 = ~(P3_ADD_547_U9 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_SUB_412_U29 = ~(P3_SUB_412_U28 & P3_SUB_412_U8); 
assign P3_SUB_412_U46 = ~P3_SUB_412_U20; 
assign P3_SUB_412_U51 = ~P3_SUB_412_U21; 
assign P3_SUB_412_U56 = ~P3_SUB_412_U22; 
assign P3_SUB_412_U61 = ~P3_SUB_412_U23; 
assign P3_SUB_412_U63 = ~(P3_SUB_412_U23 & P3_SUB_412_U7); 
assign P3_SUB_504_U29 = ~(P3_SUB_504_U28 & P3_SUB_504_U8); 
assign P3_SUB_504_U46 = ~P3_SUB_504_U20; 
assign P3_SUB_504_U51 = ~P3_SUB_504_U21; 
assign P3_SUB_504_U56 = ~P3_SUB_504_U22; 
assign P3_SUB_504_U61 = ~P3_SUB_504_U23; 
assign P3_SUB_504_U63 = ~(P3_SUB_504_U23 & P3_SUB_504_U7); 
assign P3_SUB_401_U31 = ~(P3_SUB_401_U30 & P3_SUB_401_U10); 
assign P3_SUB_401_U49 = ~P3_SUB_401_U23; 
assign P3_SUB_401_U54 = ~P3_SUB_401_U24; 
assign P3_SUB_401_U59 = ~P3_SUB_401_U25; 
assign P3_SUB_401_U64 = ~P3_SUB_401_U26; 
assign P3_SUB_401_U66 = ~(P3_SUB_401_U26 & P3_SUB_401_U9); 
assign P3_SUB_390_U31 = ~(P3_SUB_390_U30 & P3_SUB_390_U10); 
assign P3_SUB_390_U49 = ~P3_SUB_390_U23; 
assign P3_SUB_390_U54 = ~P3_SUB_390_U24; 
assign P3_SUB_390_U59 = ~P3_SUB_390_U25; 
assign P3_SUB_390_U64 = ~P3_SUB_390_U26; 
assign P3_SUB_390_U66 = ~(P3_SUB_390_U26 & P3_SUB_390_U9); 
assign P3_ADD_495_U9 = ~(P3_ADD_495_U18 & P3_ADD_495_U17); 
assign P3_ADD_495_U14 = ~P3_ADD_495_U12; 
assign P3_ADD_495_U15 = ~(P3_ADD_495_U12 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_ADD_494_U68 = ~(P3_ADD_494_U136 & P3_ADD_494_U135); 
assign P3_ADD_494_U95 = ~P3_ADD_494_U8; 
assign P3_ADD_494_U133 = ~(P3_ADD_494_U8 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_536_U68 = ~(P3_ADD_536_U136 & P3_ADD_536_U135); 
assign P3_ADD_536_U95 = ~P3_ADD_536_U8; 
assign P3_ADD_536_U133 = ~(P3_ADD_536_U8 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P2_R2027_U74 = ~(P2_R2027_U147 & P2_R2027_U146); 
assign P2_R2027_U99 = ~P2_R2027_U9; 
assign P2_R2027_U140 = ~(P2_R2027_U9 & P2_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P2_R2337_U66 = ~(P2_R2337_U134 & P2_R2337_U133); 
assign P2_R2337_U67 = ~(P2_R2337_U136 & P2_R2337_U135); 
assign P2_R2337_U96 = ~P2_R2337_U9; 
assign P2_R2337_U131 = ~(P2_R2337_U9 & P2_PHYADDRPOINTER_REG_5__SCAN_IN); 
assign P2_R2147_U8 = ~(P2_R2147_U18 & P2_R2147_U17); 
assign P2_R2238_U31 = ~(P2_R2238_U30 & P2_R2238_U10); 
assign P2_R2238_U49 = ~P2_R2238_U23; 
assign P2_R2238_U54 = ~P2_R2238_U24; 
assign P2_R2238_U59 = ~P2_R2238_U25; 
assign P2_R2238_U64 = ~P2_R2238_U26; 
assign P2_R2238_U66 = ~(P2_R2238_U26 & P2_R2238_U9); 
assign P2_R1957_U71 = ~P2_U3682; 
assign P2_R1957_U72 = ~P2_U3683; 
assign P2_R1957_U104 = P2_U3682 | P2_U3683; 
assign P2_SUB_450_U29 = ~(P2_SUB_450_U28 & P2_SUB_450_U8); 
assign P2_SUB_450_U46 = ~P2_SUB_450_U21; 
assign P2_SUB_450_U51 = ~P2_SUB_450_U22; 
assign P2_SUB_450_U56 = ~P2_SUB_450_U23; 
assign P2_SUB_450_U61 = ~P2_SUB_450_U24; 
assign P2_SUB_450_U63 = ~(P2_SUB_450_U24 & P2_SUB_450_U7); 
assign P2_ADD_394_U98 = ~P2_ADD_394_U8; 
assign P2_ADD_394_U153 = ~(P2_ADD_394_U8 & P2_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P2_ADD_394_U172 = ~(P2_ADD_394_U97 & P2_ADD_394_U7); 
assign P2_ADD_371_1212_U6 = P2_ADD_371_1212_U89 & P2_ADD_371_1212_U11; 
assign P2_ADD_371_1212_U96 = P2_ADD_371_1212_U11 & P2_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P1_R2027_U57 = ~(P1_R2027_U154 & P1_R2027_U153); 
assign P1_R2027_U60 = ~(P1_R2027_U160 & P1_R2027_U159); 
assign P1_R2027_U112 = ~P1_R2027_U13; 
assign P1_R2027_U127 = ~P1_R2027_U97; 
assign P1_R2027_U150 = ~(P1_R2027_U13 & P1_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P1_R2027_U151 = ~(P1_R2027_U97 & P1_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P1_R2337_U68 = ~(P1_R2337_U136 & P1_R2337_U135); 
assign P1_R2337_U95 = ~P1_R2337_U8; 
assign P1_R2337_U133 = ~(P1_R2337_U8 & P1_PHYADDRPOINTER_REG_4__SCAN_IN); 
assign P1_R2096_U68 = ~(P1_R2096_U136 & P1_R2096_U135); 
assign P1_R2096_U95 = ~P1_R2096_U8; 
assign P1_R2096_U133 = ~(P1_R2096_U8 & P1_REIP_REG_4__SCAN_IN); 
assign P1_R2238_U31 = ~(P1_R2238_U30 & P1_R2238_U10); 
assign P1_R2238_U49 = ~P1_R2238_U23; 
assign P1_R2238_U54 = ~P1_R2238_U24; 
assign P1_R2238_U59 = ~P1_R2238_U25; 
assign P1_R2238_U64 = ~P1_R2238_U26; 
assign P1_R2238_U66 = ~(P1_R2238_U26 & P1_R2238_U9); 
assign P1_SUB_450_U31 = ~(P1_SUB_450_U30 & P1_SUB_450_U10); 
assign P1_SUB_450_U49 = ~P1_SUB_450_U23; 
assign P1_SUB_450_U54 = ~P1_SUB_450_U24; 
assign P1_SUB_450_U59 = ~P1_SUB_450_U25; 
assign P1_SUB_450_U64 = ~P1_SUB_450_U26; 
assign P1_SUB_450_U66 = ~(P1_SUB_450_U26 & P1_SUB_450_U9); 
assign P1_ADD_405_U98 = ~P1_ADD_405_U8; 
assign P1_ADD_405_U153 = ~(P1_ADD_405_U8 & P1_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P1_ADD_405_U172 = ~(P1_ADD_405_U97 & P1_ADD_405_U7); 
assign P1_ADD_515_U85 = ~(P1_ADD_515_U170 & P1_ADD_515_U169); 
assign P1_ADD_515_U95 = ~P1_ADD_515_U8; 
assign P1_ADD_515_U151 = ~(P1_ADD_515_U8 & P1_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign U214 = ~(U383 & U381 & R165_U6 & P1_W_R_N_REG_SCAN_IN & P1_M_IO_N_REG_SCAN_IN); 
assign U248 = ~R165_U6; 
assign U249 = ~R170_U6; 
assign U387 = ~(R170_U6 & U208); 
assign U486 = ~(U386 & P2_DATAO_REG_0__SCAN_IN); 
assign U488 = ~(U386 & P2_DATAO_REG_1__SCAN_IN); 
assign U490 = ~(U386 & P2_DATAO_REG_2__SCAN_IN); 
assign U492 = ~(U386 & P2_DATAO_REG_3__SCAN_IN); 
assign U494 = ~(U386 & P2_DATAO_REG_4__SCAN_IN); 
assign U496 = ~(U386 & P2_DATAO_REG_5__SCAN_IN); 
assign U498 = ~(U386 & P2_DATAO_REG_6__SCAN_IN); 
assign U500 = ~(U386 & P2_DATAO_REG_7__SCAN_IN); 
assign U502 = ~(U386 & P2_DATAO_REG_8__SCAN_IN); 
assign U504 = ~(U386 & P2_DATAO_REG_9__SCAN_IN); 
assign U506 = ~(U386 & P2_DATAO_REG_10__SCAN_IN); 
assign U508 = ~(U386 & P2_DATAO_REG_11__SCAN_IN); 
assign U510 = ~(U386 & P2_DATAO_REG_12__SCAN_IN); 
assign U512 = ~(U386 & P2_DATAO_REG_13__SCAN_IN); 
assign U514 = ~(U386 & P2_DATAO_REG_14__SCAN_IN); 
assign U516 = ~(U386 & P2_DATAO_REG_15__SCAN_IN); 
assign U518 = ~(U386 & P2_DATAO_REG_16__SCAN_IN); 
assign U520 = ~(U386 & P2_DATAO_REG_17__SCAN_IN); 
assign U522 = ~(U386 & P2_DATAO_REG_18__SCAN_IN); 
assign U524 = ~(U386 & P2_DATAO_REG_19__SCAN_IN); 
assign U526 = ~(U386 & P2_DATAO_REG_20__SCAN_IN); 
assign U528 = ~(U386 & P2_DATAO_REG_21__SCAN_IN); 
assign U530 = ~(U386 & P2_DATAO_REG_22__SCAN_IN); 
assign U532 = ~(U386 & P2_DATAO_REG_23__SCAN_IN); 
assign U534 = ~(U386 & P2_DATAO_REG_24__SCAN_IN); 
assign U536 = ~(U386 & P2_DATAO_REG_25__SCAN_IN); 
assign U538 = ~(U386 & P2_DATAO_REG_26__SCAN_IN); 
assign U540 = ~(U386 & P2_DATAO_REG_27__SCAN_IN); 
assign U542 = ~(U386 & P2_DATAO_REG_28__SCAN_IN); 
assign U544 = ~(U386 & P2_DATAO_REG_29__SCAN_IN); 
assign U546 = ~(U386 & P2_DATAO_REG_30__SCAN_IN); 
assign U548 = ~(U386 & P2_DATAO_REG_31__SCAN_IN); 
assign U550 = ~(R170_U6 & BUF1_REG_9__SCAN_IN); 
assign U552 = ~(R170_U6 & BUF1_REG_8__SCAN_IN); 
assign U554 = ~(R170_U6 & BUF1_REG_7__SCAN_IN); 
assign U556 = ~(R170_U6 & BUF1_REG_6__SCAN_IN); 
assign U558 = ~(R170_U6 & BUF1_REG_5__SCAN_IN); 
assign U560 = ~(R170_U6 & BUF1_REG_4__SCAN_IN); 
assign U562 = ~(R170_U6 & BUF1_REG_3__SCAN_IN); 
assign U564 = ~(R170_U6 & BUF1_REG_31__SCAN_IN); 
assign U566 = ~(R170_U6 & BUF1_REG_30__SCAN_IN); 
assign U568 = ~(R170_U6 & BUF1_REG_2__SCAN_IN); 
assign U570 = ~(R170_U6 & BUF1_REG_29__SCAN_IN); 
assign U572 = ~(R170_U6 & BUF1_REG_28__SCAN_IN); 
assign U574 = ~(R170_U6 & BUF1_REG_27__SCAN_IN); 
assign U576 = ~(R170_U6 & BUF1_REG_26__SCAN_IN); 
assign U578 = ~(R170_U6 & BUF1_REG_25__SCAN_IN); 
assign U580 = ~(R170_U6 & BUF1_REG_24__SCAN_IN); 
assign U582 = ~(R170_U6 & BUF1_REG_23__SCAN_IN); 
assign U584 = ~(R170_U6 & BUF1_REG_22__SCAN_IN); 
assign U586 = ~(R170_U6 & BUF1_REG_21__SCAN_IN); 
assign U588 = ~(R170_U6 & BUF1_REG_20__SCAN_IN); 
assign U590 = ~(R170_U6 & BUF1_REG_1__SCAN_IN); 
assign U592 = ~(R170_U6 & BUF1_REG_19__SCAN_IN); 
assign U594 = ~(R170_U6 & BUF1_REG_18__SCAN_IN); 
assign U596 = ~(R170_U6 & BUF1_REG_17__SCAN_IN); 
assign U598 = ~(R170_U6 & BUF1_REG_16__SCAN_IN); 
assign U600 = ~(R170_U6 & BUF1_REG_15__SCAN_IN); 
assign U602 = ~(R170_U6 & BUF1_REG_14__SCAN_IN); 
assign U604 = ~(R170_U6 & BUF1_REG_13__SCAN_IN); 
assign U606 = ~(R170_U6 & BUF1_REG_12__SCAN_IN); 
assign U608 = ~(R170_U6 & BUF1_REG_11__SCAN_IN); 
assign U610 = ~(R170_U6 & BUF1_REG_10__SCAN_IN); 
assign U612 = ~(R170_U6 & BUF1_REG_0__SCAN_IN); 
assign U614 = ~(R165_U6 & BUF1_REG_9__SCAN_IN); 
assign U616 = ~(R165_U6 & BUF1_REG_8__SCAN_IN); 
assign U618 = ~(R165_U6 & BUF1_REG_7__SCAN_IN); 
assign U620 = ~(R165_U6 & BUF1_REG_6__SCAN_IN); 
assign U622 = ~(R165_U6 & BUF1_REG_5__SCAN_IN); 
assign U624 = ~(R165_U6 & BUF1_REG_4__SCAN_IN); 
assign U626 = ~(R165_U6 & BUF1_REG_3__SCAN_IN); 
assign U628 = ~(R165_U6 & BUF1_REG_31__SCAN_IN); 
assign U630 = ~(R165_U6 & BUF1_REG_30__SCAN_IN); 
assign U632 = ~(R165_U6 & BUF1_REG_2__SCAN_IN); 
assign U634 = ~(R165_U6 & BUF1_REG_29__SCAN_IN); 
assign U636 = ~(R165_U6 & BUF1_REG_28__SCAN_IN); 
assign U638 = ~(R165_U6 & BUF1_REG_27__SCAN_IN); 
assign U640 = ~(R165_U6 & BUF1_REG_26__SCAN_IN); 
assign U642 = ~(R165_U6 & BUF1_REG_25__SCAN_IN); 
assign U644 = ~(R165_U6 & BUF1_REG_24__SCAN_IN); 
assign U646 = ~(R165_U6 & BUF1_REG_23__SCAN_IN); 
assign U648 = ~(R165_U6 & BUF1_REG_22__SCAN_IN); 
assign U650 = ~(R165_U6 & BUF1_REG_21__SCAN_IN); 
assign U652 = ~(R165_U6 & BUF1_REG_20__SCAN_IN); 
assign U654 = ~(R165_U6 & BUF1_REG_1__SCAN_IN); 
assign U656 = ~(R165_U6 & BUF1_REG_19__SCAN_IN); 
assign U658 = ~(R165_U6 & BUF1_REG_18__SCAN_IN); 
assign U660 = ~(R165_U6 & BUF1_REG_17__SCAN_IN); 
assign U662 = ~(R165_U6 & BUF1_REG_16__SCAN_IN); 
assign U664 = ~(R165_U6 & BUF1_REG_15__SCAN_IN); 
assign U666 = ~(R165_U6 & BUF1_REG_14__SCAN_IN); 
assign U668 = ~(R165_U6 & BUF1_REG_13__SCAN_IN); 
assign U670 = ~(R165_U6 & BUF1_REG_12__SCAN_IN); 
assign U672 = ~(R165_U6 & BUF1_REG_11__SCAN_IN); 
assign U674 = ~(R165_U6 & BUF1_REG_10__SCAN_IN); 
assign U676 = ~(R165_U6 & BUF1_REG_0__SCAN_IN); 
assign U678 = ~(U384 & P3_ADDRESS_REG_9__SCAN_IN); 
assign U680 = ~(U384 & P3_ADDRESS_REG_8__SCAN_IN); 
assign U682 = ~(U384 & P3_ADDRESS_REG_7__SCAN_IN); 
assign U684 = ~(U384 & P3_ADDRESS_REG_6__SCAN_IN); 
assign U686 = ~(U384 & P3_ADDRESS_REG_5__SCAN_IN); 
assign U688 = ~(U384 & P3_ADDRESS_REG_4__SCAN_IN); 
assign U690 = ~(U384 & P3_ADDRESS_REG_3__SCAN_IN); 
assign U692 = ~(U384 & P3_ADDRESS_REG_2__SCAN_IN); 
assign U694 = ~(U384 & P3_ADDRESS_REG_29__SCAN_IN); 
assign U696 = ~(U384 & P3_ADDRESS_REG_28__SCAN_IN); 
assign U698 = ~(U384 & P3_ADDRESS_REG_27__SCAN_IN); 
assign U700 = ~(U384 & P3_ADDRESS_REG_26__SCAN_IN); 
assign U702 = ~(U384 & P3_ADDRESS_REG_25__SCAN_IN); 
assign U704 = ~(U384 & P3_ADDRESS_REG_24__SCAN_IN); 
assign U706 = ~(U384 & P3_ADDRESS_REG_23__SCAN_IN); 
assign U708 = ~(U384 & P3_ADDRESS_REG_22__SCAN_IN); 
assign U710 = ~(U384 & P3_ADDRESS_REG_21__SCAN_IN); 
assign U712 = ~(U384 & P3_ADDRESS_REG_20__SCAN_IN); 
assign U714 = ~(U384 & P3_ADDRESS_REG_1__SCAN_IN); 
assign U716 = ~(U384 & P3_ADDRESS_REG_19__SCAN_IN); 
assign U718 = ~(U384 & P3_ADDRESS_REG_18__SCAN_IN); 
assign U720 = ~(U384 & P3_ADDRESS_REG_17__SCAN_IN); 
assign U722 = ~(U384 & P3_ADDRESS_REG_16__SCAN_IN); 
assign U724 = ~(U384 & P3_ADDRESS_REG_15__SCAN_IN); 
assign U726 = ~(U384 & P3_ADDRESS_REG_14__SCAN_IN); 
assign U728 = ~(U384 & P3_ADDRESS_REG_13__SCAN_IN); 
assign U730 = ~(U384 & P3_ADDRESS_REG_12__SCAN_IN); 
assign U732 = ~(U384 & P3_ADDRESS_REG_11__SCAN_IN); 
assign U734 = ~(U384 & P3_ADDRESS_REG_10__SCAN_IN); 
assign U736 = ~(U384 & P3_ADDRESS_REG_0__SCAN_IN); 
assign P3_U2471 = P3_U4468 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P3_U2476 = P3_U4469 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign P3_U2480 = P3_U4468 & P3_U3100; 
assign P3_U2484 = P3_U4469 & P3_U3100; 
assign P3_U2583 = P3_U7775 & P3_U4468; 
assign P3_U2584 = P3_U7775 & P3_U2472; 
assign P3_U2585 = P3_U7775 & P3_U2474; 
assign P3_U2586 = P3_U7775 & P3_U4469; 
assign P3_U2587 = P3_U7775 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P3_U2592 = P3_U4468 & P3_U3268; 
assign P3_U2595 = P3_U4469 & P3_U3268; 
assign P3_U2597 = P3_U2596 & P3_U4332; 
assign P3_U2598 = P3_U2596 & P3_U2466; 
assign P3_U2599 = P3_U2596 & P3_U2468; 
assign P3_U2600 = P3_U2596 & P3_U4467; 
assign P3_U2635 = ~(P3_U8025 & P3_U8024 & P3_U4335); 
assign P3_U3134 = ~(P3_U4649 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_U3158 = ~(P3_U4642 & P3_U3128); 
assign P3_U3180 = ~(P3_U4649 & P3_U3133); 
assign P3_U3265 = ~(P3_U3099 & P3_U3224); 
assign P3_U3266 = ~(P3_U3223 & P3_U7515); 
assign P3_U3273 = ~(P3_U8036 & P3_U8035); 
assign P3_U3274 = ~(P3_U7921 & P3_U7920); 
assign P3_U3275 = ~(P3_U7923 & P3_U7922); 
assign P3_U3276 = ~(P3_U7925 & P3_U7924); 
assign P3_U3277 = ~(P3_U7927 & P3_U7926); 
assign P3_U3278 = ~(P3_U7936 & P3_U7935); 
assign P3_U3287 = ~(P3_U7984 & P3_U7983); 
assign P3_U3294 = ~(P3_U8017 & P3_U8016); 
assign P3_U3297 = ~(P3_U8027 & P3_U8026); 
assign P3_U3309 = P3_U4447 & P3_STATE_REG_0__SCAN_IN; 
assign P3_U3311 = P3_U4458 & P3_U3078; 
assign P3_U3317 = P3_U4487 & P3_U4486 & P3_U4485 & P3_U4484; 
assign P3_U3322 = P3_U4504 & P3_U4503 & P3_U4502 & P3_U4501; 
assign P3_U3327 = P3_U4521 & P3_U4520 & P3_U4519 & P3_U4518; 
assign P3_U3332 = P3_U4555 & P3_U4554 & P3_U4553 & P3_U4552; 
assign P3_U3337 = P3_U4572 & P3_U4571 & P3_U4570 & P3_U4569; 
assign P3_U3342 = P3_U4538 & P3_U4537 & P3_U4536 & P3_U4535; 
assign P3_U3347 = P3_U4606 & P3_U4605 & P3_U4604 & P3_U4603; 
assign P3_U3352 = P3_U4589 & P3_U4588 & P3_U4587 & P3_U4586; 
assign P3_U3363 = P3_U4631 & P3_U3124; 
assign P3_U4291 = ~P3_U3267; 
assign P3_U4293 = ~P3_U3105; 
assign P3_U4312 = ~P3_U3127; 
assign P3_U4320 = ~P3_U3080; 
assign P3_U4321 = ~P3_U3078; 
assign P3_U4327 = ~(P3_U4149 & P3_U4307); 
assign P3_U4336 = ~(P3_U4347 & P3_U3121); 
assign P3_U4342 = ~P3_U3150; 
assign P3_U4455 = ~(P3_U4453 & P3_U4454); 
assign P3_U4463 = ~(P3_U4462 & P3_U3076); 
assign P3_U4471 = ~P3_U3099; 
assign P3_U4476 = ~(P3_U2479 & P3_INSTQUEUE_REG_4__0__SCAN_IN); 
assign P3_U4477 = ~(P3_U2478 & P3_INSTQUEUE_REG_5__0__SCAN_IN); 
assign P3_U4478 = ~(P3_U2477 & P3_INSTQUEUE_REG_6__0__SCAN_IN); 
assign P3_U4481 = ~(P3_U2475 & P3_INSTQUEUE_REG_9__0__SCAN_IN); 
assign P3_U4482 = ~(P3_U2473 & P3_INSTQUEUE_REG_10__0__SCAN_IN); 
assign P3_U4493 = ~(P3_U2479 & P3_INSTQUEUE_REG_4__1__SCAN_IN); 
assign P3_U4494 = ~(P3_U2478 & P3_INSTQUEUE_REG_5__1__SCAN_IN); 
assign P3_U4495 = ~(P3_U2477 & P3_INSTQUEUE_REG_6__1__SCAN_IN); 
assign P3_U4498 = ~(P3_U2475 & P3_INSTQUEUE_REG_9__1__SCAN_IN); 
assign P3_U4499 = ~(P3_U2473 & P3_INSTQUEUE_REG_10__1__SCAN_IN); 
assign P3_U4510 = ~(P3_U2479 & P3_INSTQUEUE_REG_4__4__SCAN_IN); 
assign P3_U4511 = ~(P3_U2478 & P3_INSTQUEUE_REG_5__4__SCAN_IN); 
assign P3_U4512 = ~(P3_U2477 & P3_INSTQUEUE_REG_6__4__SCAN_IN); 
assign P3_U4515 = ~(P3_U2475 & P3_INSTQUEUE_REG_9__4__SCAN_IN); 
assign P3_U4516 = ~(P3_U2473 & P3_INSTQUEUE_REG_10__4__SCAN_IN); 
assign P3_U4527 = ~(P3_U2479 & P3_INSTQUEUE_REG_4__2__SCAN_IN); 
assign P3_U4528 = ~(P3_U2478 & P3_INSTQUEUE_REG_5__2__SCAN_IN); 
assign P3_U4529 = ~(P3_U2477 & P3_INSTQUEUE_REG_6__2__SCAN_IN); 
assign P3_U4532 = ~(P3_U2475 & P3_INSTQUEUE_REG_9__2__SCAN_IN); 
assign P3_U4533 = ~(P3_U2473 & P3_INSTQUEUE_REG_10__2__SCAN_IN); 
assign P3_U4544 = ~(P3_U2479 & P3_INSTQUEUE_REG_4__3__SCAN_IN); 
assign P3_U4545 = ~(P3_U2478 & P3_INSTQUEUE_REG_5__3__SCAN_IN); 
assign P3_U4546 = ~(P3_U2477 & P3_INSTQUEUE_REG_6__3__SCAN_IN); 
assign P3_U4549 = ~(P3_U2475 & P3_INSTQUEUE_REG_9__3__SCAN_IN); 
assign P3_U4550 = ~(P3_U2473 & P3_INSTQUEUE_REG_10__3__SCAN_IN); 
assign P3_U4561 = ~(P3_U2479 & P3_INSTQUEUE_REG_4__7__SCAN_IN); 
assign P3_U4562 = ~(P3_U2478 & P3_INSTQUEUE_REG_5__7__SCAN_IN); 
assign P3_U4563 = ~(P3_U2477 & P3_INSTQUEUE_REG_6__7__SCAN_IN); 
assign P3_U4566 = ~(P3_U2475 & P3_INSTQUEUE_REG_9__7__SCAN_IN); 
assign P3_U4567 = ~(P3_U2473 & P3_INSTQUEUE_REG_10__7__SCAN_IN); 
assign P3_U4578 = ~(P3_U2479 & P3_INSTQUEUE_REG_4__5__SCAN_IN); 
assign P3_U4579 = ~(P3_U2478 & P3_INSTQUEUE_REG_5__5__SCAN_IN); 
assign P3_U4580 = ~(P3_U2477 & P3_INSTQUEUE_REG_6__5__SCAN_IN); 
assign P3_U4583 = ~(P3_U2475 & P3_INSTQUEUE_REG_9__5__SCAN_IN); 
assign P3_U4584 = ~(P3_U2473 & P3_INSTQUEUE_REG_10__5__SCAN_IN); 
assign P3_U4595 = ~(P3_U2479 & P3_INSTQUEUE_REG_4__6__SCAN_IN); 
assign P3_U4596 = ~(P3_U2478 & P3_INSTQUEUE_REG_5__6__SCAN_IN); 
assign P3_U4597 = ~(P3_U2477 & P3_INSTQUEUE_REG_6__6__SCAN_IN); 
assign P3_U4600 = ~(P3_U2475 & P3_INSTQUEUE_REG_9__6__SCAN_IN); 
assign P3_U4601 = ~(P3_U2473 & P3_INSTQUEUE_REG_10__6__SCAN_IN); 
assign P3_U4653 = ~P3_U3138; 
assign P3_U4768 = ~P3_U3154; 
assign P3_U4775 = ~(P3_U3154 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U4975 = ~P3_U3173; 
assign P3_U4982 = ~(P3_U3173 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U5179 = ~P3_U3190; 
assign P3_U5186 = ~(P3_U3190 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U5239 = ~(P3_U2489 & P3_U3136); 
assign P3_U5290 = ~(P3_U2489 & P3_U3136); 
assign P3_U5341 = ~(P3_U2489 & P3_U3136); 
assign P3_U5383 = ~P3_U3202; 
assign P3_U5390 = ~(P3_U3202 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U5392 = ~(P3_U2489 & P3_U3136); 
assign P3_U5442 = ~(P3_U2489 & P3_U3136); 
assign P3_U5506 = ~P3_U3224; 
assign P3_U5548 = ~P3_U3225; 
assign P3_U5555 = ~(P3_U4345 & P3_U3225); 
assign P3_U5576 = ~(P3_U7988 & P3_STATE2_REG_1__SCAN_IN); 
assign P3_U7373 = ~(P3_U7372 & P3_U3121); 
assign P3_U7382 = ~(P3_U4347 & P3_STATE2_REG_0__SCAN_IN); 
assign P3_U7781 = ~(P3_U2594 & P3_INSTQUEUE_REG_13__7__SCAN_IN); 
assign P3_U7782 = ~(P3_U2593 & P3_INSTQUEUE_REG_14__7__SCAN_IN); 
assign P3_U7797 = ~(P3_U2594 & P3_INSTQUEUE_REG_13__6__SCAN_IN); 
assign P3_U7798 = ~(P3_U2593 & P3_INSTQUEUE_REG_14__6__SCAN_IN); 
assign P3_U7813 = ~(P3_U2594 & P3_INSTQUEUE_REG_13__5__SCAN_IN); 
assign P3_U7814 = ~(P3_U2593 & P3_INSTQUEUE_REG_14__5__SCAN_IN); 
assign P3_U7829 = ~(P3_U2594 & P3_INSTQUEUE_REG_13__4__SCAN_IN); 
assign P3_U7830 = ~(P3_U2593 & P3_INSTQUEUE_REG_14__4__SCAN_IN); 
assign P3_U7845 = ~(P3_U2594 & P3_INSTQUEUE_REG_13__3__SCAN_IN); 
assign P3_U7846 = ~(P3_U2593 & P3_INSTQUEUE_REG_14__3__SCAN_IN); 
assign P3_U7861 = ~(P3_U2594 & P3_INSTQUEUE_REG_13__2__SCAN_IN); 
assign P3_U7862 = ~(P3_U2593 & P3_INSTQUEUE_REG_14__2__SCAN_IN); 
assign P3_U7877 = ~(P3_U2594 & P3_INSTQUEUE_REG_13__1__SCAN_IN); 
assign P3_U7878 = ~(P3_U2593 & P3_INSTQUEUE_REG_14__1__SCAN_IN); 
assign P3_U7893 = ~(P3_U2594 & P3_INSTQUEUE_REG_13__0__SCAN_IN); 
assign P3_U7894 = ~(P3_U2593 & P3_INSTQUEUE_REG_14__0__SCAN_IN); 
assign P3_U7912 = ~(P3_U7911 & P3_U3088); 
assign P3_U7913 = ~(P3_U4449 & P3_U4446 & P3_STATE_REG_1__SCAN_IN); 
assign P3_U7914 = ~(P3_U7904 & P3_STATE_REG_2__SCAN_IN); 
assign P3_U7915 = ~(P3_U4446 & P3_STATE_REG_1__SCAN_IN); 
assign P3_U7930 = ~(P3_U7929 & P3_U7928); 
assign P3_U7962 = ~P3_U3269; 
assign P3_U7964 = ~(P3_U3269 & P3_U3138); 
assign P3_U8003 = ~(P3_U3291 & P3_U4307); 
assign P3_U8009 = ~(P3_U8008 & P3_U8007); 
assign P3_U8013 = ~(P3_U4307 & P3_REIP_REG_1__SCAN_IN); 
assign P3_U8015 = ~(P3_U4307 & P3_U7367); 
assign P3_U8043 = ~(P3_U7988 & P3_FLUSH_REG_SCAN_IN); 
assign P2_U2440 = P2_U3580 & P2_U3428; 
assign P2_U2445 = P2_U4650 & P2_U3307; 
assign P2_U2516 = P2_U5616 & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P2_U2518 = P2_U5616 & P2_U3272; 
assign P2_U2529 = P2_U3582 & P2_U3581; 
assign P2_U2532 = P2_U8100 & P2_U3581; 
assign P2_U2539 = ~(P2_R2147_U8 | P2_R2147_U4); 
assign P2_U2542 = P2_U3529 & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P2_U2553 = P2_R2147_U8 & P2_U3531; 
assign P2_U2556 = P2_R2147_U4 & P2_R2147_U8; 
assign P2_U2563 = P2_U8100 & P2_U3272; 
assign P2_U2566 = P2_U8100 & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign P2_U2817 = ~(P2_U8140 & P2_U8139 & P2_U4463); 
assign P2_U3526 = ~P2_R2147_U8; 
assign P2_U3548 = ~(P2_U4438 & P2_REIP_REG_1__SCAN_IN); 
assign P2_U3583 = ~(P2_U8148 & P2_U8147); 
assign P2_U3585 = ~(P2_U7900 & P2_U7899); 
assign P2_U3586 = ~(P2_U7902 & P2_U7901); 
assign P2_U3587 = ~(P2_U7904 & P2_U7903); 
assign P2_U3588 = ~(P2_U7906 & P2_U7905); 
assign P2_U3589 = ~(P2_U7916 & P2_U7915); 
assign P2_U3608 = ~(P2_U8130 & P2_U8129); 
assign P2_U3611 = ~(P2_U8142 & P2_U8141); 
assign P2_U3671 = ~(P2_U8398 & P2_U8397); 
assign P2_U3691 = P2_U4583 & P2_U3260; 
assign P2_U3693 = P2_U7799 & P2_U7783 & P2_U7767 & P2_U7751; 
assign P2_U3695 = P2_U7798 & P2_U7782 & P2_U7766 & P2_U7750; 
assign P2_U3697 = P2_U7797 & P2_U7781 & P2_U7765 & P2_U7749; 
assign P2_U3699 = P2_U7796 & P2_U7780 & P2_U7764 & P2_U7748; 
assign P2_U3701 = P2_U7795 & P2_U7779 & P2_U7763 & P2_U7747; 
assign P2_U3703 = P2_U7794 & P2_U7778 & P2_U7762 & P2_U7746; 
assign P2_U3705 = P2_U7801 & P2_U7785 & P2_U7769 & P2_U7753; 
assign P2_U3707 = P2_U7800 & P2_U7784 & P2_U7768 & P2_U7752; 
assign P2_U3720 = P2_U4465 & P2_U4453; 
assign P2_U4188 = P2_U6842 & P2_U3313 & P2_U6841; 
assign P2_U4411 = ~P2_U3290; 
assign P2_U4449 = ~P2_U3261; 
assign P2_U4450 = ~P2_U3260; 
assign P2_U4452 = ~(P2_U4182 & P2_U4438); 
assign P2_U4578 = ~(P2_U4570 & P2_U4577 & P2_STATE_REG_0__SCAN_IN); 
assign P2_U4581 = ~(P2_U4580 & P2_STATE_REG_2__SCAN_IN); 
assign P2_U4582 = ~(P2_U7910 & P2_U7909 & P2_U7892); 
assign P2_U4588 = ~(P2_U4587 & P2_U3258); 
assign P2_U4623 = ~(P2_U4622 & P2_U4621); 
assign P2_U4647 = ~P2_U3428; 
assign P2_U4711 = ~P2_U3336; 
assign P2_U4720 = ~(P2_U3336 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U4769 = ~P2_U3350; 
assign P2_U4779 = ~(P2_U3350 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U4884 = ~P2_U3377; 
assign P2_U4894 = ~(P2_U3377 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U4942 = ~P2_U3390; 
assign P2_U4951 = ~(P2_U3390 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U4999 = ~P2_U3401; 
assign P2_U5009 = ~(P2_U3401 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U5057 = ~P2_U3413; 
assign P2_U5066 = ~(P2_U3413 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U5170 = ~P2_U3439; 
assign P2_U5179 = ~(P2_U3439 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U5227 = ~P2_U3450; 
assign P2_U5237 = ~(P2_U3450 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U5400 = ~P2_U3485; 
assign P2_U5409 = ~(P2_U3485 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U5457 = ~P2_U3496; 
assign P2_U5467 = ~(P2_U3496 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U5672 = ~(P2_U4461 & P2_U3284); 
assign P2_U6569 = ~(P2_U4461 & P2_U3284); 
assign P2_U6855 = ~(P2_U4461 & P2_STATE2_REG_0__SCAN_IN); 
assign P2_U7140 = ~(P2_U4430 & P2_U3428); 
assign P2_U7151 = ~(P2_U4430 & P2_U3580); 
assign P2_U7891 = ~(P2_U4572 & P2_U4569 & P2_STATE_REG_1__SCAN_IN); 
assign P2_U7893 = ~(P2_U4569 & P2_STATE_REG_1__SCAN_IN); 
assign P2_U8067 = ~P2_U3580; 
assign P2_U8082 = ~P2_U3581; 
assign P2_U8124 = ~(P2_U3606 & P2_U4438); 
assign P2_U8126 = ~(P2_U3607 & P2_U4438); 
assign P2_U8128 = ~(P2_U4438 & P2_REIP_REG_0__SCAN_IN); 
assign P2_U8154 = ~(P2_U8152 & P2_U3431); 
assign P2_U8156 = ~(P2_U8152 & P2_U3465); 
assign P2_U8158 = ~(P2_U8152 & P2_U3454); 
assign P2_U8160 = ~(P2_U8152 & P2_U3511); 
assign P2_U8162 = ~(P2_U8152 & P2_U3477); 
assign P2_U8164 = ~(P2_U8152 & P2_U3500); 
assign P2_U8166 = ~(P2_U8152 & P2_U3488); 
assign P2_U8168 = ~(P2_U8152 & P2_U3442); 
assign P2_U8170 = ~(P2_U8152 & P2_U3432); 
assign P2_U8172 = ~(P2_U8152 & P2_U3466); 
assign P2_U8174 = ~(P2_U8152 & P2_U3455); 
assign P2_U8176 = ~(P2_U8152 & P2_U3512); 
assign P2_U8178 = ~(P2_U8152 & P2_U3478); 
assign P2_U8180 = ~(P2_U8152 & P2_U3501); 
assign P2_U8182 = ~(P2_U8152 & P2_U3489); 
assign P2_U8184 = ~(P2_U8152 & P2_U3443); 
assign P2_U8186 = ~(P2_U8152 & P2_U3433); 
assign P2_U8188 = ~(P2_U8152 & P2_U3467); 
assign P2_U8190 = ~(P2_U8152 & P2_U3456); 
assign P2_U8192 = ~(P2_U8152 & P2_U3513); 
assign P2_U8194 = ~(P2_U8152 & P2_U3479); 
assign P2_U8196 = ~(P2_U8152 & P2_U3502); 
assign P2_U8198 = ~(P2_U8152 & P2_U3490); 
assign P2_U8200 = ~(P2_U8152 & P2_U3444); 
assign P2_U8202 = ~(P2_U8152 & P2_U3434); 
assign P2_U8204 = ~(P2_U8152 & P2_U3468); 
assign P2_U8206 = ~(P2_U8152 & P2_U3457); 
assign P2_U8208 = ~(P2_U8152 & P2_U3514); 
assign P2_U8210 = ~(P2_U8152 & P2_U3480); 
assign P2_U8212 = ~(P2_U8152 & P2_U3503); 
assign P2_U8214 = ~(P2_U8152 & P2_U3491); 
assign P2_U8216 = ~(P2_U8152 & P2_U3445); 
assign P2_U8218 = ~(P2_U8152 & P2_U3435); 
assign P2_U8220 = ~(P2_U8152 & P2_U3469); 
assign P2_U8222 = ~(P2_U8152 & P2_U3458); 
assign P2_U8224 = ~(P2_U8152 & P2_U3515); 
assign P2_U8226 = ~(P2_U8152 & P2_U3481); 
assign P2_U8228 = ~(P2_U8152 & P2_U3504); 
assign P2_U8230 = ~(P2_U8152 & P2_U3492); 
assign P2_U8232 = ~(P2_U8152 & P2_U3446); 
assign P2_U8234 = ~(P2_U8152 & P2_U3436); 
assign P2_U8236 = ~(P2_U8152 & P2_U3470); 
assign P2_U8238 = ~(P2_U8152 & P2_U3459); 
assign P2_U8240 = ~(P2_U8152 & P2_U3516); 
assign P2_U8242 = ~(P2_U8152 & P2_U3482); 
assign P2_U8244 = ~(P2_U8152 & P2_U3505); 
assign P2_U8246 = ~(P2_U8152 & P2_U3493); 
assign P2_U8248 = ~(P2_U8152 & P2_U3447); 
assign P2_U8250 = ~(P2_U8152 & P2_U3437); 
assign P2_U8252 = ~(P2_U8152 & P2_U3471); 
assign P2_U8254 = ~(P2_U8152 & P2_U3460); 
assign P2_U8256 = ~(P2_U8152 & P2_U3517); 
assign P2_U8258 = ~(P2_U8152 & P2_U3483); 
assign P2_U8260 = ~(P2_U8152 & P2_U3506); 
assign P2_U8262 = ~(P2_U8152 & P2_U3494); 
assign P2_U8264 = ~(P2_U8152 & P2_U3448); 
assign P2_U8266 = ~(P2_U8152 & P2_U3438); 
assign P2_U8268 = ~(P2_U8152 & P2_U3472); 
assign P2_U8270 = ~(P2_U8152 & P2_U3461); 
assign P2_U8272 = ~(P2_U8152 & P2_U3518); 
assign P2_U8274 = ~(P2_U8152 & P2_U3484); 
assign P2_U8276 = ~(P2_U8152 & P2_U3507); 
assign P2_U8278 = ~(P2_U8152 & P2_U3495); 
assign P2_U8280 = ~(P2_U8152 & P2_U3449); 
assign P2_U8371 = ~(P2_R2337_U66 & P2_U3284); 
assign P2_U8375 = ~(P2_R2337_U67 & P2_U3284); 
assign P1_U2432 = P1_U3455 & P1_U3360; 
assign P1_U2437 = P1_U4543 & P1_U3301; 
assign P1_U2535 = P1_U5511 & P1_U3438; 
assign P1_U2540 = P1_U3438 & P1_U3401; 
assign P1_U2565 = P1_U7065 & P1_U4379; 
assign P1_U2566 = P1_U7065 & P1_U2460; 
assign P1_U2567 = P1_U7065 & P1_U2462; 
assign P1_U2568 = P1_U7065 & P1_U4380; 
assign P1_U2569 = P1_U7065 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign P1_U2579 = P1_U2578 & P1_U3498; 
assign P1_U2580 = P1_U2578 & P1_U2454; 
assign P1_U2581 = P1_U2578 & P1_U2456; 
assign P1_U2582 = P1_U2578 & P1_U4378; 
assign P1_U2605 = P1_U3533 & P1_U2607 & P1_U3532 & P1_U3531 & P1_U3530; 
assign P1_U2608 = P1_U7787 & P1_U7786; 
assign P1_U2804 = ~(P1_U7769 & P1_U7768 & P1_U4243); 
assign P1_U3442 = ~(P1_U5479 & P1_U5478); 
assign P1_U3457 = ~(P1_U7789 & P1_U7788); 
assign P1_U3458 = ~(P1_U7634 & P1_U7633); 
assign P1_U3459 = ~(P1_U7636 & P1_U7635); 
assign P1_U3460 = ~(P1_U7638 & P1_U7637); 
assign P1_U3461 = ~(P1_U7640 & P1_U7639); 
assign P1_U3462 = ~(P1_U7649 & P1_U7648); 
assign P1_U3470 = ~(P1_U7711 & P1_U7710); 
assign P1_U3483 = ~(P1_U7761 & P1_U7760); 
assign P1_U3486 = ~(P1_U7771 & P1_U7770); 
assign P1_U3495 = P1_U4370 & P1_U3250; 
assign P1_U3508 = P1_U4386 & P1_U4385 & P1_U4384 & P1_U4383; 
assign P1_U3509 = P1_U4390 & P1_U4389 & P1_U4388 & P1_U4387; 
assign P1_U3510 = P1_U4394 & P1_U4393 & P1_U4392 & P1_U4391; 
assign P1_U3511 = P1_U4398 & P1_U4397 & P1_U4396 & P1_U4395; 
assign P1_U3512 = P1_U4436 & P1_U4435 & P1_U4434 & P1_U4433; 
assign P1_U3513 = P1_U4440 & P1_U4439 & P1_U4438 & P1_U4437; 
assign P1_U3514 = P1_U4444 & P1_U4443 & P1_U4442 & P1_U4441; 
assign P1_U3515 = P1_U4448 & P1_U4447 & P1_U4446 & P1_U4445; 
assign P1_U3516 = P1_U4419 & P1_U4418 & P1_U4417 & P1_U4416; 
assign P1_U3517 = P1_U4423 & P1_U4422 & P1_U4421 & P1_U4420; 
assign P1_U3518 = P1_U4427 & P1_U4426 & P1_U4425 & P1_U4424; 
assign P1_U3519 = P1_U4431 & P1_U4430 & P1_U4429 & P1_U4428; 
assign P1_U3536 = P1_U4453 & P1_U4452 & P1_U4451 & P1_U4450; 
assign P1_U3537 = P1_U4455 & P1_U4454 & P1_U4456; 
assign P1_U3560 = P1_U4481 & P1_U4480 & P1_U4479 & P1_U4478; 
assign P1_U3561 = P1_U4485 & P1_U4484 & P1_U4483 & P1_U4482; 
assign P1_U3562 = P1_U4489 & P1_U4488 & P1_U4487 & P1_U4486; 
assign P1_U3563 = P1_U4493 & P1_U4492 & P1_U4491 & P1_U4490; 
assign P1_U3564 = P1_U4464 & P1_U4463 & P1_U4462 & P1_U4461; 
assign P1_U3565 = P1_U4468 & P1_U4467 & P1_U4466 & P1_U4465; 
assign P1_U3566 = P1_U4472 & P1_U4471 & P1_U4470 & P1_U4469; 
assign P1_U3567 = P1_U4476 & P1_U4475 & P1_U4474 & P1_U4473; 
assign P1_U3569 = P1_U4419 & P1_U4418 & P1_U4417 & P1_U4416; 
assign P1_U3570 = P1_U4423 & P1_U4422 & P1_U4421 & P1_U4420; 
assign P1_U3571 = P1_U4427 & P1_U4426 & P1_U4425 & P1_U4424; 
assign P1_U3572 = P1_U4431 & P1_U4430 & P1_U4429 & P1_U4428; 
assign P1_U3582 = P1_U4515 & P1_U3297; 
assign P1_U3887 = P1_U4241 & P1_U4244 & P1_U6362; 
assign P1_U4112 = P1_U7218 & P1_U7217; 
assign P1_U4173 = ~(P1_U3576 & P1_U2607 & P1_U3575 & P1_U3574 & P1_U3573); 
assign P1_U4232 = ~P1_U3252; 
assign P1_U4233 = ~P1_U3250; 
assign P1_U4240 = ~(P1_U3963 & P1_U4220); 
assign P1_U4368 = ~(P1_U4359 & P1_U4367 & P1_STATE_REG_0__SCAN_IN); 
assign P1_U4375 = ~(P1_U4374 & P1_U3248); 
assign P1_U4400 = ~P1_U3278; 
assign P1_U4497 = ~P1_U3272; 
assign P1_U4540 = ~P1_U3360; 
assign P1_U4602 = ~P1_U3324; 
assign P1_U4610 = ~(P1_U3324 & P1_STATE2_REG_3__SCAN_IN); 
assign P1_U4660 = ~P1_U3330; 
assign P1_U4669 = ~(P1_U3330 & P1_STATE2_REG_3__SCAN_IN); 
assign P1_U4775 = ~P1_U3341; 
assign P1_U4784 = ~(P1_U3341 & P1_STATE2_REG_3__SCAN_IN); 
assign P1_U4833 = ~P1_U3346; 
assign P1_U4841 = ~(P1_U3346 & P1_STATE2_REG_3__SCAN_IN); 
assign P1_U4890 = ~P1_U3349; 
assign P1_U4899 = ~(P1_U3349 & P1_STATE2_REG_3__SCAN_IN); 
assign P1_U4948 = ~P1_U3353; 
assign P1_U4956 = ~(P1_U3353 & P1_STATE2_REG_3__SCAN_IN); 
assign P1_U5061 = ~P1_U3363; 
assign P1_U5069 = ~(P1_U3363 & P1_STATE2_REG_3__SCAN_IN); 
assign P1_U5118 = ~P1_U3366; 
assign P1_U5127 = ~(P1_U3366 & P1_STATE2_REG_3__SCAN_IN); 
assign P1_U5291 = ~P1_U3377; 
assign P1_U5299 = ~(P1_U3377 & P1_STATE2_REG_3__SCAN_IN); 
assign P1_U5348 = ~P1_U3380; 
assign P1_U5357 = ~(P1_U3380 & P1_STATE2_REG_3__SCAN_IN); 
assign P1_U5483 = ~P1_U3438; 
assign P1_U5534 = ~(P1_U7715 & P1_STATE2_REG_1__SCAN_IN); 
assign P1_U6612 = ~(P1_U4255 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U6778 = ~(P1_R2337_U68 & P1_U2352); 
assign P1_U7070 = ~(P1_U2577 & P1_INSTQUEUE_REG_12__7__SCAN_IN); 
assign P1_U7071 = ~(P1_U2576 & P1_INSTQUEUE_REG_13__7__SCAN_IN); 
assign P1_U7072 = ~(P1_U2575 & P1_INSTQUEUE_REG_14__7__SCAN_IN); 
assign P1_U7073 = ~(P1_U2574 & P1_INSTQUEUE_REG_15__7__SCAN_IN); 
assign P1_U7097 = ~(P1_U4203 & P1_U3360); 
assign P1_U7102 = ~(P1_U2577 & P1_INSTQUEUE_REG_12__6__SCAN_IN); 
assign P1_U7103 = ~(P1_U2576 & P1_INSTQUEUE_REG_13__6__SCAN_IN); 
assign P1_U7104 = ~(P1_U2575 & P1_INSTQUEUE_REG_14__6__SCAN_IN); 
assign P1_U7105 = ~(P1_U2574 & P1_INSTQUEUE_REG_15__6__SCAN_IN); 
assign P1_U7119 = ~(P1_U2577 & P1_INSTQUEUE_REG_12__5__SCAN_IN); 
assign P1_U7120 = ~(P1_U2576 & P1_INSTQUEUE_REG_13__5__SCAN_IN); 
assign P1_U7121 = ~(P1_U2575 & P1_INSTQUEUE_REG_14__5__SCAN_IN); 
assign P1_U7122 = ~(P1_U2574 & P1_INSTQUEUE_REG_15__5__SCAN_IN); 
assign P1_U7136 = ~(P1_U2577 & P1_INSTQUEUE_REG_12__4__SCAN_IN); 
assign P1_U7137 = ~(P1_U2576 & P1_INSTQUEUE_REG_13__4__SCAN_IN); 
assign P1_U7138 = ~(P1_U2575 & P1_INSTQUEUE_REG_14__4__SCAN_IN); 
assign P1_U7139 = ~(P1_U2574 & P1_INSTQUEUE_REG_15__4__SCAN_IN); 
assign P1_U7151 = ~(P1_U2577 & P1_INSTQUEUE_REG_12__3__SCAN_IN); 
assign P1_U7152 = ~(P1_U2576 & P1_INSTQUEUE_REG_13__3__SCAN_IN); 
assign P1_U7153 = ~(P1_U2575 & P1_INSTQUEUE_REG_14__3__SCAN_IN); 
assign P1_U7154 = ~(P1_U2574 & P1_INSTQUEUE_REG_15__3__SCAN_IN); 
assign P1_U7168 = ~(P1_U2577 & P1_INSTQUEUE_REG_12__2__SCAN_IN); 
assign P1_U7169 = ~(P1_U2576 & P1_INSTQUEUE_REG_13__2__SCAN_IN); 
assign P1_U7170 = ~(P1_U2575 & P1_INSTQUEUE_REG_14__2__SCAN_IN); 
assign P1_U7171 = ~(P1_U2574 & P1_INSTQUEUE_REG_15__2__SCAN_IN); 
assign P1_U7185 = ~(P1_U2577 & P1_INSTQUEUE_REG_12__1__SCAN_IN); 
assign P1_U7186 = ~(P1_U2576 & P1_INSTQUEUE_REG_13__1__SCAN_IN); 
assign P1_U7187 = ~(P1_U2575 & P1_INSTQUEUE_REG_14__1__SCAN_IN); 
assign P1_U7188 = ~(P1_U2574 & P1_INSTQUEUE_REG_15__1__SCAN_IN); 
assign P1_U7202 = ~(P1_U2577 & P1_INSTQUEUE_REG_12__0__SCAN_IN); 
assign P1_U7203 = ~(P1_U2576 & P1_INSTQUEUE_REG_13__0__SCAN_IN); 
assign P1_U7204 = ~(P1_U2575 & P1_INSTQUEUE_REG_14__0__SCAN_IN); 
assign P1_U7205 = ~(P1_U2574 & P1_INSTQUEUE_REG_15__0__SCAN_IN); 
assign P1_U7216 = ~(P1_U4203 & P1_U3455); 
assign P1_U7470 = ~(P1_U4110 & P1_U7218); 
assign P1_U7495 = ~(P1_U4071 & P1_U2607 & P1_U4070 & P1_U4069 & P1_U4068); 
assign P1_U7622 = ~(P1_U7621 & P1_U3261); 
assign P1_U7623 = ~(P1_U4361 & P1_U4358 & P1_STATE_REG_1__SCAN_IN); 
assign P1_U7624 = ~(P1_U7468 & P1_STATE_REG_2__SCAN_IN); 
assign P1_U7625 = ~(P1_U4358 & P1_STATE_REG_1__SCAN_IN); 
assign P1_U7643 = ~(P1_U7642 & P1_U7641); 
assign P1_U7696 = ~P1_U3455; 
assign P1_U7747 = ~(P1_U3480 & P1_U4220); 
assign P1_U7753 = ~(P1_U7752 & P1_U7751); 
assign P1_U7757 = ~(P1_U4220 & P1_REIP_REG_1__SCAN_IN); 
assign P1_U7759 = ~(P1_U4220 & P1_U6599); 
assign P1_U7794 = ~(P1_U7715 & P1_STATE2_REG_1__SCAN_IN & P1_FLUSH_REG_SCAN_IN); 
assign P3_ADD_526_U16 = ~(P3_ADD_526_U83 & P3_ADD_526_U112); 
assign P3_ADD_526_U96 = ~(P3_ADD_526_U112 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_526_U149 = ~(P3_ADD_526_U112 & P3_ADD_526_U12); 
assign P3_ADD_526_U152 = ~(P3_ADD_526_U127 & P3_ADD_526_U8); 
assign P3_ADD_552_U16 = ~(P3_ADD_552_U83 & P3_ADD_552_U112); 
assign P3_ADD_552_U96 = ~(P3_ADD_552_U112 & P3_EBX_REG_5__SCAN_IN); 
assign P3_ADD_552_U149 = ~(P3_ADD_552_U112 & P3_ADD_552_U12); 
assign P3_ADD_552_U152 = ~(P3_ADD_552_U127 & P3_ADD_552_U8); 
assign P3_ADD_546_U16 = ~(P3_ADD_546_U83 & P3_ADD_546_U112); 
assign P3_ADD_546_U96 = ~(P3_ADD_546_U112 & P3_EAX_REG_5__SCAN_IN); 
assign P3_ADD_546_U149 = ~(P3_ADD_546_U112 & P3_ADD_546_U12); 
assign P3_ADD_546_U152 = ~(P3_ADD_546_U127 & P3_ADD_546_U8); 
assign P3_ADD_476_U10 = ~(P3_ADD_476_U95 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_476_U134 = ~(P3_ADD_476_U95 & P3_ADD_476_U9); 
assign P3_ADD_531_U11 = ~(P3_ADD_531_U99 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_531_U141 = ~(P3_ADD_531_U99 & P3_ADD_531_U10); 
assign P3_SUB_320_U17 = P3_SUB_320_U105 & P3_SUB_320_U21; 
assign P3_SUB_320_U58 = ~P3_ADD_318_U68; 
assign P3_SUB_320_U83 = ~P3_SUB_320_U21; 
assign P3_SUB_320_U134 = ~(P3_ADD_318_U68 & P3_SUB_320_U21); 
assign P3_ADD_505_U12 = ~(P3_ADD_505_U19 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_ADD_505_U24 = ~(P3_ADD_505_U19 & P3_ADD_505_U11); 
assign P3_ADD_318_U10 = ~(P3_ADD_318_U95 & P3_PHYADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_318_U134 = ~(P3_ADD_318_U95 & P3_ADD_318_U9); 
assign P3_SUB_370_U32 = ~(P3_SUB_370_U31 & P3_SUB_370_U29); 
assign P3_SUB_370_U65 = ~(P3_SUB_370_U64 & P3_SUB_370_U30); 
assign P3_ADD_315_U10 = ~(P3_ADD_315_U92 & P3_PHYADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_315_U128 = ~(P3_ADD_315_U92 & P3_ADD_315_U9); 
assign P3_ADD_467_U10 = ~(P3_ADD_467_U95 & P3_REIP_REG_4__SCAN_IN); 
assign P3_ADD_467_U134 = ~(P3_ADD_467_U95 & P3_ADD_467_U9); 
assign P3_ADD_430_U10 = ~(P3_ADD_430_U95 & P3_REIP_REG_4__SCAN_IN); 
assign P3_ADD_430_U134 = ~(P3_ADD_430_U95 & P3_ADD_430_U9); 
assign P3_ADD_380_U11 = ~(P3_ADD_380_U99 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_380_U141 = ~(P3_ADD_380_U99 & P3_ADD_380_U10); 
assign P3_ADD_344_U11 = ~(P3_ADD_344_U99 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_344_U141 = ~(P3_ADD_344_U99 & P3_ADD_344_U10); 
assign P3_ADD_339_U10 = ~(P3_ADD_339_U95 & P3_PHYADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_339_U134 = ~(P3_ADD_339_U95 & P3_ADD_339_U9); 
assign P3_ADD_541_U10 = ~(P3_ADD_541_U95 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_541_U134 = ~(P3_ADD_541_U95 & P3_ADD_541_U9); 
assign P3_SUB_355_U32 = ~(P3_SUB_355_U31 & P3_SUB_355_U29); 
assign P3_SUB_355_U65 = ~(P3_SUB_355_U64 & P3_SUB_355_U30); 
assign P3_SUB_450_U30 = ~(P3_SUB_450_U29 & P3_SUB_450_U26); 
assign P3_SUB_450_U62 = ~(P3_SUB_450_U61 & P3_SUB_450_U28); 
assign P3_ADD_486_U12 = ~(P3_ADD_486_U19 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_ADD_486_U24 = ~(P3_ADD_486_U19 & P3_ADD_486_U11); 
assign P3_SUB_485_U30 = ~(P3_SUB_485_U29 & P3_SUB_485_U26); 
assign P3_SUB_485_U62 = ~(P3_SUB_485_U61 & P3_SUB_485_U28); 
assign P3_ADD_515_U10 = ~(P3_ADD_515_U95 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_515_U134 = ~(P3_ADD_515_U95 & P3_ADD_515_U9); 
assign P3_ADD_394_U10 = ~(P3_ADD_394_U98 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_394_U93 = P3_ADD_394_U140 & P3_ADD_394_U139; 
assign P3_ADD_394_U138 = ~(P3_ADD_394_U98 & P3_ADD_394_U9); 
assign P3_SUB_414_U18 = P3_SUB_414_U92 & P3_SUB_414_U22; 
assign P3_SUB_414_U23 = ~(P3_SUB_414_U26 & P3_SUB_414_U56 & P3_SUB_414_U84); 
assign P3_SUB_414_U89 = ~(P3_SUB_414_U84 & P3_SUB_414_U56); 
assign P3_SUB_414_U133 = ~(P3_SUB_414_U84 & P3_SUB_414_U56); 
assign P3_ADD_441_U10 = ~(P3_ADD_441_U95 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_441_U134 = ~(P3_ADD_441_U95 & P3_ADD_441_U9); 
assign P3_ADD_349_U11 = ~(P3_ADD_349_U99 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_349_U141 = ~(P3_ADD_349_U99 & P3_ADD_349_U10); 
assign P3_ADD_405_U10 = ~(P3_ADD_405_U98 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_405_U93 = P3_ADD_405_U140 & P3_ADD_405_U139; 
assign P3_ADD_405_U138 = ~(P3_ADD_405_U98 & P3_ADD_405_U9); 
assign P3_ADD_553_U11 = ~(P3_ADD_553_U99 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_553_U141 = ~(P3_ADD_553_U99 & P3_ADD_553_U10); 
assign P3_ADD_558_U11 = ~(P3_ADD_558_U99 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_558_U141 = ~(P3_ADD_558_U99 & P3_ADD_558_U10); 
assign P3_ADD_385_U11 = ~(P3_ADD_385_U99 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_385_U141 = ~(P3_ADD_385_U99 & P3_ADD_385_U10); 
assign P3_ADD_547_U11 = ~(P3_ADD_547_U99 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_547_U141 = ~(P3_ADD_547_U99 & P3_ADD_547_U10); 
assign P3_SUB_412_U30 = ~(P3_SUB_412_U29 & P3_SUB_412_U26); 
assign P3_SUB_412_U62 = ~(P3_SUB_412_U61 & P3_SUB_412_U28); 
assign P3_SUB_504_U30 = ~(P3_SUB_504_U29 & P3_SUB_504_U26); 
assign P3_SUB_504_U62 = ~(P3_SUB_504_U61 & P3_SUB_504_U28); 
assign P3_SUB_401_U32 = ~(P3_SUB_401_U31 & P3_SUB_401_U29); 
assign P3_SUB_401_U65 = ~(P3_SUB_401_U64 & P3_SUB_401_U30); 
assign P3_SUB_390_U32 = ~(P3_SUB_390_U31 & P3_SUB_390_U29); 
assign P3_SUB_390_U65 = ~(P3_SUB_390_U64 & P3_SUB_390_U30); 
assign P3_ADD_495_U16 = ~(P3_ADD_495_U14 & P3_ADD_495_U11); 
assign P3_ADD_494_U10 = ~(P3_ADD_494_U95 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_494_U134 = ~(P3_ADD_494_U95 & P3_ADD_494_U9); 
assign P3_ADD_536_U10 = ~(P3_ADD_536_U95 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_536_U134 = ~(P3_ADD_536_U95 & P3_ADD_536_U9); 
assign P2_R2027_U11 = ~(P2_R2027_U99 & P2_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P2_R2027_U141 = ~(P2_R2027_U99 & P2_R2027_U10); 
assign P2_R2337_U11 = ~(P2_R2337_U96 & P2_PHYADDRPOINTER_REG_5__SCAN_IN); 
assign P2_R2337_U132 = ~(P2_R2337_U96 & P2_R2337_U10); 
assign P2_R2238_U32 = ~(P2_R2238_U31 & P2_R2238_U29); 
assign P2_R2238_U65 = ~(P2_R2238_U64 & P2_R2238_U30); 
assign P2_R1957_U148 = ~(P2_U3682 & P2_R1957_U72); 
assign P2_R1957_U149 = ~(P2_U3683 & P2_R1957_U71); 
assign P2_SUB_450_U30 = ~(P2_SUB_450_U29 & P2_SUB_450_U27); 
assign P2_SUB_450_U62 = ~(P2_SUB_450_U61 & P2_SUB_450_U28); 
assign P2_ADD_394_U10 = ~(P2_ADD_394_U98 & P2_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P2_ADD_394_U95 = P2_ADD_394_U172 & P2_ADD_394_U171; 
assign P2_ADD_394_U154 = ~(P2_ADD_394_U98 & P2_ADD_394_U9); 
assign P2_ADD_371_1212_U9 = P2_ADD_371_1212_U6 & P2_ADD_371_1212_U90; 
assign P2_ADD_371_1212_U97 = P2_ADD_371_1212_U6 & P2_ADD_371_1212_U98; 
assign P2_ADD_371_1212_U99 = P2_ADD_371_1212_U6 & P2_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P1_R2027_U16 = ~(P1_R2027_U83 & P1_R2027_U112); 
assign P1_R2027_U96 = ~(P1_R2027_U112 & P1_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P1_R2027_U149 = ~(P1_R2027_U112 & P1_R2027_U12); 
assign P1_R2027_U152 = ~(P1_R2027_U127 & P1_R2027_U8); 
assign P1_R2337_U10 = ~(P1_R2337_U95 & P1_PHYADDRPOINTER_REG_4__SCAN_IN); 
assign P1_R2337_U134 = ~(P1_R2337_U95 & P1_R2337_U9); 
assign P1_R2096_U10 = ~(P1_R2096_U95 & P1_REIP_REG_4__SCAN_IN); 
assign P1_R2096_U134 = ~(P1_R2096_U95 & P1_R2096_U9); 
assign P1_R2238_U32 = ~(P1_R2238_U31 & P1_R2238_U29); 
assign P1_R2238_U65 = ~(P1_R2238_U64 & P1_R2238_U30); 
assign P1_SUB_450_U32 = ~(P1_SUB_450_U31 & P1_SUB_450_U29); 
assign P1_SUB_450_U65 = ~(P1_SUB_450_U64 & P1_SUB_450_U30); 
assign P1_ADD_405_U10 = ~(P1_ADD_405_U98 & P1_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P1_ADD_405_U95 = P1_ADD_405_U172 & P1_ADD_405_U171; 
assign P1_ADD_405_U154 = ~(P1_ADD_405_U98 & P1_ADD_405_U9); 
assign P1_ADD_515_U10 = ~(P1_ADD_515_U95 & P1_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P1_ADD_515_U152 = ~(P1_ADD_515_U95 & P1_ADD_515_U9); 
assign U212 = ~(U208 & R170_U6 & U214); 
assign U250 = ~(U214 & U387); 
assign U251 = ~(U486 & U485); 
assign U252 = ~(U488 & U487); 
assign U253 = ~(U490 & U489); 
assign U254 = ~(U492 & U491); 
assign U255 = ~(U494 & U493); 
assign U256 = ~(U496 & U495); 
assign U257 = ~(U498 & U497); 
assign U258 = ~(U500 & U499); 
assign U259 = ~(U502 & U501); 
assign U260 = ~(U504 & U503); 
assign U261 = ~(U506 & U505); 
assign U262 = ~(U508 & U507); 
assign U263 = ~(U510 & U509); 
assign U264 = ~(U512 & U511); 
assign U265 = ~(U514 & U513); 
assign U266 = ~(U516 & U515); 
assign U267 = ~(U518 & U517); 
assign U268 = ~(U520 & U519); 
assign U269 = ~(U522 & U521); 
assign U270 = ~(U524 & U523); 
assign U271 = ~(U526 & U525); 
assign U272 = ~(U528 & U527); 
assign U273 = ~(U530 & U529); 
assign U274 = ~(U532 & U531); 
assign U275 = ~(U534 & U533); 
assign U276 = ~(U536 & U535); 
assign U277 = ~(U538 & U537); 
assign U278 = ~(U540 & U539); 
assign U279 = ~(U542 & U541); 
assign U280 = ~(U544 & U543); 
assign U281 = ~(U546 & U545); 
assign U282 = ~(U548 & U547); 
assign U347 = ~(U678 & U677); 
assign U348 = ~(U680 & U679); 
assign U349 = ~(U682 & U681); 
assign U350 = ~(U684 & U683); 
assign U351 = ~(U686 & U685); 
assign U352 = ~(U688 & U687); 
assign U353 = ~(U690 & U689); 
assign U354 = ~(U692 & U691); 
assign U355 = ~(U694 & U693); 
assign U356 = ~(U696 & U695); 
assign U357 = ~(U698 & U697); 
assign U358 = ~(U700 & U699); 
assign U359 = ~(U702 & U701); 
assign U360 = ~(U704 & U703); 
assign U361 = ~(U706 & U705); 
assign U362 = ~(U708 & U707); 
assign U363 = ~(U710 & U709); 
assign U364 = ~(U712 & U711); 
assign U365 = ~(U714 & U713); 
assign U366 = ~(U716 & U715); 
assign U367 = ~(U718 & U717); 
assign U368 = ~(U720 & U719); 
assign U369 = ~(U722 & U721); 
assign U370 = ~(U724 & U723); 
assign U371 = ~(U726 & U725); 
assign U372 = ~(U728 & U727); 
assign U373 = ~(U730 & U729); 
assign U374 = ~(U732 & U731); 
assign U375 = ~(U734 & U733); 
assign U376 = ~(U736 & U735); 
assign U385 = ~U214; 
assign U549 = ~(U249 & BUF2_REG_9__SCAN_IN); 
assign U551 = ~(U249 & BUF2_REG_8__SCAN_IN); 
assign U553 = ~(U249 & BUF2_REG_7__SCAN_IN); 
assign U555 = ~(U249 & BUF2_REG_6__SCAN_IN); 
assign U557 = ~(U249 & BUF2_REG_5__SCAN_IN); 
assign U559 = ~(U249 & BUF2_REG_4__SCAN_IN); 
assign U561 = ~(U249 & BUF2_REG_3__SCAN_IN); 
assign U563 = ~(U249 & BUF2_REG_31__SCAN_IN); 
assign U565 = ~(U249 & BUF2_REG_30__SCAN_IN); 
assign U567 = ~(U249 & BUF2_REG_2__SCAN_IN); 
assign U569 = ~(U249 & BUF2_REG_29__SCAN_IN); 
assign U571 = ~(U249 & BUF2_REG_28__SCAN_IN); 
assign U573 = ~(U249 & BUF2_REG_27__SCAN_IN); 
assign U575 = ~(U249 & BUF2_REG_26__SCAN_IN); 
assign U577 = ~(U249 & BUF2_REG_25__SCAN_IN); 
assign U579 = ~(U249 & BUF2_REG_24__SCAN_IN); 
assign U581 = ~(U249 & BUF2_REG_23__SCAN_IN); 
assign U583 = ~(U249 & BUF2_REG_22__SCAN_IN); 
assign U585 = ~(U249 & BUF2_REG_21__SCAN_IN); 
assign U587 = ~(U249 & BUF2_REG_20__SCAN_IN); 
assign U589 = ~(U249 & BUF2_REG_1__SCAN_IN); 
assign U591 = ~(U249 & BUF2_REG_19__SCAN_IN); 
assign U593 = ~(U249 & BUF2_REG_18__SCAN_IN); 
assign U595 = ~(U249 & BUF2_REG_17__SCAN_IN); 
assign U597 = ~(U249 & BUF2_REG_16__SCAN_IN); 
assign U599 = ~(U249 & BUF2_REG_15__SCAN_IN); 
assign U601 = ~(U249 & BUF2_REG_14__SCAN_IN); 
assign U603 = ~(U249 & BUF2_REG_13__SCAN_IN); 
assign U605 = ~(U249 & BUF2_REG_12__SCAN_IN); 
assign U607 = ~(U249 & BUF2_REG_11__SCAN_IN); 
assign U609 = ~(U249 & BUF2_REG_10__SCAN_IN); 
assign U611 = ~(U249 & BUF2_REG_0__SCAN_IN); 
assign U613 = ~(DATAI_9_ & U248); 
assign U615 = ~(DATAI_8_ & U248); 
assign U617 = ~(DATAI_7_ & U248); 
assign U619 = ~(DATAI_6_ & U248); 
assign U621 = ~(DATAI_5_ & U248); 
assign U623 = ~(DATAI_4_ & U248); 
assign U625 = ~(DATAI_3_ & U248); 
assign U627 = ~(DATAI_31_ & U248); 
assign U629 = ~(DATAI_30_ & U248); 
assign U631 = ~(DATAI_2_ & U248); 
assign U633 = ~(DATAI_29_ & U248); 
assign U635 = ~(DATAI_28_ & U248); 
assign U637 = ~(DATAI_27_ & U248); 
assign U639 = ~(DATAI_26_ & U248); 
assign U641 = ~(DATAI_25_ & U248); 
assign U643 = ~(DATAI_24_ & U248); 
assign U645 = ~(DATAI_23_ & U248); 
assign U647 = ~(DATAI_22_ & U248); 
assign U649 = ~(DATAI_21_ & U248); 
assign U651 = ~(DATAI_20_ & U248); 
assign U653 = ~(DATAI_1_ & U248); 
assign U655 = ~(DATAI_19_ & U248); 
assign U657 = ~(DATAI_18_ & U248); 
assign U659 = ~(DATAI_17_ & U248); 
assign U661 = ~(DATAI_16_ & U248); 
assign U663 = ~(DATAI_15_ & U248); 
assign U665 = ~(DATAI_14_ & U248); 
assign U667 = ~(DATAI_13_ & U248); 
assign U669 = ~(DATAI_12_ & U248); 
assign U671 = ~(DATAI_11_ & U248); 
assign U673 = ~(DATAI_10_ & U248); 
assign U675 = ~(DATAI_0_ & U248); 
assign P3_U2379 = P3_U4322 & P3_U4312; 
assign P3_U2381 = P3_U4312 & P3_STATE2_REG_3__SCAN_IN; 
assign P3_U2413 = P3_U4312 & BUF2_REG_0__SCAN_IN; 
assign P3_U2414 = P3_U4312 & BUF2_REG_1__SCAN_IN; 
assign P3_U2415 = P3_U4312 & BUF2_REG_2__SCAN_IN; 
assign P3_U2416 = P3_U4312 & BUF2_REG_3__SCAN_IN; 
assign P3_U2417 = P3_U4312 & BUF2_REG_4__SCAN_IN; 
assign P3_U2418 = P3_U4312 & BUF2_REG_5__SCAN_IN; 
assign P3_U2419 = P3_U4312 & BUF2_REG_6__SCAN_IN; 
assign P3_U2420 = P3_U4312 & BUF2_REG_7__SCAN_IN; 
assign P3_U2533 = P3_U5548 & P3_U3265; 
assign P3_U2538 = P3_U3265 & P3_U3225; 
assign P3_U2543 = P3_U3272 & P3_U3266; 
assign P3_U2548 = P3_U8034 & P3_U3266; 
assign P3_U2573 = P3_U4291 & P3_U3273; 
assign P3_U2578 = P3_U3273 & P3_U3267; 
assign P3_U2588 = P3_U2587 & P3_U4332; 
assign P3_U2589 = P3_U2587 & P3_U2466; 
assign P3_U2590 = P3_U2587 & P3_U2468; 
assign P3_U2591 = P3_U2587 & P3_U4467; 
assign P3_U2638 = ~(P3_U8013 & P3_U8012 & P3_U4327); 
assign P3_U2639 = ~(P3_U8003 & P3_U8002 & P3_U4327); 
assign P3_U3106 = ~(P3_U4293 & P3_U2630); 
assign P3_U3139 = ~(P3_U3180 & P3_U4651); 
assign P3_U3141 = ~(P3_U3150 & P3_U3158); 
assign P3_U3293 = ~(P3_U8015 & P3_U8014); 
assign P3_U3302 = ~(P3_U8043 & P3_U8042); 
assign P3_U3353 = P3_U2352 & P3_U4293; 
assign P3_U3387 = P3_U4723 & P3_U4312; 
assign P3_U3405 = P3_U4775 & P3_U4312; 
assign P3_U3423 = P3_U4826 & P3_U4312; 
assign P3_U3440 = P3_U4878 & P3_U4312; 
assign P3_U3458 = P3_U4930 & P3_U4312; 
assign P3_U3476 = P3_U4982 & P3_U4312; 
assign P3_U3493 = P3_U5033 & P3_U4312; 
assign P3_U3528 = P3_U5134 & P3_U4312; 
assign P3_U3546 = P3_U5186 & P3_U4312; 
assign P3_U3564 = P3_U5237 & P3_U4312; 
assign P3_U3582 = P3_U5288 & P3_U4312; 
assign P3_U3599 = P3_U5339 & P3_U4312; 
assign P3_U3617 = P3_U5390 & P3_U4312; 
assign P3_U3635 = P3_U5440 & P3_U4312; 
assign P3_U3684 = P3_U5576 & P3_U5574; 
assign P3_U3986 = P3_U4293 & P3_U2390; 
assign P3_U4030 = P3_U4329 & P3_U4328 & P3_U4336; 
assign P3_U4151 = P3_U7373 & P3_U3135; 
assign P3_U4343 = ~P3_U3158; 
assign P3_U4355 = ~(P3_U4321 & P3_REIP_REG_31__SCAN_IN); 
assign P3_U4356 = ~(P3_U4320 & P3_REIP_REG_30__SCAN_IN); 
assign P3_U4358 = ~(P3_U4321 & P3_REIP_REG_30__SCAN_IN); 
assign P3_U4359 = ~(P3_U4320 & P3_REIP_REG_29__SCAN_IN); 
assign P3_U4361 = ~(P3_U4321 & P3_REIP_REG_29__SCAN_IN); 
assign P3_U4362 = ~(P3_U4320 & P3_REIP_REG_28__SCAN_IN); 
assign P3_U4364 = ~(P3_U4321 & P3_REIP_REG_28__SCAN_IN); 
assign P3_U4365 = ~(P3_U4320 & P3_REIP_REG_27__SCAN_IN); 
assign P3_U4367 = ~(P3_U4321 & P3_REIP_REG_27__SCAN_IN); 
assign P3_U4368 = ~(P3_U4320 & P3_REIP_REG_26__SCAN_IN); 
assign P3_U4370 = ~(P3_U4321 & P3_REIP_REG_26__SCAN_IN); 
assign P3_U4371 = ~(P3_U4320 & P3_REIP_REG_25__SCAN_IN); 
assign P3_U4373 = ~(P3_U4321 & P3_REIP_REG_25__SCAN_IN); 
assign P3_U4374 = ~(P3_U4320 & P3_REIP_REG_24__SCAN_IN); 
assign P3_U4376 = ~(P3_U4321 & P3_REIP_REG_24__SCAN_IN); 
assign P3_U4377 = ~(P3_U4320 & P3_REIP_REG_23__SCAN_IN); 
assign P3_U4379 = ~(P3_U4321 & P3_REIP_REG_23__SCAN_IN); 
assign P3_U4380 = ~(P3_U4320 & P3_REIP_REG_22__SCAN_IN); 
assign P3_U4382 = ~(P3_U4321 & P3_REIP_REG_22__SCAN_IN); 
assign P3_U4383 = ~(P3_U4320 & P3_REIP_REG_21__SCAN_IN); 
assign P3_U4385 = ~(P3_U4321 & P3_REIP_REG_21__SCAN_IN); 
assign P3_U4386 = ~(P3_U4320 & P3_REIP_REG_20__SCAN_IN); 
assign P3_U4388 = ~(P3_U4321 & P3_REIP_REG_20__SCAN_IN); 
assign P3_U4389 = ~(P3_U4320 & P3_REIP_REG_19__SCAN_IN); 
assign P3_U4391 = ~(P3_U4321 & P3_REIP_REG_19__SCAN_IN); 
assign P3_U4392 = ~(P3_U4320 & P3_REIP_REG_18__SCAN_IN); 
assign P3_U4394 = ~(P3_U4321 & P3_REIP_REG_18__SCAN_IN); 
assign P3_U4395 = ~(P3_U4320 & P3_REIP_REG_17__SCAN_IN); 
assign P3_U4397 = ~(P3_U4321 & P3_REIP_REG_17__SCAN_IN); 
assign P3_U4398 = ~(P3_U4320 & P3_REIP_REG_16__SCAN_IN); 
assign P3_U4400 = ~(P3_U4321 & P3_REIP_REG_16__SCAN_IN); 
assign P3_U4401 = ~(P3_U4320 & P3_REIP_REG_15__SCAN_IN); 
assign P3_U4403 = ~(P3_U4321 & P3_REIP_REG_15__SCAN_IN); 
assign P3_U4404 = ~(P3_U4320 & P3_REIP_REG_14__SCAN_IN); 
assign P3_U4406 = ~(P3_U4321 & P3_REIP_REG_14__SCAN_IN); 
assign P3_U4407 = ~(P3_U4320 & P3_REIP_REG_13__SCAN_IN); 
assign P3_U4409 = ~(P3_U4321 & P3_REIP_REG_13__SCAN_IN); 
assign P3_U4410 = ~(P3_U4320 & P3_REIP_REG_12__SCAN_IN); 
assign P3_U4412 = ~(P3_U4321 & P3_REIP_REG_12__SCAN_IN); 
assign P3_U4413 = ~(P3_U4320 & P3_REIP_REG_11__SCAN_IN); 
assign P3_U4415 = ~(P3_U4321 & P3_REIP_REG_11__SCAN_IN); 
assign P3_U4416 = ~(P3_U4320 & P3_REIP_REG_10__SCAN_IN); 
assign P3_U4418 = ~(P3_U4321 & P3_REIP_REG_10__SCAN_IN); 
assign P3_U4419 = ~(P3_U4320 & P3_REIP_REG_9__SCAN_IN); 
assign P3_U4421 = ~(P3_U4321 & P3_REIP_REG_9__SCAN_IN); 
assign P3_U4422 = ~(P3_U4320 & P3_REIP_REG_8__SCAN_IN); 
assign P3_U4424 = ~(P3_U4321 & P3_REIP_REG_8__SCAN_IN); 
assign P3_U4425 = ~(P3_U4320 & P3_REIP_REG_7__SCAN_IN); 
assign P3_U4427 = ~(P3_U4321 & P3_REIP_REG_7__SCAN_IN); 
assign P3_U4428 = ~(P3_U4320 & P3_REIP_REG_6__SCAN_IN); 
assign P3_U4430 = ~(P3_U4321 & P3_REIP_REG_6__SCAN_IN); 
assign P3_U4431 = ~(P3_U4320 & P3_REIP_REG_5__SCAN_IN); 
assign P3_U4433 = ~(P3_U4321 & P3_REIP_REG_5__SCAN_IN); 
assign P3_U4434 = ~(P3_U4320 & P3_REIP_REG_4__SCAN_IN); 
assign P3_U4436 = ~(P3_U4321 & P3_REIP_REG_4__SCAN_IN); 
assign P3_U4437 = ~(P3_U4320 & P3_REIP_REG_3__SCAN_IN); 
assign P3_U4439 = ~(P3_U4321 & P3_REIP_REG_3__SCAN_IN); 
assign P3_U4440 = ~(P3_U4320 & P3_REIP_REG_2__SCAN_IN); 
assign P3_U4442 = ~(P3_U4321 & P3_REIP_REG_2__SCAN_IN); 
assign P3_U4443 = ~(P3_U4320 & P3_REIP_REG_1__SCAN_IN); 
assign P3_U4451 = ~(P3_U7912 & P3_U4450 & P3_U7913); 
assign P3_U4456 = ~(P3_U3309 & P3_U4455); 
assign P3_U4459 = ~(P3_U3312 & P3_U7915); 
assign P3_U4472 = ~(P3_U2484 & P3_INSTQUEUE_REG_0__0__SCAN_IN); 
assign P3_U4475 = ~(P3_U2480 & P3_INSTQUEUE_REG_3__0__SCAN_IN); 
assign P3_U4479 = ~(P3_U4471 & P3_INSTQUEUE_REG_7__0__SCAN_IN); 
assign P3_U4480 = ~(P3_U2476 & P3_INSTQUEUE_REG_8__0__SCAN_IN); 
assign P3_U4483 = ~(P3_U2471 & P3_INSTQUEUE_REG_11__0__SCAN_IN); 
assign P3_U4489 = ~(P3_U2484 & P3_INSTQUEUE_REG_0__1__SCAN_IN); 
assign P3_U4492 = ~(P3_U2480 & P3_INSTQUEUE_REG_3__1__SCAN_IN); 
assign P3_U4496 = ~(P3_U4471 & P3_INSTQUEUE_REG_7__1__SCAN_IN); 
assign P3_U4497 = ~(P3_U2476 & P3_INSTQUEUE_REG_8__1__SCAN_IN); 
assign P3_U4500 = ~(P3_U2471 & P3_INSTQUEUE_REG_11__1__SCAN_IN); 
assign P3_U4506 = ~(P3_U2484 & P3_INSTQUEUE_REG_0__4__SCAN_IN); 
assign P3_U4509 = ~(P3_U2480 & P3_INSTQUEUE_REG_3__4__SCAN_IN); 
assign P3_U4513 = ~(P3_U4471 & P3_INSTQUEUE_REG_7__4__SCAN_IN); 
assign P3_U4514 = ~(P3_U2476 & P3_INSTQUEUE_REG_8__4__SCAN_IN); 
assign P3_U4517 = ~(P3_U2471 & P3_INSTQUEUE_REG_11__4__SCAN_IN); 
assign P3_U4523 = ~(P3_U2484 & P3_INSTQUEUE_REG_0__2__SCAN_IN); 
assign P3_U4526 = ~(P3_U2480 & P3_INSTQUEUE_REG_3__2__SCAN_IN); 
assign P3_U4530 = ~(P3_U4471 & P3_INSTQUEUE_REG_7__2__SCAN_IN); 
assign P3_U4531 = ~(P3_U2476 & P3_INSTQUEUE_REG_8__2__SCAN_IN); 
assign P3_U4534 = ~(P3_U2471 & P3_INSTQUEUE_REG_11__2__SCAN_IN); 
assign P3_U4540 = ~(P3_U2484 & P3_INSTQUEUE_REG_0__3__SCAN_IN); 
assign P3_U4543 = ~(P3_U2480 & P3_INSTQUEUE_REG_3__3__SCAN_IN); 
assign P3_U4547 = ~(P3_U4471 & P3_INSTQUEUE_REG_7__3__SCAN_IN); 
assign P3_U4548 = ~(P3_U2476 & P3_INSTQUEUE_REG_8__3__SCAN_IN); 
assign P3_U4551 = ~(P3_U2471 & P3_INSTQUEUE_REG_11__3__SCAN_IN); 
assign P3_U4557 = ~(P3_U2484 & P3_INSTQUEUE_REG_0__7__SCAN_IN); 
assign P3_U4560 = ~(P3_U2480 & P3_INSTQUEUE_REG_3__7__SCAN_IN); 
assign P3_U4564 = ~(P3_U4471 & P3_INSTQUEUE_REG_7__7__SCAN_IN); 
assign P3_U4565 = ~(P3_U2476 & P3_INSTQUEUE_REG_8__7__SCAN_IN); 
assign P3_U4568 = ~(P3_U2471 & P3_INSTQUEUE_REG_11__7__SCAN_IN); 
assign P3_U4574 = ~(P3_U2484 & P3_INSTQUEUE_REG_0__5__SCAN_IN); 
assign P3_U4577 = ~(P3_U2480 & P3_INSTQUEUE_REG_3__5__SCAN_IN); 
assign P3_U4581 = ~(P3_U4471 & P3_INSTQUEUE_REG_7__5__SCAN_IN); 
assign P3_U4582 = ~(P3_U2476 & P3_INSTQUEUE_REG_8__5__SCAN_IN); 
assign P3_U4585 = ~(P3_U2471 & P3_INSTQUEUE_REG_11__5__SCAN_IN); 
assign P3_U4591 = ~(P3_U2484 & P3_INSTQUEUE_REG_0__6__SCAN_IN); 
assign P3_U4594 = ~(P3_U2480 & P3_INSTQUEUE_REG_3__6__SCAN_IN); 
assign P3_U4598 = ~(P3_U4471 & P3_INSTQUEUE_REG_7__6__SCAN_IN); 
assign P3_U4599 = ~(P3_U2476 & P3_INSTQUEUE_REG_8__6__SCAN_IN); 
assign P3_U4602 = ~(P3_U2471 & P3_INSTQUEUE_REG_11__6__SCAN_IN); 
assign P3_U4650 = ~P3_U3180; 
assign P3_U4654 = ~(P3_U4653 & P3_U3269); 
assign P3_U4662 = ~P3_U3134; 
assign P3_U4671 = ~(P3_U3134 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U5082 = ~(P3_U3180 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U5543 = ~P3_U3265; 
assign P3_U5544 = ~(P3_U4345 & P3_U3265); 
assign P3_U5554 = ~(P3_U3286 & P3_U3287 & P3_STATE2_REG_1__SCAN_IN); 
assign P3_U7516 = ~P3_U3266; 
assign P3_U7776 = ~(P3_U2600 & P3_INSTQUEUE_REG_8__7__SCAN_IN); 
assign P3_U7777 = ~(P3_U2599 & P3_INSTQUEUE_REG_9__7__SCAN_IN); 
assign P3_U7778 = ~(P3_U2598 & P3_INSTQUEUE_REG_10__7__SCAN_IN); 
assign P3_U7779 = ~(P3_U2597 & P3_INSTQUEUE_REG_11__7__SCAN_IN); 
assign P3_U7780 = ~(P3_U2595 & P3_INSTQUEUE_REG_12__7__SCAN_IN); 
assign P3_U7783 = ~(P3_U2592 & P3_INSTQUEUE_REG_15__7__SCAN_IN); 
assign P3_U7788 = ~(P3_U2586 & P3_INSTQUEUE_REG_4__7__SCAN_IN); 
assign P3_U7789 = ~(P3_U2585 & P3_INSTQUEUE_REG_5__7__SCAN_IN); 
assign P3_U7790 = ~(P3_U2584 & P3_INSTQUEUE_REG_6__7__SCAN_IN); 
assign P3_U7791 = ~(P3_U2583 & P3_INSTQUEUE_REG_7__7__SCAN_IN); 
assign P3_U7792 = ~(P3_U2600 & P3_INSTQUEUE_REG_8__6__SCAN_IN); 
assign P3_U7793 = ~(P3_U2599 & P3_INSTQUEUE_REG_9__6__SCAN_IN); 
assign P3_U7794 = ~(P3_U2598 & P3_INSTQUEUE_REG_10__6__SCAN_IN); 
assign P3_U7795 = ~(P3_U2597 & P3_INSTQUEUE_REG_11__6__SCAN_IN); 
assign P3_U7796 = ~(P3_U2595 & P3_INSTQUEUE_REG_12__6__SCAN_IN); 
assign P3_U7799 = ~(P3_U2592 & P3_INSTQUEUE_REG_15__6__SCAN_IN); 
assign P3_U7804 = ~(P3_U2586 & P3_INSTQUEUE_REG_4__6__SCAN_IN); 
assign P3_U7805 = ~(P3_U2585 & P3_INSTQUEUE_REG_5__6__SCAN_IN); 
assign P3_U7806 = ~(P3_U2584 & P3_INSTQUEUE_REG_6__6__SCAN_IN); 
assign P3_U7807 = ~(P3_U2583 & P3_INSTQUEUE_REG_7__6__SCAN_IN); 
assign P3_U7808 = ~(P3_U2600 & P3_INSTQUEUE_REG_8__5__SCAN_IN); 
assign P3_U7809 = ~(P3_U2599 & P3_INSTQUEUE_REG_9__5__SCAN_IN); 
assign P3_U7810 = ~(P3_U2598 & P3_INSTQUEUE_REG_10__5__SCAN_IN); 
assign P3_U7811 = ~(P3_U2597 & P3_INSTQUEUE_REG_11__5__SCAN_IN); 
assign P3_U7812 = ~(P3_U2595 & P3_INSTQUEUE_REG_12__5__SCAN_IN); 
assign P3_U7815 = ~(P3_U2592 & P3_INSTQUEUE_REG_15__5__SCAN_IN); 
assign P3_U7820 = ~(P3_U2586 & P3_INSTQUEUE_REG_4__5__SCAN_IN); 
assign P3_U7821 = ~(P3_U2585 & P3_INSTQUEUE_REG_5__5__SCAN_IN); 
assign P3_U7822 = ~(P3_U2584 & P3_INSTQUEUE_REG_6__5__SCAN_IN); 
assign P3_U7823 = ~(P3_U2583 & P3_INSTQUEUE_REG_7__5__SCAN_IN); 
assign P3_U7824 = ~(P3_U2600 & P3_INSTQUEUE_REG_8__4__SCAN_IN); 
assign P3_U7825 = ~(P3_U2599 & P3_INSTQUEUE_REG_9__4__SCAN_IN); 
assign P3_U7826 = ~(P3_U2598 & P3_INSTQUEUE_REG_10__4__SCAN_IN); 
assign P3_U7827 = ~(P3_U2597 & P3_INSTQUEUE_REG_11__4__SCAN_IN); 
assign P3_U7828 = ~(P3_U2595 & P3_INSTQUEUE_REG_12__4__SCAN_IN); 
assign P3_U7831 = ~(P3_U2592 & P3_INSTQUEUE_REG_15__4__SCAN_IN); 
assign P3_U7836 = ~(P3_U2586 & P3_INSTQUEUE_REG_4__4__SCAN_IN); 
assign P3_U7837 = ~(P3_U2585 & P3_INSTQUEUE_REG_5__4__SCAN_IN); 
assign P3_U7838 = ~(P3_U2584 & P3_INSTQUEUE_REG_6__4__SCAN_IN); 
assign P3_U7839 = ~(P3_U2583 & P3_INSTQUEUE_REG_7__4__SCAN_IN); 
assign P3_U7840 = ~(P3_U2600 & P3_INSTQUEUE_REG_8__3__SCAN_IN); 
assign P3_U7841 = ~(P3_U2599 & P3_INSTQUEUE_REG_9__3__SCAN_IN); 
assign P3_U7842 = ~(P3_U2598 & P3_INSTQUEUE_REG_10__3__SCAN_IN); 
assign P3_U7843 = ~(P3_U2597 & P3_INSTQUEUE_REG_11__3__SCAN_IN); 
assign P3_U7844 = ~(P3_U2595 & P3_INSTQUEUE_REG_12__3__SCAN_IN); 
assign P3_U7847 = ~(P3_U2592 & P3_INSTQUEUE_REG_15__3__SCAN_IN); 
assign P3_U7852 = ~(P3_U2586 & P3_INSTQUEUE_REG_4__3__SCAN_IN); 
assign P3_U7853 = ~(P3_U2585 & P3_INSTQUEUE_REG_5__3__SCAN_IN); 
assign P3_U7854 = ~(P3_U2584 & P3_INSTQUEUE_REG_6__3__SCAN_IN); 
assign P3_U7855 = ~(P3_U2583 & P3_INSTQUEUE_REG_7__3__SCAN_IN); 
assign P3_U7856 = ~(P3_U2600 & P3_INSTQUEUE_REG_8__2__SCAN_IN); 
assign P3_U7857 = ~(P3_U2599 & P3_INSTQUEUE_REG_9__2__SCAN_IN); 
assign P3_U7858 = ~(P3_U2598 & P3_INSTQUEUE_REG_10__2__SCAN_IN); 
assign P3_U7859 = ~(P3_U2597 & P3_INSTQUEUE_REG_11__2__SCAN_IN); 
assign P3_U7860 = ~(P3_U2595 & P3_INSTQUEUE_REG_12__2__SCAN_IN); 
assign P3_U7863 = ~(P3_U2592 & P3_INSTQUEUE_REG_15__2__SCAN_IN); 
assign P3_U7868 = ~(P3_U2586 & P3_INSTQUEUE_REG_4__2__SCAN_IN); 
assign P3_U7869 = ~(P3_U2585 & P3_INSTQUEUE_REG_5__2__SCAN_IN); 
assign P3_U7870 = ~(P3_U2584 & P3_INSTQUEUE_REG_6__2__SCAN_IN); 
assign P3_U7871 = ~(P3_U2583 & P3_INSTQUEUE_REG_7__2__SCAN_IN); 
assign P3_U7872 = ~(P3_U2600 & P3_INSTQUEUE_REG_8__1__SCAN_IN); 
assign P3_U7873 = ~(P3_U2599 & P3_INSTQUEUE_REG_9__1__SCAN_IN); 
assign P3_U7874 = ~(P3_U2598 & P3_INSTQUEUE_REG_10__1__SCAN_IN); 
assign P3_U7875 = ~(P3_U2597 & P3_INSTQUEUE_REG_11__1__SCAN_IN); 
assign P3_U7876 = ~(P3_U2595 & P3_INSTQUEUE_REG_12__1__SCAN_IN); 
assign P3_U7879 = ~(P3_U2592 & P3_INSTQUEUE_REG_15__1__SCAN_IN); 
assign P3_U7884 = ~(P3_U2586 & P3_INSTQUEUE_REG_4__1__SCAN_IN); 
assign P3_U7885 = ~(P3_U2585 & P3_INSTQUEUE_REG_5__1__SCAN_IN); 
assign P3_U7886 = ~(P3_U2584 & P3_INSTQUEUE_REG_6__1__SCAN_IN); 
assign P3_U7887 = ~(P3_U2583 & P3_INSTQUEUE_REG_7__1__SCAN_IN); 
assign P3_U7888 = ~(P3_U2600 & P3_INSTQUEUE_REG_8__0__SCAN_IN); 
assign P3_U7889 = ~(P3_U2599 & P3_INSTQUEUE_REG_9__0__SCAN_IN); 
assign P3_U7890 = ~(P3_U2598 & P3_INSTQUEUE_REG_10__0__SCAN_IN); 
assign P3_U7891 = ~(P3_U2597 & P3_INSTQUEUE_REG_11__0__SCAN_IN); 
assign P3_U7892 = ~(P3_U2595 & P3_INSTQUEUE_REG_12__0__SCAN_IN); 
assign P3_U7895 = ~(P3_U2592 & P3_INSTQUEUE_REG_15__0__SCAN_IN); 
assign P3_U7900 = ~(P3_U2586 & P3_INSTQUEUE_REG_4__0__SCAN_IN); 
assign P3_U7901 = ~(P3_U2585 & P3_INSTQUEUE_REG_5__0__SCAN_IN); 
assign P3_U7902 = ~(P3_U2584 & P3_INSTQUEUE_REG_6__0__SCAN_IN); 
assign P3_U7903 = ~(P3_U2583 & P3_INSTQUEUE_REG_7__0__SCAN_IN); 
assign P3_U7931 = ~(P3_U7914 & P3_U4449 & P3_STATE_REG_1__SCAN_IN); 
assign P3_U7932 = ~(P3_U7930 & P3_U3076); 
assign P3_U7937 = ~P3_U3278; 
assign P3_U7939 = ~(P3_U3279 & P3_U3278); 
assign P3_U7940 = ~(P3_U3278 & P3_U4464); 
assign P3_U7963 = ~(P3_U7962 & P3_U4653); 
assign P3_U7985 = ~P3_U3287; 
assign P3_U8011 = ~(P3_U8009 & P3_U4307); 
assign P3_U8021 = ~(BS16 & P3_U3278); 
assign P3_U8037 = ~P3_U3273; 
assign P3_U8039 = ~(P3_U3287 & P3_U3286 & P3_FLUSH_REG_SCAN_IN); 
assign P2_U2359 = P2_U4411 & P2_U3265; 
assign P2_U2441 = P2_U4647 & P2_U3580; 
assign P2_U2442 = P2_U8067 & P2_U3428; 
assign P2_U2443 = P2_U4647 & P2_U8067; 
assign P2_U2515 = P2_U8082 & P2_U8100; 
assign P2_U2520 = P2_U8082 & P2_U3582; 
assign P2_U2530 = P2_U2525 & P2_U2529; 
assign P2_U2531 = P2_U2523 & P2_U2529; 
assign P2_U2533 = P2_U2525 & P2_U2532; 
assign P2_U2534 = P2_U2523 & P2_U2532; 
assign P2_U2535 = P2_U2529 & P2_U2518; 
assign P2_U2536 = P2_U2529 & P2_U2516; 
assign P2_U2537 = P2_U2518 & P2_U2532; 
assign P2_U2538 = P2_U2516 & P2_U2532; 
assign P2_U2541 = P2_U2539 & P2_U2540; 
assign P2_U2543 = P2_U2539 & P2_U2542; 
assign P2_U2544 = P2_R2147_U4 & P2_U3526; 
assign P2_U2548 = P2_U2539 & P2_U2547; 
assign P2_U2550 = P2_U2539 & P2_U2549; 
assign P2_U2554 = P2_U2540 & P2_U2553; 
assign P2_U2555 = P2_U2542 & P2_U2553; 
assign P2_U2557 = P2_U2540 & P2_U2556; 
assign P2_U2558 = P2_U2542 & P2_U2556; 
assign P2_U2559 = P2_U2553 & P2_U2547; 
assign P2_U2560 = P2_U2553 & P2_U2549; 
assign P2_U2561 = P2_U2547 & P2_U2556; 
assign P2_U2562 = P2_U2549 & P2_U2556; 
assign P2_U2564 = P2_U4409 & P2_U3583; 
assign P2_U2572 = P2_U3583 & P2_U3553; 
assign P2_U2616 = ~(P2_U3706 & P2_U3705); 
assign P2_U2617 = ~(P2_U3694 & P2_U3693); 
assign P2_U2820 = ~(P2_U8128 & P2_U8127 & P2_U3548); 
assign P2_U2821 = ~(P2_U3548 & P2_U4452 & P2_U6837); 
assign P2_U2823 = ~(P2_U8124 & P2_U8123 & P2_U4452); 
assign P2_U3245 = ~(P2_U2440 & P2_U3243); 
assign P2_U3246 = ~(P2_U2440 & P2_U4650); 
assign P2_U3253 = ~(P2_U3708 & P2_U3707); 
assign P2_U3255 = ~(P2_U3696 & P2_U3695); 
assign P2_U3278 = ~(P2_U3700 & P2_U3699); 
assign P2_U3279 = ~(P2_U3702 & P2_U3701); 
assign P2_U3280 = ~(P2_U3704 & P2_U3703); 
assign P2_U3521 = ~(P2_U3698 & P2_U3697); 
assign P2_U3658 = ~(P2_U8372 & P2_U8371); 
assign P2_U3660 = ~(P2_U8376 & P2_U8375); 
assign P2_U3690 = P2_U4578 & P2_U3261; 
assign P2_U4069 = P2_U4454 & P2_U4453 & P2_U6569; 
assign P2_U4398 = P2_U8126 & P2_U8125; 
assign P2_U4477 = ~P2_U3548; 
assign P2_U4478 = ~(P2_U4450 & P2_REIP_REG_31__SCAN_IN); 
assign P2_U4479 = ~(P2_U4449 & P2_REIP_REG_30__SCAN_IN); 
assign P2_U4481 = ~(P2_U4450 & P2_REIP_REG_30__SCAN_IN); 
assign P2_U4482 = ~(P2_U4449 & P2_REIP_REG_29__SCAN_IN); 
assign P2_U4484 = ~(P2_U4450 & P2_REIP_REG_29__SCAN_IN); 
assign P2_U4485 = ~(P2_U4449 & P2_REIP_REG_28__SCAN_IN); 
assign P2_U4487 = ~(P2_U4450 & P2_REIP_REG_28__SCAN_IN); 
assign P2_U4488 = ~(P2_U4449 & P2_REIP_REG_27__SCAN_IN); 
assign P2_U4490 = ~(P2_U4450 & P2_REIP_REG_27__SCAN_IN); 
assign P2_U4491 = ~(P2_U4449 & P2_REIP_REG_26__SCAN_IN); 
assign P2_U4493 = ~(P2_U4450 & P2_REIP_REG_26__SCAN_IN); 
assign P2_U4494 = ~(P2_U4449 & P2_REIP_REG_25__SCAN_IN); 
assign P2_U4496 = ~(P2_U4450 & P2_REIP_REG_25__SCAN_IN); 
assign P2_U4497 = ~(P2_U4449 & P2_REIP_REG_24__SCAN_IN); 
assign P2_U4499 = ~(P2_U4450 & P2_REIP_REG_24__SCAN_IN); 
assign P2_U4500 = ~(P2_U4449 & P2_REIP_REG_23__SCAN_IN); 
assign P2_U4502 = ~(P2_U4450 & P2_REIP_REG_23__SCAN_IN); 
assign P2_U4503 = ~(P2_U4449 & P2_REIP_REG_22__SCAN_IN); 
assign P2_U4505 = ~(P2_U4450 & P2_REIP_REG_22__SCAN_IN); 
assign P2_U4506 = ~(P2_U4449 & P2_REIP_REG_21__SCAN_IN); 
assign P2_U4508 = ~(P2_U4450 & P2_REIP_REG_21__SCAN_IN); 
assign P2_U4509 = ~(P2_U4449 & P2_REIP_REG_20__SCAN_IN); 
assign P2_U4511 = ~(P2_U4450 & P2_REIP_REG_20__SCAN_IN); 
assign P2_U4512 = ~(P2_U4449 & P2_REIP_REG_19__SCAN_IN); 
assign P2_U4514 = ~(P2_U4450 & P2_REIP_REG_19__SCAN_IN); 
assign P2_U4515 = ~(P2_U4449 & P2_REIP_REG_18__SCAN_IN); 
assign P2_U4517 = ~(P2_U4450 & P2_REIP_REG_18__SCAN_IN); 
assign P2_U4518 = ~(P2_U4449 & P2_REIP_REG_17__SCAN_IN); 
assign P2_U4520 = ~(P2_U4450 & P2_REIP_REG_17__SCAN_IN); 
assign P2_U4521 = ~(P2_U4449 & P2_REIP_REG_16__SCAN_IN); 
assign P2_U4523 = ~(P2_U4450 & P2_REIP_REG_16__SCAN_IN); 
assign P2_U4524 = ~(P2_U4449 & P2_REIP_REG_15__SCAN_IN); 
assign P2_U4526 = ~(P2_U4450 & P2_REIP_REG_15__SCAN_IN); 
assign P2_U4527 = ~(P2_U4449 & P2_REIP_REG_14__SCAN_IN); 
assign P2_U4529 = ~(P2_U4450 & P2_REIP_REG_14__SCAN_IN); 
assign P2_U4530 = ~(P2_U4449 & P2_REIP_REG_13__SCAN_IN); 
assign P2_U4532 = ~(P2_U4450 & P2_REIP_REG_13__SCAN_IN); 
assign P2_U4533 = ~(P2_U4449 & P2_REIP_REG_12__SCAN_IN); 
assign P2_U4535 = ~(P2_U4450 & P2_REIP_REG_12__SCAN_IN); 
assign P2_U4536 = ~(P2_U4449 & P2_REIP_REG_11__SCAN_IN); 
assign P2_U4538 = ~(P2_U4450 & P2_REIP_REG_11__SCAN_IN); 
assign P2_U4539 = ~(P2_U4449 & P2_REIP_REG_10__SCAN_IN); 
assign P2_U4541 = ~(P2_U4450 & P2_REIP_REG_10__SCAN_IN); 
assign P2_U4542 = ~(P2_U4449 & P2_REIP_REG_9__SCAN_IN); 
assign P2_U4544 = ~(P2_U4450 & P2_REIP_REG_9__SCAN_IN); 
assign P2_U4545 = ~(P2_U4449 & P2_REIP_REG_8__SCAN_IN); 
assign P2_U4547 = ~(P2_U4450 & P2_REIP_REG_8__SCAN_IN); 
assign P2_U4548 = ~(P2_U4449 & P2_REIP_REG_7__SCAN_IN); 
assign P2_U4550 = ~(P2_U4450 & P2_REIP_REG_7__SCAN_IN); 
assign P2_U4551 = ~(P2_U4449 & P2_REIP_REG_6__SCAN_IN); 
assign P2_U4553 = ~(P2_U4450 & P2_REIP_REG_6__SCAN_IN); 
assign P2_U4554 = ~(P2_U4449 & P2_REIP_REG_5__SCAN_IN); 
assign P2_U4556 = ~(P2_U4450 & P2_REIP_REG_5__SCAN_IN); 
assign P2_U4557 = ~(P2_U4449 & P2_REIP_REG_4__SCAN_IN); 
assign P2_U4559 = ~(P2_U4450 & P2_REIP_REG_4__SCAN_IN); 
assign P2_U4560 = ~(P2_U4449 & P2_REIP_REG_3__SCAN_IN); 
assign P2_U4562 = ~(P2_U4450 & P2_REIP_REG_3__SCAN_IN); 
assign P2_U4563 = ~(P2_U4449 & P2_REIP_REG_2__SCAN_IN); 
assign P2_U4565 = ~(P2_U4450 & P2_REIP_REG_2__SCAN_IN); 
assign P2_U4566 = ~(P2_U4449 & P2_REIP_REG_1__SCAN_IN); 
assign P2_U4573 = ~(P2_U4392 & P2_U7891); 
assign P2_U4584 = ~(P2_U3692 & P2_U7893); 
assign P2_U4624 = ~(P2_U4623 & P2_STATE2_REG_1__SCAN_IN); 
assign P2_U4651 = ~(P2_U2440 & P2_U2444); 
assign P2_U4770 = ~(P2_U2445 & P2_U2440); 
assign P2_U6844 = ~(P2_U4411 & P2_STATEBS16_REG_SCAN_IN); 
assign P2_U6847 = ~(P2_U4411 & P2_U3265); 
assign P2_U7754 = ~(P2_U8154 & P2_U8153 & P2_U4592); 
assign P2_U7755 = ~(P2_U8170 & P2_U8169 & P2_U4592); 
assign P2_U7756 = ~(P2_U8186 & P2_U8185 & P2_U4592); 
assign P2_U7757 = ~(P2_U8202 & P2_U8201 & P2_U4592); 
assign P2_U7758 = ~(P2_U8218 & P2_U8217 & P2_U4592); 
assign P2_U7759 = ~(P2_U8234 & P2_U8233 & P2_U4592); 
assign P2_U7760 = ~(P2_U8250 & P2_U8249 & P2_U4592); 
assign P2_U7761 = ~(P2_U8266 & P2_U8265 & P2_U4592); 
assign P2_U7770 = ~(P2_U8156 & P2_U8155 & P2_U4593); 
assign P2_U7771 = ~(P2_U8172 & P2_U8171 & P2_U4593); 
assign P2_U7772 = ~(P2_U8188 & P2_U8187 & P2_U4593); 
assign P2_U7773 = ~(P2_U8204 & P2_U8203 & P2_U4593); 
assign P2_U7774 = ~(P2_U8220 & P2_U8219 & P2_U4593); 
assign P2_U7775 = ~(P2_U8236 & P2_U8235 & P2_U4593); 
assign P2_U7776 = ~(P2_U8252 & P2_U8251 & P2_U4593); 
assign P2_U7777 = ~(P2_U8268 & P2_U8267 & P2_U4593); 
assign P2_U7786 = ~(P2_U8158 & P2_U8157 & P2_U2456); 
assign P2_U7787 = ~(P2_U8174 & P2_U8173 & P2_U2456); 
assign P2_U7788 = ~(P2_U8190 & P2_U8189 & P2_U2456); 
assign P2_U7789 = ~(P2_U8206 & P2_U8205 & P2_U2456); 
assign P2_U7790 = ~(P2_U8222 & P2_U8221 & P2_U2456); 
assign P2_U7791 = ~(P2_U8238 & P2_U8237 & P2_U2456); 
assign P2_U7792 = ~(P2_U8254 & P2_U8253 & P2_U2456); 
assign P2_U7793 = ~(P2_U8270 & P2_U8269 & P2_U2456); 
assign P2_U7802 = ~(P2_U8160 & P2_U8159 & P2_U2454); 
assign P2_U7803 = ~(P2_U8176 & P2_U8175 & P2_U2454); 
assign P2_U7804 = ~(P2_U8192 & P2_U8191 & P2_U2454); 
assign P2_U7805 = ~(P2_U8208 & P2_U8207 & P2_U2454); 
assign P2_U7806 = ~(P2_U8224 & P2_U8223 & P2_U2454); 
assign P2_U7807 = ~(P2_U8240 & P2_U8239 & P2_U2454); 
assign P2_U7808 = ~(P2_U8256 & P2_U8255 & P2_U2454); 
assign P2_U7809 = ~(P2_U8272 & P2_U8271 & P2_U2454); 
assign P2_U7818 = ~(P2_U8162 & P2_U8161 & P2_U4590); 
assign P2_U7819 = ~(P2_U8178 & P2_U8177 & P2_U4590); 
assign P2_U7820 = ~(P2_U8194 & P2_U8193 & P2_U4590); 
assign P2_U7821 = ~(P2_U8210 & P2_U8209 & P2_U4590); 
assign P2_U7822 = ~(P2_U8226 & P2_U8225 & P2_U4590); 
assign P2_U7823 = ~(P2_U8242 & P2_U8241 & P2_U4590); 
assign P2_U7824 = ~(P2_U8258 & P2_U8257 & P2_U4590); 
assign P2_U7825 = ~(P2_U8274 & P2_U8273 & P2_U4590); 
assign P2_U7834 = ~(P2_U8164 & P2_U8163 & P2_U2453); 
assign P2_U7835 = ~(P2_U8180 & P2_U8179 & P2_U2453); 
assign P2_U7836 = ~(P2_U8196 & P2_U8195 & P2_U2453); 
assign P2_U7837 = ~(P2_U8212 & P2_U8211 & P2_U2453); 
assign P2_U7838 = ~(P2_U8228 & P2_U8227 & P2_U2453); 
assign P2_U7839 = ~(P2_U8244 & P2_U8243 & P2_U2453); 
assign P2_U7840 = ~(P2_U8260 & P2_U8259 & P2_U2453); 
assign P2_U7841 = ~(P2_U8276 & P2_U8275 & P2_U2453); 
assign P2_U7850 = ~(P2_U8166 & P2_U8165 & P2_U2452); 
assign P2_U7851 = ~(P2_U8182 & P2_U8181 & P2_U2452); 
assign P2_U7852 = ~(P2_U8198 & P2_U8197 & P2_U2452); 
assign P2_U7853 = ~(P2_U8214 & P2_U8213 & P2_U2452); 
assign P2_U7854 = ~(P2_U8230 & P2_U8229 & P2_U2452); 
assign P2_U7855 = ~(P2_U8246 & P2_U8245 & P2_U2452); 
assign P2_U7856 = ~(P2_U8262 & P2_U8261 & P2_U2452); 
assign P2_U7857 = ~(P2_U8278 & P2_U8277 & P2_U2452); 
assign P2_U7874 = ~(P2_U8168 & P2_U8167 & P2_U2455); 
assign P2_U7875 = ~(P2_U8184 & P2_U8183 & P2_U2455); 
assign P2_U7876 = ~(P2_U8200 & P2_U8199 & P2_U2455); 
assign P2_U7877 = ~(P2_U8216 & P2_U8215 & P2_U2455); 
assign P2_U7878 = ~(P2_U8232 & P2_U8231 & P2_U2455); 
assign P2_U7879 = ~(P2_U8248 & P2_U8247 & P2_U2455); 
assign P2_U7880 = ~(P2_U8264 & P2_U8263 & P2_U2455); 
assign P2_U7881 = ~(P2_U8280 & P2_U8279 & P2_U2455); 
assign P2_U7911 = ~(P2_U4581 & P2_U4572 & P2_STATE_REG_1__SCAN_IN); 
assign P2_U7912 = ~(P2_U4582 & P2_U3258); 
assign P2_U7917 = ~P2_U3589; 
assign P2_U7919 = ~(P2_U3590 & P2_U3589); 
assign P2_U7920 = ~(P2_U3589 & P2_U4589); 
assign P2_U8136 = ~(BS16 & P2_U3589); 
assign P2_U8149 = ~P2_U3583; 
assign P1_U2433 = P1_U4540 & P1_U3455; 
assign P1_U2434 = P1_U7696 & P1_U3360; 
assign P1_U2435 = P1_U4540 & P1_U7696; 
assign P1_U2450 = P1_U4400 & P1_STATE2_REG_0__SCAN_IN; 
assign P1_U2522 = P1_U5483 & P1_U5511; 
assign P1_U2530 = P1_U5483 & P1_U3401; 
assign P1_U2536 = P1_U2535 & P1_U2521; 
assign P1_U2537 = P1_U2535 & P1_U2524; 
assign P1_U2538 = P1_U2535 & P1_U2526; 
assign P1_U2539 = P1_U2535 & P1_U2528; 
assign P1_U2541 = P1_U2521 & P1_U2540; 
assign P1_U2542 = P1_U2524 & P1_U2540; 
assign P1_U2543 = P1_U2526 & P1_U2540; 
assign P1_U2544 = P1_U2528 & P1_U2540; 
assign P1_U2555 = P1_U7720 & P1_U3442; 
assign P1_U2560 = P1_U3456 & P1_U3442; 
assign P1_U2570 = P1_U2569 & P1_U3498; 
assign P1_U2571 = P1_U2569 & P1_U2454; 
assign P1_U2572 = P1_U2569 & P1_U2456; 
assign P1_U2573 = P1_U2569 & P1_U4378; 
assign P1_U2593 = P1_U4184 & P1_U3457; 
assign P1_U2598 = P1_U3457 & P1_U3452; 
assign P1_U2807 = ~(P1_U7757 & P1_U7756 & P1_U4240); 
assign P1_U2808 = ~(P1_U7747 & P1_U7746 & P1_U4240); 
assign P1_U3236 = ~(P1_U2432 & P1_U3235); 
assign P1_U3237 = ~(P1_U2432 & P1_U4543); 
assign P1_U3271 = ~(P1_U3567 & P1_U3566 & P1_U3565 & P1_U3564); 
assign P1_U3276 = ~(P1_U3519 & P1_U3518 & P1_U3517 & P1_U3516); 
assign P1_U3277 = ~(P1_U3539 & P1_U4170 & P1_U3538 & P1_U3537 & P1_U3536); 
assign P1_U3283 = ~(P1_U3511 & P1_U3510 & P1_U3509 & P1_U3508); 
assign P1_U3284 = ~(P1_U3563 & P1_U3562 & P1_U3561 & P1_U3560); 
assign P1_U3391 = ~(P1_U3515 & P1_U3514 & P1_U3513 & P1_U3512); 
assign P1_U3415 = ~(P1_U4400 & P1_U4173); 
assign P1_U3453 = ~(P1_U2605 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U3482 = ~(P1_U7759 & P1_U7758); 
assign P1_U3494 = P1_U4368 & P1_U3252; 
assign P1_U3733 = P1_U4497 & P1_U3257; 
assign P1_U4064 = P1_U7073 & P1_U7072 & P1_U7071 & P1_U7070; 
assign P1_U4078 = P1_U7097 & P1_U7095; 
assign P1_U4080 = P1_U7105 & P1_U7104 & P1_U7103 & P1_U7102; 
assign P1_U4084 = P1_U7122 & P1_U7121 & P1_U7120 & P1_U7119; 
assign P1_U4088 = P1_U7139 & P1_U7138 & P1_U7137 & P1_U7136; 
assign P1_U4093 = P1_U7154 & P1_U7153 & P1_U7152 & P1_U7151; 
assign P1_U4097 = P1_U7171 & P1_U7170 & P1_U7169 & P1_U7168; 
assign P1_U4101 = P1_U7188 & P1_U7187 & P1_U7186 & P1_U7185; 
assign P1_U4105 = P1_U7205 & P1_U7204 & P1_U7203 & P1_U7202; 
assign P1_U4109 = P1_U7216 & P1_U7215; 
assign P1_U4160 = P1_U4173 & P1_STATE2_REG_0__SCAN_IN; 
assign P1_U4171 = ~(P1_U3572 & P1_U3571 & P1_U3570 & P1_U3569); 
assign P1_U4267 = ~(P1_U4233 & P1_REIP_REG_31__SCAN_IN); 
assign P1_U4268 = ~(P1_U4232 & P1_REIP_REG_30__SCAN_IN); 
assign P1_U4270 = ~(P1_U4233 & P1_REIP_REG_30__SCAN_IN); 
assign P1_U4271 = ~(P1_U4232 & P1_REIP_REG_29__SCAN_IN); 
assign P1_U4273 = ~(P1_U4233 & P1_REIP_REG_29__SCAN_IN); 
assign P1_U4274 = ~(P1_U4232 & P1_REIP_REG_28__SCAN_IN); 
assign P1_U4276 = ~(P1_U4233 & P1_REIP_REG_28__SCAN_IN); 
assign P1_U4277 = ~(P1_U4232 & P1_REIP_REG_27__SCAN_IN); 
assign P1_U4279 = ~(P1_U4233 & P1_REIP_REG_27__SCAN_IN); 
assign P1_U4280 = ~(P1_U4232 & P1_REIP_REG_26__SCAN_IN); 
assign P1_U4282 = ~(P1_U4233 & P1_REIP_REG_26__SCAN_IN); 
assign P1_U4283 = ~(P1_U4232 & P1_REIP_REG_25__SCAN_IN); 
assign P1_U4285 = ~(P1_U4233 & P1_REIP_REG_25__SCAN_IN); 
assign P1_U4286 = ~(P1_U4232 & P1_REIP_REG_24__SCAN_IN); 
assign P1_U4288 = ~(P1_U4233 & P1_REIP_REG_24__SCAN_IN); 
assign P1_U4289 = ~(P1_U4232 & P1_REIP_REG_23__SCAN_IN); 
assign P1_U4291 = ~(P1_U4233 & P1_REIP_REG_23__SCAN_IN); 
assign P1_U4292 = ~(P1_U4232 & P1_REIP_REG_22__SCAN_IN); 
assign P1_U4294 = ~(P1_U4233 & P1_REIP_REG_22__SCAN_IN); 
assign P1_U4295 = ~(P1_U4232 & P1_REIP_REG_21__SCAN_IN); 
assign P1_U4297 = ~(P1_U4233 & P1_REIP_REG_21__SCAN_IN); 
assign P1_U4298 = ~(P1_U4232 & P1_REIP_REG_20__SCAN_IN); 
assign P1_U4300 = ~(P1_U4233 & P1_REIP_REG_20__SCAN_IN); 
assign P1_U4301 = ~(P1_U4232 & P1_REIP_REG_19__SCAN_IN); 
assign P1_U4303 = ~(P1_U4233 & P1_REIP_REG_19__SCAN_IN); 
assign P1_U4304 = ~(P1_U4232 & P1_REIP_REG_18__SCAN_IN); 
assign P1_U4306 = ~(P1_U4233 & P1_REIP_REG_18__SCAN_IN); 
assign P1_U4307 = ~(P1_U4232 & P1_REIP_REG_17__SCAN_IN); 
assign P1_U4309 = ~(P1_U4233 & P1_REIP_REG_17__SCAN_IN); 
assign P1_U4310 = ~(P1_U4232 & P1_REIP_REG_16__SCAN_IN); 
assign P1_U4312 = ~(P1_U4233 & P1_REIP_REG_16__SCAN_IN); 
assign P1_U4313 = ~(P1_U4232 & P1_REIP_REG_15__SCAN_IN); 
assign P1_U4315 = ~(P1_U4233 & P1_REIP_REG_15__SCAN_IN); 
assign P1_U4316 = ~(P1_U4232 & P1_REIP_REG_14__SCAN_IN); 
assign P1_U4318 = ~(P1_U4233 & P1_REIP_REG_14__SCAN_IN); 
assign P1_U4319 = ~(P1_U4232 & P1_REIP_REG_13__SCAN_IN); 
assign P1_U4321 = ~(P1_U4233 & P1_REIP_REG_13__SCAN_IN); 
assign P1_U4322 = ~(P1_U4232 & P1_REIP_REG_12__SCAN_IN); 
assign P1_U4324 = ~(P1_U4233 & P1_REIP_REG_12__SCAN_IN); 
assign P1_U4325 = ~(P1_U4232 & P1_REIP_REG_11__SCAN_IN); 
assign P1_U4327 = ~(P1_U4233 & P1_REIP_REG_11__SCAN_IN); 
assign P1_U4328 = ~(P1_U4232 & P1_REIP_REG_10__SCAN_IN); 
assign P1_U4330 = ~(P1_U4233 & P1_REIP_REG_10__SCAN_IN); 
assign P1_U4331 = ~(P1_U4232 & P1_REIP_REG_9__SCAN_IN); 
assign P1_U4333 = ~(P1_U4233 & P1_REIP_REG_9__SCAN_IN); 
assign P1_U4334 = ~(P1_U4232 & P1_REIP_REG_8__SCAN_IN); 
assign P1_U4336 = ~(P1_U4233 & P1_REIP_REG_8__SCAN_IN); 
assign P1_U4337 = ~(P1_U4232 & P1_REIP_REG_7__SCAN_IN); 
assign P1_U4339 = ~(P1_U4233 & P1_REIP_REG_7__SCAN_IN); 
assign P1_U4340 = ~(P1_U4232 & P1_REIP_REG_6__SCAN_IN); 
assign P1_U4342 = ~(P1_U4233 & P1_REIP_REG_6__SCAN_IN); 
assign P1_U4343 = ~(P1_U4232 & P1_REIP_REG_5__SCAN_IN); 
assign P1_U4345 = ~(P1_U4233 & P1_REIP_REG_5__SCAN_IN); 
assign P1_U4346 = ~(P1_U4232 & P1_REIP_REG_4__SCAN_IN); 
assign P1_U4348 = ~(P1_U4233 & P1_REIP_REG_4__SCAN_IN); 
assign P1_U4349 = ~(P1_U4232 & P1_REIP_REG_3__SCAN_IN); 
assign P1_U4351 = ~(P1_U4233 & P1_REIP_REG_3__SCAN_IN); 
assign P1_U4352 = ~(P1_U4232 & P1_REIP_REG_2__SCAN_IN); 
assign P1_U4354 = ~(P1_U4233 & P1_REIP_REG_2__SCAN_IN); 
assign P1_U4355 = ~(P1_U4232 & P1_REIP_REG_1__SCAN_IN); 
assign P1_U4363 = ~(P1_U7622 & P1_U4362 & P1_U7623); 
assign P1_U4371 = ~(P1_U3496 & P1_U7625); 
assign P1_U4415 = ~P1_U4173; 
assign P1_U4544 = ~(P1_U2432 & P1_U2436); 
assign P1_U4663 = ~(P1_U2437 & P1_U2432); 
assign P1_U5480 = ~P1_U3442; 
assign P1_U5488 = ~(P1_U4400 & P1_U2605); 
assign P1_U5515 = ~(P1_U2446 & P1_U3470); 
assign P1_U6604 = ~(P1_U4497 & P1_STATEBS16_REG_SCAN_IN); 
assign P1_U7066 = ~(P1_U2582 & P1_INSTQUEUE_REG_8__7__SCAN_IN); 
assign P1_U7067 = ~(P1_U2581 & P1_INSTQUEUE_REG_9__7__SCAN_IN); 
assign P1_U7068 = ~(P1_U2580 & P1_INSTQUEUE_REG_10__7__SCAN_IN); 
assign P1_U7069 = ~(P1_U2579 & P1_INSTQUEUE_REG_11__7__SCAN_IN); 
assign P1_U7078 = ~(P1_U2568 & P1_INSTQUEUE_REG_4__7__SCAN_IN); 
assign P1_U7079 = ~(P1_U2567 & P1_INSTQUEUE_REG_5__7__SCAN_IN); 
assign P1_U7080 = ~(P1_U2566 & P1_INSTQUEUE_REG_6__7__SCAN_IN); 
assign P1_U7081 = ~(P1_U2565 & P1_INSTQUEUE_REG_7__7__SCAN_IN); 
assign P1_U7098 = ~(P1_U2582 & P1_INSTQUEUE_REG_8__6__SCAN_IN); 
assign P1_U7099 = ~(P1_U2581 & P1_INSTQUEUE_REG_9__6__SCAN_IN); 
assign P1_U7100 = ~(P1_U2580 & P1_INSTQUEUE_REG_10__6__SCAN_IN); 
assign P1_U7101 = ~(P1_U2579 & P1_INSTQUEUE_REG_11__6__SCAN_IN); 
assign P1_U7110 = ~(P1_U2568 & P1_INSTQUEUE_REG_4__6__SCAN_IN); 
assign P1_U7111 = ~(P1_U2567 & P1_INSTQUEUE_REG_5__6__SCAN_IN); 
assign P1_U7112 = ~(P1_U2566 & P1_INSTQUEUE_REG_6__6__SCAN_IN); 
assign P1_U7113 = ~(P1_U2565 & P1_INSTQUEUE_REG_7__6__SCAN_IN); 
assign P1_U7115 = ~(P1_U2582 & P1_INSTQUEUE_REG_8__5__SCAN_IN); 
assign P1_U7116 = ~(P1_U2581 & P1_INSTQUEUE_REG_9__5__SCAN_IN); 
assign P1_U7117 = ~(P1_U2580 & P1_INSTQUEUE_REG_10__5__SCAN_IN); 
assign P1_U7118 = ~(P1_U2579 & P1_INSTQUEUE_REG_11__5__SCAN_IN); 
assign P1_U7127 = ~(P1_U2568 & P1_INSTQUEUE_REG_4__5__SCAN_IN); 
assign P1_U7128 = ~(P1_U2567 & P1_INSTQUEUE_REG_5__5__SCAN_IN); 
assign P1_U7129 = ~(P1_U2566 & P1_INSTQUEUE_REG_6__5__SCAN_IN); 
assign P1_U7130 = ~(P1_U2565 & P1_INSTQUEUE_REG_7__5__SCAN_IN); 
assign P1_U7132 = ~(P1_U2582 & P1_INSTQUEUE_REG_8__4__SCAN_IN); 
assign P1_U7133 = ~(P1_U2581 & P1_INSTQUEUE_REG_9__4__SCAN_IN); 
assign P1_U7134 = ~(P1_U2580 & P1_INSTQUEUE_REG_10__4__SCAN_IN); 
assign P1_U7135 = ~(P1_U2579 & P1_INSTQUEUE_REG_11__4__SCAN_IN); 
assign P1_U7143 = ~(P1_U2568 & P1_INSTQUEUE_REG_4__4__SCAN_IN); 
assign P1_U7144 = ~(P1_U2567 & P1_INSTQUEUE_REG_5__4__SCAN_IN); 
assign P1_U7145 = ~(P1_U2566 & P1_INSTQUEUE_REG_6__4__SCAN_IN); 
assign P1_U7146 = ~(P1_U2565 & P1_INSTQUEUE_REG_7__4__SCAN_IN); 
assign P1_U7147 = ~(P1_U2582 & P1_INSTQUEUE_REG_8__3__SCAN_IN); 
assign P1_U7148 = ~(P1_U2581 & P1_INSTQUEUE_REG_9__3__SCAN_IN); 
assign P1_U7149 = ~(P1_U2580 & P1_INSTQUEUE_REG_10__3__SCAN_IN); 
assign P1_U7150 = ~(P1_U2579 & P1_INSTQUEUE_REG_11__3__SCAN_IN); 
assign P1_U7159 = ~(P1_U2568 & P1_INSTQUEUE_REG_4__3__SCAN_IN); 
assign P1_U7160 = ~(P1_U2567 & P1_INSTQUEUE_REG_5__3__SCAN_IN); 
assign P1_U7161 = ~(P1_U2566 & P1_INSTQUEUE_REG_6__3__SCAN_IN); 
assign P1_U7162 = ~(P1_U2565 & P1_INSTQUEUE_REG_7__3__SCAN_IN); 
assign P1_U7164 = ~(P1_U2582 & P1_INSTQUEUE_REG_8__2__SCAN_IN); 
assign P1_U7165 = ~(P1_U2581 & P1_INSTQUEUE_REG_9__2__SCAN_IN); 
assign P1_U7166 = ~(P1_U2580 & P1_INSTQUEUE_REG_10__2__SCAN_IN); 
assign P1_U7167 = ~(P1_U2579 & P1_INSTQUEUE_REG_11__2__SCAN_IN); 
assign P1_U7176 = ~(P1_U2568 & P1_INSTQUEUE_REG_4__2__SCAN_IN); 
assign P1_U7177 = ~(P1_U2567 & P1_INSTQUEUE_REG_5__2__SCAN_IN); 
assign P1_U7178 = ~(P1_U2566 & P1_INSTQUEUE_REG_6__2__SCAN_IN); 
assign P1_U7179 = ~(P1_U2565 & P1_INSTQUEUE_REG_7__2__SCAN_IN); 
assign P1_U7181 = ~(P1_U2582 & P1_INSTQUEUE_REG_8__1__SCAN_IN); 
assign P1_U7182 = ~(P1_U2581 & P1_INSTQUEUE_REG_9__1__SCAN_IN); 
assign P1_U7183 = ~(P1_U2580 & P1_INSTQUEUE_REG_10__1__SCAN_IN); 
assign P1_U7184 = ~(P1_U2579 & P1_INSTQUEUE_REG_11__1__SCAN_IN); 
assign P1_U7193 = ~(P1_U2568 & P1_INSTQUEUE_REG_4__1__SCAN_IN); 
assign P1_U7194 = ~(P1_U2567 & P1_INSTQUEUE_REG_5__1__SCAN_IN); 
assign P1_U7195 = ~(P1_U2566 & P1_INSTQUEUE_REG_6__1__SCAN_IN); 
assign P1_U7196 = ~(P1_U2565 & P1_INSTQUEUE_REG_7__1__SCAN_IN); 
assign P1_U7198 = ~(P1_U2582 & P1_INSTQUEUE_REG_8__0__SCAN_IN); 
assign P1_U7199 = ~(P1_U2581 & P1_INSTQUEUE_REG_9__0__SCAN_IN); 
assign P1_U7200 = ~(P1_U2580 & P1_INSTQUEUE_REG_10__0__SCAN_IN); 
assign P1_U7201 = ~(P1_U2579 & P1_INSTQUEUE_REG_11__0__SCAN_IN); 
assign P1_U7210 = ~(P1_U2568 & P1_INSTQUEUE_REG_4__0__SCAN_IN); 
assign P1_U7211 = ~(P1_U2567 & P1_INSTQUEUE_REG_5__0__SCAN_IN); 
assign P1_U7212 = ~(P1_U2566 & P1_INSTQUEUE_REG_6__0__SCAN_IN); 
assign P1_U7213 = ~(P1_U2565 & P1_INSTQUEUE_REG_7__0__SCAN_IN); 
assign P1_U7380 = ~(P1_U4173 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U7461 = ~(P1_U2446 & P1_U3470 & P1_FLUSH_REG_SCAN_IN); 
assign P1_U7478 = ~(P1_U2608 & P1_U3266); 
assign P1_U7491 = ~(P1_U4108 & P1_U7216); 
assign P1_U7644 = ~(P1_U7624 & P1_U4361 & P1_STATE_REG_1__SCAN_IN); 
assign P1_U7645 = ~(P1_U7643 & P1_U3248); 
assign P1_U7650 = ~P1_U3462; 
assign P1_U7652 = ~(P1_U3463 & P1_U3462); 
assign P1_U7653 = ~(P1_U3462 & P1_U4376); 
assign P1_U7712 = ~P1_U3470; 
assign P1_U7755 = ~(P1_U7753 & P1_U4220); 
assign P1_U7765 = ~(BS16 & P1_U3462); 
assign P1_U7790 = ~P1_U3457; 
assign P3_ADD_526_U55 = ~(P3_ADD_526_U150 & P3_ADD_526_U149); 
assign P3_ADD_526_U56 = ~(P3_ADD_526_U152 & P3_ADD_526_U151); 
assign P3_ADD_526_U118 = ~P3_ADD_526_U16; 
assign P3_ADD_526_U126 = ~P3_ADD_526_U96; 
assign P3_ADD_526_U146 = ~(P3_ADD_526_U16 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_526_U147 = ~(P3_ADD_526_U96 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_552_U55 = ~(P3_ADD_552_U150 & P3_ADD_552_U149); 
assign P3_ADD_552_U56 = ~(P3_ADD_552_U152 & P3_ADD_552_U151); 
assign P3_ADD_552_U118 = ~P3_ADD_552_U16; 
assign P3_ADD_552_U126 = ~P3_ADD_552_U96; 
assign P3_ADD_552_U146 = ~(P3_ADD_552_U16 & P3_EBX_REG_7__SCAN_IN); 
assign P3_ADD_552_U147 = ~(P3_ADD_552_U96 & P3_EBX_REG_6__SCAN_IN); 
assign P3_ADD_546_U55 = ~(P3_ADD_546_U150 & P3_ADD_546_U149); 
assign P3_ADD_546_U56 = ~(P3_ADD_546_U152 & P3_ADD_546_U151); 
assign P3_ADD_546_U118 = ~P3_ADD_546_U16; 
assign P3_ADD_546_U126 = ~P3_ADD_546_U96; 
assign P3_ADD_546_U146 = ~(P3_ADD_546_U16 & P3_EAX_REG_7__SCAN_IN); 
assign P3_ADD_546_U147 = ~(P3_ADD_546_U96 & P3_EAX_REG_6__SCAN_IN); 
assign P3_ADD_476_U67 = ~(P3_ADD_476_U134 & P3_ADD_476_U133); 
assign P3_ADD_476_U96 = ~P3_ADD_476_U10; 
assign P3_ADD_476_U131 = ~(P3_ADD_476_U10 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_531_U71 = ~(P3_ADD_531_U141 & P3_ADD_531_U140); 
assign P3_ADD_531_U100 = ~P3_ADD_531_U11; 
assign P3_ADD_531_U138 = ~(P3_ADD_531_U11 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_SUB_320_U91 = ~(P3_SUB_320_U83 & P3_SUB_320_U58); 
assign P3_SUB_320_U135 = ~(P3_SUB_320_U83 & P3_SUB_320_U58); 
assign P3_ADD_505_U15 = ~(P3_ADD_505_U24 & P3_ADD_505_U23); 
assign P3_ADD_505_U20 = ~P3_ADD_505_U12; 
assign P3_ADD_505_U21 = ~(P3_ADD_505_U12 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_ADD_318_U67 = ~(P3_ADD_318_U134 & P3_ADD_318_U133); 
assign P3_ADD_318_U96 = ~P3_ADD_318_U10; 
assign P3_ADD_318_U131 = ~(P3_ADD_318_U10 & P3_PHYADDRPOINTER_REG_5__SCAN_IN); 
assign P3_SUB_370_U22 = ~(P3_SUB_370_U66 & P3_SUB_370_U65); 
assign P3_SUB_370_U28 = ~(P3_SUB_370_U33 & P3_SUB_370_U32); 
assign P3_ADD_315_U64 = ~(P3_ADD_315_U128 & P3_ADD_315_U127); 
assign P3_ADD_315_U93 = ~P3_ADD_315_U10; 
assign P3_ADD_315_U125 = ~(P3_ADD_315_U10 & P3_PHYADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_467_U67 = ~(P3_ADD_467_U134 & P3_ADD_467_U133); 
assign P3_ADD_467_U96 = ~P3_ADD_467_U10; 
assign P3_ADD_467_U131 = ~(P3_ADD_467_U10 & P3_REIP_REG_5__SCAN_IN); 
assign P3_ADD_430_U67 = ~(P3_ADD_430_U134 & P3_ADD_430_U133); 
assign P3_ADD_430_U96 = ~P3_ADD_430_U10; 
assign P3_ADD_430_U131 = ~(P3_ADD_430_U10 & P3_REIP_REG_5__SCAN_IN); 
assign P3_ADD_380_U71 = ~(P3_ADD_380_U141 & P3_ADD_380_U140); 
assign P3_ADD_380_U100 = ~P3_ADD_380_U11; 
assign P3_ADD_380_U138 = ~(P3_ADD_380_U11 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_344_U71 = ~(P3_ADD_344_U141 & P3_ADD_344_U140); 
assign P3_ADD_344_U100 = ~P3_ADD_344_U11; 
assign P3_ADD_344_U138 = ~(P3_ADD_344_U11 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_339_U67 = ~(P3_ADD_339_U134 & P3_ADD_339_U133); 
assign P3_ADD_339_U96 = ~P3_ADD_339_U10; 
assign P3_ADD_339_U131 = ~(P3_ADD_339_U10 & P3_PHYADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_541_U67 = ~(P3_ADD_541_U134 & P3_ADD_541_U133); 
assign P3_ADD_541_U96 = ~P3_ADD_541_U10; 
assign P3_ADD_541_U131 = ~(P3_ADD_541_U10 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_SUB_355_U22 = ~(P3_SUB_355_U66 & P3_SUB_355_U65); 
assign P3_SUB_355_U28 = ~(P3_SUB_355_U33 & P3_SUB_355_U32); 
assign P3_SUB_450_U19 = ~(P3_SUB_450_U63 & P3_SUB_450_U62); 
assign P3_SUB_450_U25 = ~(P3_SUB_450_U31 & P3_SUB_450_U30); 
assign P3_ADD_486_U15 = ~(P3_ADD_486_U24 & P3_ADD_486_U23); 
assign P3_ADD_486_U20 = ~P3_ADD_486_U12; 
assign P3_ADD_486_U21 = ~(P3_ADD_486_U12 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_SUB_485_U19 = ~(P3_SUB_485_U63 & P3_SUB_485_U62); 
assign P3_SUB_485_U25 = ~(P3_SUB_485_U31 & P3_SUB_485_U30); 
assign P3_ADD_515_U67 = ~(P3_ADD_515_U134 & P3_ADD_515_U133); 
assign P3_ADD_515_U96 = ~P3_ADD_515_U10; 
assign P3_ADD_515_U131 = ~(P3_ADD_515_U10 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_394_U68 = ~(P3_ADD_394_U138 & P3_ADD_394_U137); 
assign P3_ADD_394_U99 = ~P3_ADD_394_U10; 
assign P3_ADD_394_U135 = ~(P3_ADD_394_U10 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_SUB_414_U57 = P3_SUB_414_U133 & P3_SUB_414_U132; 
assign P3_SUB_414_U85 = ~P3_SUB_414_U23; 
assign P3_SUB_414_U90 = ~(P3_SUB_414_U89 & P3_EBX_REG_6__SCAN_IN); 
assign P3_SUB_414_U130 = ~(P3_SUB_414_U23 & P3_EBX_REG_7__SCAN_IN); 
assign P3_ADD_441_U67 = ~(P3_ADD_441_U134 & P3_ADD_441_U133); 
assign P3_ADD_441_U96 = ~P3_ADD_441_U10; 
assign P3_ADD_441_U131 = ~(P3_ADD_441_U10 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_349_U71 = ~(P3_ADD_349_U141 & P3_ADD_349_U140); 
assign P3_ADD_349_U100 = ~P3_ADD_349_U11; 
assign P3_ADD_349_U138 = ~(P3_ADD_349_U11 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_405_U68 = ~(P3_ADD_405_U138 & P3_ADD_405_U137); 
assign P3_ADD_405_U99 = ~P3_ADD_405_U10; 
assign P3_ADD_405_U135 = ~(P3_ADD_405_U10 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_553_U71 = ~(P3_ADD_553_U141 & P3_ADD_553_U140); 
assign P3_ADD_553_U100 = ~P3_ADD_553_U11; 
assign P3_ADD_553_U138 = ~(P3_ADD_553_U11 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_558_U71 = ~(P3_ADD_558_U141 & P3_ADD_558_U140); 
assign P3_ADD_558_U100 = ~P3_ADD_558_U11; 
assign P3_ADD_558_U138 = ~(P3_ADD_558_U11 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_385_U71 = ~(P3_ADD_385_U141 & P3_ADD_385_U140); 
assign P3_ADD_385_U100 = ~P3_ADD_385_U11; 
assign P3_ADD_385_U138 = ~(P3_ADD_385_U11 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_547_U71 = ~(P3_ADD_547_U141 & P3_ADD_547_U140); 
assign P3_ADD_547_U100 = ~P3_ADD_547_U11; 
assign P3_ADD_547_U138 = ~(P3_ADD_547_U11 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_SUB_412_U19 = ~(P3_SUB_412_U63 & P3_SUB_412_U62); 
assign P3_SUB_412_U25 = ~(P3_SUB_412_U31 & P3_SUB_412_U30); 
assign P3_SUB_504_U19 = ~(P3_SUB_504_U63 & P3_SUB_504_U62); 
assign P3_SUB_504_U25 = ~(P3_SUB_504_U31 & P3_SUB_504_U30); 
assign P3_SUB_401_U22 = ~(P3_SUB_401_U66 & P3_SUB_401_U65); 
assign P3_SUB_401_U28 = ~(P3_SUB_401_U33 & P3_SUB_401_U32); 
assign P3_SUB_390_U22 = ~(P3_SUB_390_U66 & P3_SUB_390_U65); 
assign P3_SUB_390_U28 = ~(P3_SUB_390_U33 & P3_SUB_390_U32); 
assign P3_ADD_495_U8 = ~(P3_ADD_495_U16 & P3_ADD_495_U15); 
assign P3_ADD_494_U67 = ~(P3_ADD_494_U134 & P3_ADD_494_U133); 
assign P3_ADD_494_U96 = ~P3_ADD_494_U10; 
assign P3_ADD_494_U131 = ~(P3_ADD_494_U10 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_536_U67 = ~(P3_ADD_536_U134 & P3_ADD_536_U133); 
assign P3_ADD_536_U96 = ~P3_ADD_536_U10; 
assign P3_ADD_536_U131 = ~(P3_ADD_536_U10 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P2_R2027_U71 = ~(P2_R2027_U141 & P2_R2027_U140); 
assign P2_R2027_U100 = ~P2_R2027_U11; 
assign P2_R2027_U138 = ~(P2_R2027_U11 & P2_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P2_R2337_U65 = ~(P2_R2337_U132 & P2_R2337_U131); 
assign P2_R2337_U97 = ~P2_R2337_U11; 
assign P2_R2337_U129 = ~(P2_R2337_U11 & P2_PHYADDRPOINTER_REG_6__SCAN_IN); 
assign P2_R2238_U22 = ~(P2_R2238_U66 & P2_R2238_U65); 
assign P2_R2238_U28 = ~(P2_R2238_U33 & P2_R2238_U32); 
assign P2_R1957_U21 = P2_U3682 | P2_U3683 | P2_U3671; 
assign P2_R1957_U49 = ~(P2_R1957_U149 & P2_R1957_U148); 
assign P2_R1957_U105 = ~(P2_U3671 & P2_R1957_U104); 
assign P2_SUB_450_U20 = ~(P2_SUB_450_U63 & P2_SUB_450_U62); 
assign P2_SUB_450_U26 = ~(P2_SUB_450_U31 & P2_SUB_450_U30); 
assign P2_ADD_394_U76 = ~(P2_ADD_394_U154 & P2_ADD_394_U153); 
assign P2_ADD_394_U99 = ~P2_ADD_394_U10; 
assign P2_ADD_394_U159 = ~(P2_ADD_394_U10 & P2_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P2_ADD_371_1212_U8 = P2_ADD_371_1212_U9 & P2_ADD_371_1212_U91; 
assign P2_ADD_371_1212_U103 = P2_ADD_371_1212_U9 & P2_ADD_371_1212_U104; 
assign P2_ADD_371_1212_U109 = P2_ADD_371_1212_U9 & P2_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P1_R2027_U55 = ~(P1_R2027_U150 & P1_R2027_U149); 
assign P1_R2027_U56 = ~(P1_R2027_U152 & P1_R2027_U151); 
assign P1_R2027_U118 = ~P1_R2027_U16; 
assign P1_R2027_U126 = ~P1_R2027_U96; 
assign P1_R2027_U146 = ~(P1_R2027_U16 & P1_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P1_R2027_U147 = ~(P1_R2027_U96 & P1_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P1_R2337_U67 = ~(P1_R2337_U134 & P1_R2337_U133); 
assign P1_R2337_U96 = ~P1_R2337_U10; 
assign P1_R2337_U131 = ~(P1_R2337_U10 & P1_PHYADDRPOINTER_REG_5__SCAN_IN); 
assign P1_R2096_U67 = ~(P1_R2096_U134 & P1_R2096_U133); 
assign P1_R2096_U96 = ~P1_R2096_U10; 
assign P1_R2096_U131 = ~(P1_R2096_U10 & P1_REIP_REG_5__SCAN_IN); 
assign P1_R2238_U22 = ~(P1_R2238_U66 & P1_R2238_U65); 
assign P1_R2238_U28 = ~(P1_R2238_U33 & P1_R2238_U32); 
assign P1_SUB_450_U22 = ~(P1_SUB_450_U66 & P1_SUB_450_U65); 
assign P1_SUB_450_U28 = ~(P1_SUB_450_U33 & P1_SUB_450_U32); 
assign P1_ADD_405_U76 = ~(P1_ADD_405_U154 & P1_ADD_405_U153); 
assign P1_ADD_405_U99 = ~P1_ADD_405_U10; 
assign P1_ADD_405_U159 = ~(P1_ADD_405_U10 & P1_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P1_ADD_515_U76 = ~(P1_ADD_515_U152 & P1_ADD_515_U151); 
assign P1_ADD_515_U96 = ~P1_ADD_515_U10; 
assign P1_ADD_515_U157 = ~(P1_ADD_515_U10 & P1_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign U207 = U250 & U214; 
assign U283 = ~(U550 & U549); 
assign U284 = ~(U552 & U551); 
assign U285 = ~(U554 & U553); 
assign U286 = ~(U556 & U555); 
assign U287 = ~(U558 & U557); 
assign U288 = ~(U560 & U559); 
assign U289 = ~(U562 & U561); 
assign U290 = ~(U564 & U563); 
assign U291 = ~(U566 & U565); 
assign U292 = ~(U568 & U567); 
assign U293 = ~(U570 & U569); 
assign U294 = ~(U572 & U571); 
assign U295 = ~(U574 & U573); 
assign U296 = ~(U576 & U575); 
assign U297 = ~(U578 & U577); 
assign U298 = ~(U580 & U579); 
assign U299 = ~(U582 & U581); 
assign U300 = ~(U584 & U583); 
assign U301 = ~(U586 & U585); 
assign U302 = ~(U588 & U587); 
assign U303 = ~(U590 & U589); 
assign U304 = ~(U592 & U591); 
assign U305 = ~(U594 & U593); 
assign U306 = ~(U596 & U595); 
assign U307 = ~(U598 & U597); 
assign U308 = ~(U600 & U599); 
assign U309 = ~(U602 & U601); 
assign U310 = ~(U604 & U603); 
assign U311 = ~(U606 & U605); 
assign U312 = ~(U608 & U607); 
assign U313 = ~(U610 & U609); 
assign U314 = ~(U612 & U611); 
assign U315 = ~(U614 & U613); 
assign U316 = ~(U616 & U615); 
assign U317 = ~(U618 & U617); 
assign U318 = ~(U620 & U619); 
assign U319 = ~(U622 & U621); 
assign U320 = ~(U624 & U623); 
assign U321 = ~(U626 & U625); 
assign U322 = ~(U628 & U627); 
assign U323 = ~(U630 & U629); 
assign U324 = ~(U632 & U631); 
assign U325 = ~(U634 & U633); 
assign U326 = ~(U636 & U635); 
assign U327 = ~(U638 & U637); 
assign U328 = ~(U640 & U639); 
assign U329 = ~(U642 & U641); 
assign U330 = ~(U644 & U643); 
assign U331 = ~(U646 & U645); 
assign U332 = ~(U648 & U647); 
assign U333 = ~(U650 & U649); 
assign U334 = ~(U652 & U651); 
assign U335 = ~(U654 & U653); 
assign U336 = ~(U656 & U655); 
assign U337 = ~(U658 & U657); 
assign U338 = ~(U660 & U659); 
assign U339 = ~(U662 & U661); 
assign U340 = ~(U664 & U663); 
assign U341 = ~(U666 & U665); 
assign U342 = ~(U668 & U667); 
assign U343 = ~(U670 & U669); 
assign U344 = ~(U672 & U671); 
assign U345 = ~(U674 & U673); 
assign U346 = ~(U676 & U675); 
assign U388 = ~U250; 
assign U390 = ~(U385 & P1_DATAO_REG_0__SCAN_IN); 
assign U393 = ~(U385 & P1_DATAO_REG_1__SCAN_IN); 
assign U396 = ~(U385 & P1_DATAO_REG_2__SCAN_IN); 
assign U399 = ~(U385 & P1_DATAO_REG_3__SCAN_IN); 
assign U402 = ~(U385 & P1_DATAO_REG_4__SCAN_IN); 
assign U405 = ~(U385 & P1_DATAO_REG_5__SCAN_IN); 
assign U408 = ~(U385 & P1_DATAO_REG_6__SCAN_IN); 
assign U411 = ~(U385 & P1_DATAO_REG_7__SCAN_IN); 
assign U414 = ~(U385 & P1_DATAO_REG_8__SCAN_IN); 
assign U417 = ~(U385 & P1_DATAO_REG_9__SCAN_IN); 
assign U420 = ~(U385 & P1_DATAO_REG_10__SCAN_IN); 
assign U423 = ~(U385 & P1_DATAO_REG_11__SCAN_IN); 
assign U426 = ~(U385 & P1_DATAO_REG_12__SCAN_IN); 
assign U429 = ~(U385 & P1_DATAO_REG_13__SCAN_IN); 
assign U432 = ~(U385 & P1_DATAO_REG_14__SCAN_IN); 
assign U435 = ~(U385 & P1_DATAO_REG_15__SCAN_IN); 
assign U438 = ~(U385 & P1_DATAO_REG_16__SCAN_IN); 
assign U441 = ~(U385 & P1_DATAO_REG_17__SCAN_IN); 
assign U444 = ~(U385 & P1_DATAO_REG_18__SCAN_IN); 
assign U447 = ~(U385 & P1_DATAO_REG_19__SCAN_IN); 
assign U450 = ~(U385 & P1_DATAO_REG_20__SCAN_IN); 
assign U453 = ~(U385 & P1_DATAO_REG_21__SCAN_IN); 
assign U456 = ~(U385 & P1_DATAO_REG_22__SCAN_IN); 
assign U459 = ~(U385 & P1_DATAO_REG_23__SCAN_IN); 
assign U462 = ~(U385 & P1_DATAO_REG_24__SCAN_IN); 
assign U465 = ~(U385 & P1_DATAO_REG_25__SCAN_IN); 
assign U468 = ~(U385 & P1_DATAO_REG_26__SCAN_IN); 
assign U471 = ~(U385 & P1_DATAO_REG_27__SCAN_IN); 
assign U474 = ~(U385 & P1_DATAO_REG_28__SCAN_IN); 
assign U477 = ~(U385 & P1_DATAO_REG_29__SCAN_IN); 
assign U480 = ~(U385 & P1_DATAO_REG_30__SCAN_IN); 
assign U483 = ~(U385 & P1_DATAO_REG_31__SCAN_IN); 
assign P3_U2421 = P3_U2379 & BUF2_REG_24__SCAN_IN; 
assign P3_U2422 = P3_U2379 & BUF2_REG_16__SCAN_IN; 
assign P3_U2423 = P3_U2379 & BUF2_REG_25__SCAN_IN; 
assign P3_U2424 = P3_U2379 & BUF2_REG_17__SCAN_IN; 
assign P3_U2425 = P3_U2379 & BUF2_REG_26__SCAN_IN; 
assign P3_U2426 = P3_U2379 & BUF2_REG_18__SCAN_IN; 
assign P3_U2427 = P3_U2379 & BUF2_REG_27__SCAN_IN; 
assign P3_U2428 = P3_U2379 & BUF2_REG_19__SCAN_IN; 
assign P3_U2429 = P3_U2379 & BUF2_REG_28__SCAN_IN; 
assign P3_U2430 = P3_U2379 & BUF2_REG_20__SCAN_IN; 
assign P3_U2431 = P3_U2379 & BUF2_REG_29__SCAN_IN; 
assign P3_U2432 = P3_U2379 & BUF2_REG_21__SCAN_IN; 
assign P3_U2433 = P3_U2379 & BUF2_REG_30__SCAN_IN; 
assign P3_U2434 = P3_U2379 & BUF2_REG_22__SCAN_IN; 
assign P3_U2435 = P3_U2379 & BUF2_REG_31__SCAN_IN; 
assign P3_U2436 = P3_U2379 & BUF2_REG_23__SCAN_IN; 
assign P3_U2457 = P3_U3269 & P3_U3139; 
assign P3_U2459 = P3_U7962 & P3_U3139; 
assign P3_U2520 = P3_U5543 & P3_U5548; 
assign P3_U2528 = P3_U5543 & P3_U3225; 
assign P3_U2534 = P3_U2533 & P3_U2519; 
assign P3_U2535 = P3_U2533 & P3_U2522; 
assign P3_U2536 = P3_U2533 & P3_U2524; 
assign P3_U2537 = P3_U2533 & P3_U2526; 
assign P3_U2539 = P3_U2519 & P3_U2538; 
assign P3_U2540 = P3_U2522 & P3_U2538; 
assign P3_U2541 = P3_U2524 & P3_U2538; 
assign P3_U2542 = P3_U2526 & P3_U2538; 
assign P3_U2544 = P3_U2543 & P3_U2468; 
assign P3_U2545 = P3_U2543 & P3_U4467; 
assign P3_U2546 = P3_U2543 & P3_U4332; 
assign P3_U2547 = P3_U2543 & P3_U2466; 
assign P3_U2549 = P3_U2548 & P3_U2468; 
assign P3_U2550 = P3_U2548 & P3_U4467; 
assign P3_U2551 = P3_U2548 & P3_U4332; 
assign P3_U2552 = P3_U2548 & P3_U2466; 
assign P3_U2553 = P3_U7516 & P3_U3272; 
assign P3_U2558 = P3_U7516 & P3_U8034; 
assign P3_U2563 = P3_U8037 & P3_U4291; 
assign P3_U2568 = P3_U8037 & P3_U3267; 
assign P3_U2574 = P3_U2573 & P3_U2522; 
assign P3_U2575 = P3_U2573 & P3_U2519; 
assign P3_U2576 = P3_U2573 & P3_U2526; 
assign P3_U2577 = P3_U2573 & P3_U2524; 
assign P3_U2579 = P3_U2578 & P3_U2522; 
assign P3_U2580 = P3_U2578 & P3_U2519; 
assign P3_U2581 = P3_U2578 & P3_U2526; 
assign P3_U2582 = P3_U2578 & P3_U2524; 
assign P3_U2633 = ~(P3_U7937 & P3_U7383); 
assign P3_U2999 = P3_U7937 & P3_DATAWIDTH_REG_31__SCAN_IN; 
assign P3_U3000 = P3_U7937 & P3_DATAWIDTH_REG_30__SCAN_IN; 
assign P3_U3001 = P3_U7937 & P3_DATAWIDTH_REG_29__SCAN_IN; 
assign P3_U3002 = P3_U7937 & P3_DATAWIDTH_REG_28__SCAN_IN; 
assign P3_U3003 = P3_U7937 & P3_DATAWIDTH_REG_27__SCAN_IN; 
assign P3_U3004 = P3_U7937 & P3_DATAWIDTH_REG_26__SCAN_IN; 
assign P3_U3005 = P3_U7937 & P3_DATAWIDTH_REG_25__SCAN_IN; 
assign P3_U3006 = P3_U7937 & P3_DATAWIDTH_REG_24__SCAN_IN; 
assign P3_U3007 = P3_U7937 & P3_DATAWIDTH_REG_23__SCAN_IN; 
assign P3_U3008 = P3_U7937 & P3_DATAWIDTH_REG_22__SCAN_IN; 
assign P3_U3009 = P3_U7937 & P3_DATAWIDTH_REG_21__SCAN_IN; 
assign P3_U3010 = P3_U7937 & P3_DATAWIDTH_REG_20__SCAN_IN; 
assign P3_U3011 = P3_U7937 & P3_DATAWIDTH_REG_19__SCAN_IN; 
assign P3_U3012 = P3_U7937 & P3_DATAWIDTH_REG_18__SCAN_IN; 
assign P3_U3013 = P3_U7937 & P3_DATAWIDTH_REG_17__SCAN_IN; 
assign P3_U3014 = P3_U7937 & P3_DATAWIDTH_REG_16__SCAN_IN; 
assign P3_U3015 = P3_U7937 & P3_DATAWIDTH_REG_15__SCAN_IN; 
assign P3_U3016 = P3_U7937 & P3_DATAWIDTH_REG_14__SCAN_IN; 
assign P3_U3017 = P3_U7937 & P3_DATAWIDTH_REG_13__SCAN_IN; 
assign P3_U3018 = P3_U7937 & P3_DATAWIDTH_REG_12__SCAN_IN; 
assign P3_U3019 = P3_U7937 & P3_DATAWIDTH_REG_11__SCAN_IN; 
assign P3_U3020 = P3_U7937 & P3_DATAWIDTH_REG_10__SCAN_IN; 
assign P3_U3021 = P3_U7937 & P3_DATAWIDTH_REG_9__SCAN_IN; 
assign P3_U3022 = P3_U7937 & P3_DATAWIDTH_REG_8__SCAN_IN; 
assign P3_U3023 = P3_U7937 & P3_DATAWIDTH_REG_7__SCAN_IN; 
assign P3_U3024 = P3_U7937 & P3_DATAWIDTH_REG_6__SCAN_IN; 
assign P3_U3025 = P3_U7937 & P3_DATAWIDTH_REG_5__SCAN_IN; 
assign P3_U3026 = P3_U7937 & P3_DATAWIDTH_REG_4__SCAN_IN; 
assign P3_U3027 = P3_U7937 & P3_DATAWIDTH_REG_3__SCAN_IN; 
assign P3_U3028 = P3_U7937 & P3_DATAWIDTH_REG_2__SCAN_IN; 
assign P3_U3030 = ~(P3_U7932 & P3_U7931 & P3_U3311); 
assign P3_U3032 = ~(P3_U4443 & P3_U4442 & P3_U4444); 
assign P3_U3033 = ~(P3_U4440 & P3_U4439 & P3_U4441); 
assign P3_U3034 = ~(P3_U4437 & P3_U4436 & P3_U4438); 
assign P3_U3035 = ~(P3_U4434 & P3_U4433 & P3_U4435); 
assign P3_U3036 = ~(P3_U4431 & P3_U4430 & P3_U4432); 
assign P3_U3037 = ~(P3_U4428 & P3_U4427 & P3_U4429); 
assign P3_U3038 = ~(P3_U4425 & P3_U4424 & P3_U4426); 
assign P3_U3039 = ~(P3_U4422 & P3_U4421 & P3_U4423); 
assign P3_U3040 = ~(P3_U4419 & P3_U4418 & P3_U4420); 
assign P3_U3041 = ~(P3_U4416 & P3_U4415 & P3_U4417); 
assign P3_U3042 = ~(P3_U4413 & P3_U4412 & P3_U4414); 
assign P3_U3043 = ~(P3_U4410 & P3_U4409 & P3_U4411); 
assign P3_U3044 = ~(P3_U4407 & P3_U4406 & P3_U4408); 
assign P3_U3045 = ~(P3_U4404 & P3_U4403 & P3_U4405); 
assign P3_U3046 = ~(P3_U4401 & P3_U4400 & P3_U4402); 
assign P3_U3047 = ~(P3_U4398 & P3_U4397 & P3_U4399); 
assign P3_U3048 = ~(P3_U4395 & P3_U4394 & P3_U4396); 
assign P3_U3049 = ~(P3_U4392 & P3_U4391 & P3_U4393); 
assign P3_U3050 = ~(P3_U4389 & P3_U4388 & P3_U4390); 
assign P3_U3051 = ~(P3_U4386 & P3_U4385 & P3_U4387); 
assign P3_U3052 = ~(P3_U4383 & P3_U4382 & P3_U4384); 
assign P3_U3053 = ~(P3_U4380 & P3_U4379 & P3_U4381); 
assign P3_U3054 = ~(P3_U4377 & P3_U4376 & P3_U4378); 
assign P3_U3055 = ~(P3_U4374 & P3_U4373 & P3_U4375); 
assign P3_U3056 = ~(P3_U4371 & P3_U4370 & P3_U4372); 
assign P3_U3057 = ~(P3_U4368 & P3_U4367 & P3_U4369); 
assign P3_U3058 = ~(P3_U4365 & P3_U4364 & P3_U4366); 
assign P3_U3059 = ~(P3_U4362 & P3_U4361 & P3_U4363); 
assign P3_U3060 = ~(P3_U4359 & P3_U4358 & P3_U4360); 
assign P3_U3061 = ~(P3_U4356 & P3_U4355 & P3_U4357); 
assign P3_U3140 = ~(P3_U3141 & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P3_U3148 = ~(P3_U3141 & P3_U3128); 
assign P3_U3270 = ~(P3_U7964 & P3_U7963); 
assign P3_U3292 = ~(P3_U8011 & P3_U8010); 
assign P3_U3300 = ~(P3_U8039 & P3_U8038); 
assign P3_U3310 = P3_U4456 & P3_U3080; 
assign P3_U3313 = P3_U4475 & P3_U4474 & P3_U4473 & P3_U4472; 
assign P3_U3314 = P3_U4479 & P3_U4478 & P3_U4477 & P3_U4476; 
assign P3_U3315 = P3_U4481 & P3_U4480; 
assign P3_U3316 = P3_U4483 & P3_U4482; 
assign P3_U3318 = P3_U4492 & P3_U4491 & P3_U4490 & P3_U4489; 
assign P3_U3319 = P3_U4496 & P3_U4495 & P3_U4494 & P3_U4493; 
assign P3_U3320 = P3_U4498 & P3_U4497; 
assign P3_U3321 = P3_U4500 & P3_U4499; 
assign P3_U3323 = P3_U4509 & P3_U4508 & P3_U4507 & P3_U4506; 
assign P3_U3324 = P3_U4513 & P3_U4512 & P3_U4511 & P3_U4510; 
assign P3_U3325 = P3_U4515 & P3_U4514; 
assign P3_U3326 = P3_U4517 & P3_U4516; 
assign P3_U3328 = P3_U4543 & P3_U4542 & P3_U4541 & P3_U4540; 
assign P3_U3329 = P3_U4547 & P3_U4546 & P3_U4545 & P3_U4544; 
assign P3_U3330 = P3_U4549 & P3_U4548; 
assign P3_U3331 = P3_U4551 & P3_U4550; 
assign P3_U3333 = P3_U4560 & P3_U4559 & P3_U4558 & P3_U4557; 
assign P3_U3334 = P3_U4564 & P3_U4563 & P3_U4562 & P3_U4561; 
assign P3_U3335 = P3_U4566 & P3_U4565; 
assign P3_U3336 = P3_U4568 & P3_U4567; 
assign P3_U3338 = P3_U4526 & P3_U4525 & P3_U4524 & P3_U4523; 
assign P3_U3339 = P3_U4530 & P3_U4529 & P3_U4528 & P3_U4527; 
assign P3_U3340 = P3_U4532 & P3_U4531; 
assign P3_U3341 = P3_U4534 & P3_U4533; 
assign P3_U3343 = P3_U4594 & P3_U4593 & P3_U4592 & P3_U4591; 
assign P3_U3344 = P3_U4598 & P3_U4597 & P3_U4596 & P3_U4595; 
assign P3_U3345 = P3_U4600 & P3_U4599; 
assign P3_U3346 = P3_U4602 & P3_U4601; 
assign P3_U3348 = P3_U4577 & P3_U4576 & P3_U4575 & P3_U4574; 
assign P3_U3349 = P3_U4581 & P3_U4580 & P3_U4579 & P3_U4578; 
assign P3_U3350 = P3_U4583 & P3_U4582; 
assign P3_U3351 = P3_U4585 & P3_U4584; 
assign P3_U3369 = P3_U4671 & P3_U4312; 
assign P3_U3510 = P3_U5082 & P3_U4312; 
assign P3_U3652 = P3_U4340 & P3_ADD_495_U8; 
assign P3_U3680 = P3_U5555 & P3_U5554; 
assign P3_U4248 = P3_U7779 & P3_U7778 & P3_U7777 & P3_U7776; 
assign P3_U4249 = P3_U7783 & P3_U7782 & P3_U7781 & P3_U7780; 
assign P3_U4251 = P3_U7791 & P3_U7790 & P3_U7789 & P3_U7788; 
assign P3_U4252 = P3_U7795 & P3_U7794 & P3_U7793 & P3_U7792; 
assign P3_U4253 = P3_U7799 & P3_U7798 & P3_U7797 & P3_U7796; 
assign P3_U4255 = P3_U7807 & P3_U7806 & P3_U7805 & P3_U7804; 
assign P3_U4256 = P3_U7811 & P3_U7810 & P3_U7809 & P3_U7808; 
assign P3_U4257 = P3_U7815 & P3_U7814 & P3_U7813 & P3_U7812; 
assign P3_U4259 = P3_U7823 & P3_U7822 & P3_U7821 & P3_U7820; 
assign P3_U4260 = P3_U7827 & P3_U7826 & P3_U7825 & P3_U7824; 
assign P3_U4261 = P3_U7831 & P3_U7830 & P3_U7829 & P3_U7828; 
assign P3_U4263 = P3_U7839 & P3_U7838 & P3_U7837 & P3_U7836; 
assign P3_U4264 = P3_U7843 & P3_U7842 & P3_U7841 & P3_U7840; 
assign P3_U4265 = P3_U7847 & P3_U7846 & P3_U7845 & P3_U7844; 
assign P3_U4267 = P3_U7855 & P3_U7854 & P3_U7853 & P3_U7852; 
assign P3_U4268 = P3_U7859 & P3_U7858 & P3_U7857 & P3_U7856; 
assign P3_U4269 = P3_U7863 & P3_U7862 & P3_U7861 & P3_U7860; 
assign P3_U4271 = P3_U7871 & P3_U7870 & P3_U7869 & P3_U7868; 
assign P3_U4272 = P3_U7875 & P3_U7874 & P3_U7873 & P3_U7872; 
assign P3_U4273 = P3_U7879 & P3_U7878 & P3_U7877 & P3_U7876; 
assign P3_U4275 = P3_U7887 & P3_U7886 & P3_U7885 & P3_U7884; 
assign P3_U4276 = P3_U7891 & P3_U7890 & P3_U7889 & P3_U7888; 
assign P3_U4277 = P3_U7895 & P3_U7894 & P3_U7893 & P3_U7892; 
assign P3_U4279 = P3_U7903 & P3_U7902 & P3_U7901 & P3_U7900; 
assign P3_U4294 = ~P3_U3106; 
assign P3_U4457 = ~(P3_U4451 & P3_STATE_REG_2__SCAN_IN); 
assign P3_U4643 = ~P3_U3141; 
assign P3_U4652 = ~P3_U3139; 
assign P3_U4655 = ~(P3_U4654 & P3_U3139); 
assign P3_U5567 = ~(P3_U3286 & P3_U7985 & P3_STATE2_REG_1__SCAN_IN); 
assign P3_U5588 = ~(P3_U4650 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U5605 = ~(P3_U5582 & P3_U3141); 
assign P3_U7784 = ~(P3_U2591 & P3_INSTQUEUE_REG_0__7__SCAN_IN); 
assign P3_U7785 = ~(P3_U2590 & P3_INSTQUEUE_REG_1__7__SCAN_IN); 
assign P3_U7786 = ~(P3_U2589 & P3_INSTQUEUE_REG_2__7__SCAN_IN); 
assign P3_U7787 = ~(P3_U2588 & P3_INSTQUEUE_REG_3__7__SCAN_IN); 
assign P3_U7800 = ~(P3_U2591 & P3_INSTQUEUE_REG_0__6__SCAN_IN); 
assign P3_U7801 = ~(P3_U2590 & P3_INSTQUEUE_REG_1__6__SCAN_IN); 
assign P3_U7802 = ~(P3_U2589 & P3_INSTQUEUE_REG_2__6__SCAN_IN); 
assign P3_U7803 = ~(P3_U2588 & P3_INSTQUEUE_REG_3__6__SCAN_IN); 
assign P3_U7816 = ~(P3_U2591 & P3_INSTQUEUE_REG_0__5__SCAN_IN); 
assign P3_U7817 = ~(P3_U2590 & P3_INSTQUEUE_REG_1__5__SCAN_IN); 
assign P3_U7818 = ~(P3_U2589 & P3_INSTQUEUE_REG_2__5__SCAN_IN); 
assign P3_U7819 = ~(P3_U2588 & P3_INSTQUEUE_REG_3__5__SCAN_IN); 
assign P3_U7832 = ~(P3_U2591 & P3_INSTQUEUE_REG_0__4__SCAN_IN); 
assign P3_U7833 = ~(P3_U2590 & P3_INSTQUEUE_REG_1__4__SCAN_IN); 
assign P3_U7834 = ~(P3_U2589 & P3_INSTQUEUE_REG_2__4__SCAN_IN); 
assign P3_U7835 = ~(P3_U2588 & P3_INSTQUEUE_REG_3__4__SCAN_IN); 
assign P3_U7848 = ~(P3_U2591 & P3_INSTQUEUE_REG_0__3__SCAN_IN); 
assign P3_U7849 = ~(P3_U2590 & P3_INSTQUEUE_REG_1__3__SCAN_IN); 
assign P3_U7850 = ~(P3_U2589 & P3_INSTQUEUE_REG_2__3__SCAN_IN); 
assign P3_U7851 = ~(P3_U2588 & P3_INSTQUEUE_REG_3__3__SCAN_IN); 
assign P3_U7864 = ~(P3_U2591 & P3_INSTQUEUE_REG_0__2__SCAN_IN); 
assign P3_U7865 = ~(P3_U2590 & P3_INSTQUEUE_REG_1__2__SCAN_IN); 
assign P3_U7866 = ~(P3_U2589 & P3_INSTQUEUE_REG_2__2__SCAN_IN); 
assign P3_U7867 = ~(P3_U2588 & P3_INSTQUEUE_REG_3__2__SCAN_IN); 
assign P3_U7880 = ~(P3_U2591 & P3_INSTQUEUE_REG_0__1__SCAN_IN); 
assign P3_U7881 = ~(P3_U2590 & P3_INSTQUEUE_REG_1__1__SCAN_IN); 
assign P3_U7882 = ~(P3_U2589 & P3_INSTQUEUE_REG_2__1__SCAN_IN); 
assign P3_U7883 = ~(P3_U2588 & P3_INSTQUEUE_REG_3__1__SCAN_IN); 
assign P3_U7896 = ~(P3_U2591 & P3_INSTQUEUE_REG_0__0__SCAN_IN); 
assign P3_U7897 = ~(P3_U2590 & P3_INSTQUEUE_REG_1__0__SCAN_IN); 
assign P3_U7898 = ~(P3_U2589 & P3_INSTQUEUE_REG_2__0__SCAN_IN); 
assign P3_U7899 = ~(P3_U2588 & P3_INSTQUEUE_REG_3__0__SCAN_IN); 
assign P3_U7934 = ~(P3_U4459 & P3_U3079); 
assign P3_U7938 = ~(P3_U7937 & P3_DATAWIDTH_REG_0__SCAN_IN); 
assign P3_U7941 = ~(P3_U7937 & P3_DATAWIDTH_REG_1__SCAN_IN); 
assign P3_U8020 = ~(P3_U7937 & P3_STATEBS16_REG_SCAN_IN); 
assign P3_U8041 = ~(P3_U3286 & P3_U7985 & P3_FLUSH_REG_SCAN_IN); 
assign P2_U2356 = P2_U3253 & P2_STATE2_REG_0__SCAN_IN; 
assign P2_U2439 = P2_U4339 & P2_U3521; 
assign P2_U2447 = P2_U2616 & P2_STATE2_REG_0__SCAN_IN; 
assign P2_U2449 = P2_U3278 & P2_U3521; 
assign P2_U2457 = P2_U3521 & P2_U3255; 
assign P2_U2517 = P2_U2515 & P2_U2516; 
assign P2_U2519 = P2_U2515 & P2_U2518; 
assign P2_U2521 = P2_U2520 & P2_U2516; 
assign P2_U2522 = P2_U2520 & P2_U2518; 
assign P2_U2524 = P2_U2515 & P2_U2523; 
assign P2_U2526 = P2_U2515 & P2_U2525; 
assign P2_U2527 = P2_U2520 & P2_U2523; 
assign P2_U2528 = P2_U2520 & P2_U2525; 
assign P2_U2545 = P2_U2544 & P2_U2540; 
assign P2_U2546 = P2_U2544 & P2_U2542; 
assign P2_U2551 = P2_U2544 & P2_U2547; 
assign P2_U2552 = P2_U2544 & P2_U2549; 
assign P2_U2565 = P2_U2564 & P2_U2563; 
assign P2_U2567 = P2_U2564 & P2_U2566; 
assign P2_U2569 = P2_U2564 & P2_U2568; 
assign P2_U2571 = P2_U2564 & P2_U2570; 
assign P2_U2573 = P2_U2572 & P2_U2563; 
assign P2_U2574 = P2_U2572 & P2_U2566; 
assign P2_U2575 = P2_U2572 & P2_U2568; 
assign P2_U2576 = P2_U2572 & P2_U2570; 
assign P2_U2577 = P2_U4409 & P2_U8149; 
assign P2_U2582 = P2_U8149 & P2_U3553; 
assign P2_U2815 = ~(P2_U7917 & P2_U6856); 
assign P2_U3179 = P2_U7917 & P2_DATAWIDTH_REG_31__SCAN_IN; 
assign P2_U3180 = P2_U7917 & P2_DATAWIDTH_REG_30__SCAN_IN; 
assign P2_U3181 = P2_U7917 & P2_DATAWIDTH_REG_29__SCAN_IN; 
assign P2_U3182 = P2_U7917 & P2_DATAWIDTH_REG_28__SCAN_IN; 
assign P2_U3183 = P2_U7917 & P2_DATAWIDTH_REG_27__SCAN_IN; 
assign P2_U3184 = P2_U7917 & P2_DATAWIDTH_REG_26__SCAN_IN; 
assign P2_U3185 = P2_U7917 & P2_DATAWIDTH_REG_25__SCAN_IN; 
assign P2_U3186 = P2_U7917 & P2_DATAWIDTH_REG_24__SCAN_IN; 
assign P2_U3187 = P2_U7917 & P2_DATAWIDTH_REG_23__SCAN_IN; 
assign P2_U3188 = P2_U7917 & P2_DATAWIDTH_REG_22__SCAN_IN; 
assign P2_U3189 = P2_U7917 & P2_DATAWIDTH_REG_21__SCAN_IN; 
assign P2_U3190 = P2_U7917 & P2_DATAWIDTH_REG_20__SCAN_IN; 
assign P2_U3191 = P2_U7917 & P2_DATAWIDTH_REG_19__SCAN_IN; 
assign P2_U3192 = P2_U7917 & P2_DATAWIDTH_REG_18__SCAN_IN; 
assign P2_U3193 = P2_U7917 & P2_DATAWIDTH_REG_17__SCAN_IN; 
assign P2_U3194 = P2_U7917 & P2_DATAWIDTH_REG_16__SCAN_IN; 
assign P2_U3195 = P2_U7917 & P2_DATAWIDTH_REG_15__SCAN_IN; 
assign P2_U3196 = P2_U7917 & P2_DATAWIDTH_REG_14__SCAN_IN; 
assign P2_U3197 = P2_U7917 & P2_DATAWIDTH_REG_13__SCAN_IN; 
assign P2_U3198 = P2_U7917 & P2_DATAWIDTH_REG_12__SCAN_IN; 
assign P2_U3199 = P2_U7917 & P2_DATAWIDTH_REG_11__SCAN_IN; 
assign P2_U3200 = P2_U7917 & P2_DATAWIDTH_REG_10__SCAN_IN; 
assign P2_U3201 = P2_U7917 & P2_DATAWIDTH_REG_9__SCAN_IN; 
assign P2_U3202 = P2_U7917 & P2_DATAWIDTH_REG_8__SCAN_IN; 
assign P2_U3203 = P2_U7917 & P2_DATAWIDTH_REG_7__SCAN_IN; 
assign P2_U3204 = P2_U7917 & P2_DATAWIDTH_REG_6__SCAN_IN; 
assign P2_U3205 = P2_U7917 & P2_DATAWIDTH_REG_5__SCAN_IN; 
assign P2_U3206 = P2_U7917 & P2_DATAWIDTH_REG_4__SCAN_IN; 
assign P2_U3207 = P2_U7917 & P2_DATAWIDTH_REG_3__SCAN_IN; 
assign P2_U3208 = P2_U7917 & P2_DATAWIDTH_REG_2__SCAN_IN; 
assign P2_U3210 = ~(P2_U7912 & P2_U7911 & P2_U3691); 
assign P2_U3212 = ~(P2_U4566 & P2_U4565 & P2_U4567); 
assign P2_U3213 = ~(P2_U4563 & P2_U4562 & P2_U4564); 
assign P2_U3214 = ~(P2_U4560 & P2_U4559 & P2_U4561); 
assign P2_U3215 = ~(P2_U4557 & P2_U4556 & P2_U4558); 
assign P2_U3216 = ~(P2_U4554 & P2_U4553 & P2_U4555); 
assign P2_U3217 = ~(P2_U4551 & P2_U4550 & P2_U4552); 
assign P2_U3218 = ~(P2_U4548 & P2_U4547 & P2_U4549); 
assign P2_U3219 = ~(P2_U4545 & P2_U4544 & P2_U4546); 
assign P2_U3220 = ~(P2_U4542 & P2_U4541 & P2_U4543); 
assign P2_U3221 = ~(P2_U4539 & P2_U4538 & P2_U4540); 
assign P2_U3222 = ~(P2_U4536 & P2_U4535 & P2_U4537); 
assign P2_U3223 = ~(P2_U4533 & P2_U4532 & P2_U4534); 
assign P2_U3224 = ~(P2_U4530 & P2_U4529 & P2_U4531); 
assign P2_U3225 = ~(P2_U4527 & P2_U4526 & P2_U4528); 
assign P2_U3226 = ~(P2_U4524 & P2_U4523 & P2_U4525); 
assign P2_U3227 = ~(P2_U4521 & P2_U4520 & P2_U4522); 
assign P2_U3228 = ~(P2_U4518 & P2_U4517 & P2_U4519); 
assign P2_U3229 = ~(P2_U4515 & P2_U4514 & P2_U4516); 
assign P2_U3230 = ~(P2_U4512 & P2_U4511 & P2_U4513); 
assign P2_U3231 = ~(P2_U4509 & P2_U4508 & P2_U4510); 
assign P2_U3232 = ~(P2_U4506 & P2_U4505 & P2_U4507); 
assign P2_U3233 = ~(P2_U4503 & P2_U4502 & P2_U4504); 
assign P2_U3234 = ~(P2_U4500 & P2_U4499 & P2_U4501); 
assign P2_U3235 = ~(P2_U4497 & P2_U4496 & P2_U4498); 
assign P2_U3236 = ~(P2_U4494 & P2_U4493 & P2_U4495); 
assign P2_U3237 = ~(P2_U4491 & P2_U4490 & P2_U4492); 
assign P2_U3238 = ~(P2_U4488 & P2_U4487 & P2_U4489); 
assign P2_U3239 = ~(P2_U4485 & P2_U4484 & P2_U4486); 
assign P2_U3240 = ~(P2_U4482 & P2_U4481 & P2_U4483); 
assign P2_U3241 = ~(P2_U4479 & P2_U4478 & P2_U4480); 
assign P2_U3247 = ~(P2_U2442 & P2_U3243); 
assign P2_U3248 = ~(P2_U2442 & P2_U4650); 
assign P2_U3249 = ~(P2_U2441 & P2_U3243); 
assign P2_U3250 = ~(P2_U2441 & P2_U4650); 
assign P2_U3251 = ~(P2_U2443 & P2_U3243); 
assign P2_U3252 = ~(P2_U2443 & P2_U4650); 
assign P2_U3286 = ~(P2_U3253 & P2_U2616); 
assign P2_U3325 = ~(P2_U3312 & P2_U4651); 
assign P2_U3355 = ~(P2_U3350 & P2_U4770); 
assign P2_U3716 = P2_U4624 & P2_U3304; 
assign P2_U4057 = P2_U2616 & P2_U4468; 
assign P2_U4189 = P2_U2374 & P2_U3253; 
assign P2_U4259 = P2_U7802 & P2_U7786 & P2_U7770 & P2_U7754; 
assign P2_U4260 = P2_U7874 & P2_U7850 & P2_U7834 & P2_U7818; 
assign P2_U4261 = P2_U7803 & P2_U7787 & P2_U7771 & P2_U7755; 
assign P2_U4262 = P2_U7875 & P2_U7851 & P2_U7835 & P2_U7819; 
assign P2_U4263 = P2_U7804 & P2_U7788 & P2_U7772 & P2_U7756; 
assign P2_U4264 = P2_U7876 & P2_U7852 & P2_U7836 & P2_U7820; 
assign P2_U4265 = P2_U7805 & P2_U7789 & P2_U7773 & P2_U7757; 
assign P2_U4266 = P2_U7877 & P2_U7853 & P2_U7837 & P2_U7821; 
assign P2_U4267 = P2_U7806 & P2_U7790 & P2_U7774 & P2_U7758; 
assign P2_U4268 = P2_U7878 & P2_U7854 & P2_U7838 & P2_U7822; 
assign P2_U4269 = P2_U7807 & P2_U7791 & P2_U7775 & P2_U7759; 
assign P2_U4270 = P2_U7879 & P2_U7855 & P2_U7839 & P2_U7823; 
assign P2_U4271 = P2_U7808 & P2_U7792 & P2_U7776 & P2_U7760; 
assign P2_U4272 = P2_U7880 & P2_U7856 & P2_U7840 & P2_U7824; 
assign P2_U4273 = P2_U7809 & P2_U7793 & P2_U7777 & P2_U7761; 
assign P2_U4274 = P2_U7881 & P2_U7857 & P2_U7841 & P2_U7825; 
assign P2_U4337 = P2_U2616 & P2_U3300; 
assign P2_U4579 = ~(P2_U4573 & P2_STATE_REG_2__SCAN_IN); 
assign P2_U4712 = ~P2_U3245; 
assign P2_U4828 = ~P2_U3246; 
assign P2_U4885 = ~(P2_U2442 & P2_U2444); 
assign P2_U5000 = ~(P2_U2442 & P2_U2445); 
assign P2_U5114 = ~(P2_U2441 & P2_U2444); 
assign P2_U5228 = ~(P2_U2441 & P2_U2445); 
assign P2_U5343 = ~(P2_U2443 & P2_U2444); 
assign P2_U5458 = ~(P2_U2443 & P2_U2445); 
assign P2_U5598 = ~(P2_U2617 & P2_U3521); 
assign P2_U6133 = ~(U211 & P2_U2616); 
assign P2_U6836 = ~(P2_U4477 & P2_REIP_REG_0__SCAN_IN); 
assign P2_U6862 = ~(P2_U2538 & P2_INSTQUEUE_REG_8__7__SCAN_IN); 
assign P2_U6863 = ~(P2_U2537 & P2_INSTQUEUE_REG_9__7__SCAN_IN); 
assign P2_U6864 = ~(P2_U2536 & P2_INSTQUEUE_REG_10__7__SCAN_IN); 
assign P2_U6865 = ~(P2_U2535 & P2_INSTQUEUE_REG_11__7__SCAN_IN); 
assign P2_U6866 = ~(P2_U2534 & P2_INSTQUEUE_REG_12__7__SCAN_IN); 
assign P2_U6867 = ~(P2_U2533 & P2_INSTQUEUE_REG_13__7__SCAN_IN); 
assign P2_U6868 = ~(P2_U2531 & P2_INSTQUEUE_REG_14__7__SCAN_IN); 
assign P2_U6869 = ~(P2_U2530 & P2_INSTQUEUE_REG_15__7__SCAN_IN); 
assign P2_U6878 = ~(P2_U2562 & P2_INSTQUEUE_REG_15__7__SCAN_IN); 
assign P2_U6879 = ~(P2_U2561 & P2_INSTQUEUE_REG_14__7__SCAN_IN); 
assign P2_U6880 = ~(P2_U2560 & P2_INSTQUEUE_REG_13__7__SCAN_IN); 
assign P2_U6881 = ~(P2_U2559 & P2_INSTQUEUE_REG_12__7__SCAN_IN); 
assign P2_U6882 = ~(P2_U2558 & P2_INSTQUEUE_REG_11__7__SCAN_IN); 
assign P2_U6883 = ~(P2_U2557 & P2_INSTQUEUE_REG_10__7__SCAN_IN); 
assign P2_U6884 = ~(P2_U2555 & P2_INSTQUEUE_REG_9__7__SCAN_IN); 
assign P2_U6885 = ~(P2_U2554 & P2_INSTQUEUE_REG_8__7__SCAN_IN); 
assign P2_U6888 = ~(P2_U2550 & P2_INSTQUEUE_REG_5__7__SCAN_IN); 
assign P2_U6889 = ~(P2_U2548 & P2_INSTQUEUE_REG_4__7__SCAN_IN); 
assign P2_U6892 = ~(P2_U2543 & P2_INSTQUEUE_REG_1__7__SCAN_IN); 
assign P2_U6893 = ~(P2_U2541 & P2_INSTQUEUE_REG_0__7__SCAN_IN); 
assign P2_U6894 = ~(P2_U2562 & P2_INSTQUEUE_REG_15__6__SCAN_IN); 
assign P2_U6895 = ~(P2_U2561 & P2_INSTQUEUE_REG_14__6__SCAN_IN); 
assign P2_U6896 = ~(P2_U2560 & P2_INSTQUEUE_REG_13__6__SCAN_IN); 
assign P2_U6897 = ~(P2_U2559 & P2_INSTQUEUE_REG_12__6__SCAN_IN); 
assign P2_U6898 = ~(P2_U2558 & P2_INSTQUEUE_REG_11__6__SCAN_IN); 
assign P2_U6899 = ~(P2_U2557 & P2_INSTQUEUE_REG_10__6__SCAN_IN); 
assign P2_U6900 = ~(P2_U2555 & P2_INSTQUEUE_REG_9__6__SCAN_IN); 
assign P2_U6901 = ~(P2_U2554 & P2_INSTQUEUE_REG_8__6__SCAN_IN); 
assign P2_U6904 = ~(P2_U2550 & P2_INSTQUEUE_REG_5__6__SCAN_IN); 
assign P2_U6905 = ~(P2_U2548 & P2_INSTQUEUE_REG_4__6__SCAN_IN); 
assign P2_U6908 = ~(P2_U2543 & P2_INSTQUEUE_REG_1__6__SCAN_IN); 
assign P2_U6909 = ~(P2_U2541 & P2_INSTQUEUE_REG_0__6__SCAN_IN); 
assign P2_U6910 = ~(P2_U2562 & P2_INSTQUEUE_REG_15__5__SCAN_IN); 
assign P2_U6911 = ~(P2_U2561 & P2_INSTQUEUE_REG_14__5__SCAN_IN); 
assign P2_U6912 = ~(P2_U2560 & P2_INSTQUEUE_REG_13__5__SCAN_IN); 
assign P2_U6913 = ~(P2_U2559 & P2_INSTQUEUE_REG_12__5__SCAN_IN); 
assign P2_U6914 = ~(P2_U2558 & P2_INSTQUEUE_REG_11__5__SCAN_IN); 
assign P2_U6915 = ~(P2_U2557 & P2_INSTQUEUE_REG_10__5__SCAN_IN); 
assign P2_U6916 = ~(P2_U2555 & P2_INSTQUEUE_REG_9__5__SCAN_IN); 
assign P2_U6917 = ~(P2_U2554 & P2_INSTQUEUE_REG_8__5__SCAN_IN); 
assign P2_U6920 = ~(P2_U2550 & P2_INSTQUEUE_REG_5__5__SCAN_IN); 
assign P2_U6921 = ~(P2_U2548 & P2_INSTQUEUE_REG_4__5__SCAN_IN); 
assign P2_U6924 = ~(P2_U2543 & P2_INSTQUEUE_REG_1__5__SCAN_IN); 
assign P2_U6925 = ~(P2_U2541 & P2_INSTQUEUE_REG_0__5__SCAN_IN); 
assign P2_U6926 = ~(P2_U2562 & P2_INSTQUEUE_REG_15__4__SCAN_IN); 
assign P2_U6927 = ~(P2_U2561 & P2_INSTQUEUE_REG_14__4__SCAN_IN); 
assign P2_U6928 = ~(P2_U2560 & P2_INSTQUEUE_REG_13__4__SCAN_IN); 
assign P2_U6929 = ~(P2_U2559 & P2_INSTQUEUE_REG_12__4__SCAN_IN); 
assign P2_U6930 = ~(P2_U2558 & P2_INSTQUEUE_REG_11__4__SCAN_IN); 
assign P2_U6931 = ~(P2_U2557 & P2_INSTQUEUE_REG_10__4__SCAN_IN); 
assign P2_U6932 = ~(P2_U2555 & P2_INSTQUEUE_REG_9__4__SCAN_IN); 
assign P2_U6933 = ~(P2_U2554 & P2_INSTQUEUE_REG_8__4__SCAN_IN); 
assign P2_U6936 = ~(P2_U2550 & P2_INSTQUEUE_REG_5__4__SCAN_IN); 
assign P2_U6937 = ~(P2_U2548 & P2_INSTQUEUE_REG_4__4__SCAN_IN); 
assign P2_U6940 = ~(P2_U2543 & P2_INSTQUEUE_REG_1__4__SCAN_IN); 
assign P2_U6941 = ~(P2_U2541 & P2_INSTQUEUE_REG_0__4__SCAN_IN); 
assign P2_U6942 = ~(P2_U2562 & P2_INSTQUEUE_REG_15__3__SCAN_IN); 
assign P2_U6943 = ~(P2_U2561 & P2_INSTQUEUE_REG_14__3__SCAN_IN); 
assign P2_U6944 = ~(P2_U2560 & P2_INSTQUEUE_REG_13__3__SCAN_IN); 
assign P2_U6945 = ~(P2_U2559 & P2_INSTQUEUE_REG_12__3__SCAN_IN); 
assign P2_U6946 = ~(P2_U2558 & P2_INSTQUEUE_REG_11__3__SCAN_IN); 
assign P2_U6947 = ~(P2_U2557 & P2_INSTQUEUE_REG_10__3__SCAN_IN); 
assign P2_U6948 = ~(P2_U2555 & P2_INSTQUEUE_REG_9__3__SCAN_IN); 
assign P2_U6949 = ~(P2_U2554 & P2_INSTQUEUE_REG_8__3__SCAN_IN); 
assign P2_U6952 = ~(P2_U2550 & P2_INSTQUEUE_REG_5__3__SCAN_IN); 
assign P2_U6953 = ~(P2_U2548 & P2_INSTQUEUE_REG_4__3__SCAN_IN); 
assign P2_U6956 = ~(P2_U2543 & P2_INSTQUEUE_REG_1__3__SCAN_IN); 
assign P2_U6957 = ~(P2_U2541 & P2_INSTQUEUE_REG_0__3__SCAN_IN); 
assign P2_U6958 = ~(P2_U2562 & P2_INSTQUEUE_REG_15__2__SCAN_IN); 
assign P2_U6959 = ~(P2_U2561 & P2_INSTQUEUE_REG_14__2__SCAN_IN); 
assign P2_U6960 = ~(P2_U2560 & P2_INSTQUEUE_REG_13__2__SCAN_IN); 
assign P2_U6961 = ~(P2_U2559 & P2_INSTQUEUE_REG_12__2__SCAN_IN); 
assign P2_U6962 = ~(P2_U2558 & P2_INSTQUEUE_REG_11__2__SCAN_IN); 
assign P2_U6963 = ~(P2_U2557 & P2_INSTQUEUE_REG_10__2__SCAN_IN); 
assign P2_U6964 = ~(P2_U2555 & P2_INSTQUEUE_REG_9__2__SCAN_IN); 
assign P2_U6965 = ~(P2_U2554 & P2_INSTQUEUE_REG_8__2__SCAN_IN); 
assign P2_U6968 = ~(P2_U2550 & P2_INSTQUEUE_REG_5__2__SCAN_IN); 
assign P2_U6969 = ~(P2_U2548 & P2_INSTQUEUE_REG_4__2__SCAN_IN); 
assign P2_U6972 = ~(P2_U2543 & P2_INSTQUEUE_REG_1__2__SCAN_IN); 
assign P2_U6973 = ~(P2_U2541 & P2_INSTQUEUE_REG_0__2__SCAN_IN); 
assign P2_U6974 = ~(P2_U2562 & P2_INSTQUEUE_REG_15__1__SCAN_IN); 
assign P2_U6975 = ~(P2_U2561 & P2_INSTQUEUE_REG_14__1__SCAN_IN); 
assign P2_U6976 = ~(P2_U2560 & P2_INSTQUEUE_REG_13__1__SCAN_IN); 
assign P2_U6977 = ~(P2_U2559 & P2_INSTQUEUE_REG_12__1__SCAN_IN); 
assign P2_U6978 = ~(P2_U2558 & P2_INSTQUEUE_REG_11__1__SCAN_IN); 
assign P2_U6979 = ~(P2_U2557 & P2_INSTQUEUE_REG_10__1__SCAN_IN); 
assign P2_U6980 = ~(P2_U2555 & P2_INSTQUEUE_REG_9__1__SCAN_IN); 
assign P2_U6981 = ~(P2_U2554 & P2_INSTQUEUE_REG_8__1__SCAN_IN); 
assign P2_U6984 = ~(P2_U2550 & P2_INSTQUEUE_REG_5__1__SCAN_IN); 
assign P2_U6985 = ~(P2_U2548 & P2_INSTQUEUE_REG_4__1__SCAN_IN); 
assign P2_U6988 = ~(P2_U2543 & P2_INSTQUEUE_REG_1__1__SCAN_IN); 
assign P2_U6989 = ~(P2_U2541 & P2_INSTQUEUE_REG_0__1__SCAN_IN); 
assign P2_U6990 = ~(P2_U2562 & P2_INSTQUEUE_REG_15__0__SCAN_IN); 
assign P2_U6991 = ~(P2_U2561 & P2_INSTQUEUE_REG_14__0__SCAN_IN); 
assign P2_U6992 = ~(P2_U2560 & P2_INSTQUEUE_REG_13__0__SCAN_IN); 
assign P2_U6993 = ~(P2_U2559 & P2_INSTQUEUE_REG_12__0__SCAN_IN); 
assign P2_U6994 = ~(P2_U2558 & P2_INSTQUEUE_REG_11__0__SCAN_IN); 
assign P2_U6995 = ~(P2_U2557 & P2_INSTQUEUE_REG_10__0__SCAN_IN); 
assign P2_U6996 = ~(P2_U2555 & P2_INSTQUEUE_REG_9__0__SCAN_IN); 
assign P2_U6997 = ~(P2_U2554 & P2_INSTQUEUE_REG_8__0__SCAN_IN); 
assign P2_U7000 = ~(P2_U2550 & P2_INSTQUEUE_REG_5__0__SCAN_IN); 
assign P2_U7001 = ~(P2_U2548 & P2_INSTQUEUE_REG_4__0__SCAN_IN); 
assign P2_U7004 = ~(P2_U2543 & P2_INSTQUEUE_REG_1__0__SCAN_IN); 
assign P2_U7005 = ~(P2_U2541 & P2_INSTQUEUE_REG_0__0__SCAN_IN); 
assign P2_U7201 = ~(P2_U2538 & P2_INSTQUEUE_REG_8__6__SCAN_IN); 
assign P2_U7202 = ~(P2_U2537 & P2_INSTQUEUE_REG_9__6__SCAN_IN); 
assign P2_U7203 = ~(P2_U2536 & P2_INSTQUEUE_REG_10__6__SCAN_IN); 
assign P2_U7204 = ~(P2_U2535 & P2_INSTQUEUE_REG_11__6__SCAN_IN); 
assign P2_U7205 = ~(P2_U2534 & P2_INSTQUEUE_REG_12__6__SCAN_IN); 
assign P2_U7206 = ~(P2_U2533 & P2_INSTQUEUE_REG_13__6__SCAN_IN); 
assign P2_U7207 = ~(P2_U2531 & P2_INSTQUEUE_REG_14__6__SCAN_IN); 
assign P2_U7208 = ~(P2_U2530 & P2_INSTQUEUE_REG_15__6__SCAN_IN); 
assign P2_U7235 = ~(P2_U2538 & P2_INSTQUEUE_REG_8__5__SCAN_IN); 
assign P2_U7236 = ~(P2_U2537 & P2_INSTQUEUE_REG_9__5__SCAN_IN); 
assign P2_U7237 = ~(P2_U2536 & P2_INSTQUEUE_REG_10__5__SCAN_IN); 
assign P2_U7238 = ~(P2_U2535 & P2_INSTQUEUE_REG_11__5__SCAN_IN); 
assign P2_U7239 = ~(P2_U2534 & P2_INSTQUEUE_REG_12__5__SCAN_IN); 
assign P2_U7240 = ~(P2_U2533 & P2_INSTQUEUE_REG_13__5__SCAN_IN); 
assign P2_U7241 = ~(P2_U2531 & P2_INSTQUEUE_REG_14__5__SCAN_IN); 
assign P2_U7242 = ~(P2_U2530 & P2_INSTQUEUE_REG_15__5__SCAN_IN); 
assign P2_U7269 = ~(P2_U2538 & P2_INSTQUEUE_REG_8__4__SCAN_IN); 
assign P2_U7270 = ~(P2_U2537 & P2_INSTQUEUE_REG_9__4__SCAN_IN); 
assign P2_U7271 = ~(P2_U2536 & P2_INSTQUEUE_REG_10__4__SCAN_IN); 
assign P2_U7272 = ~(P2_U2535 & P2_INSTQUEUE_REG_11__4__SCAN_IN); 
assign P2_U7273 = ~(P2_U2534 & P2_INSTQUEUE_REG_12__4__SCAN_IN); 
assign P2_U7274 = ~(P2_U2533 & P2_INSTQUEUE_REG_13__4__SCAN_IN); 
assign P2_U7275 = ~(P2_U2531 & P2_INSTQUEUE_REG_14__4__SCAN_IN); 
assign P2_U7276 = ~(P2_U2530 & P2_INSTQUEUE_REG_15__4__SCAN_IN); 
assign P2_U7303 = ~(P2_U2538 & P2_INSTQUEUE_REG_8__3__SCAN_IN); 
assign P2_U7304 = ~(P2_U2537 & P2_INSTQUEUE_REG_9__3__SCAN_IN); 
assign P2_U7305 = ~(P2_U2536 & P2_INSTQUEUE_REG_10__3__SCAN_IN); 
assign P2_U7306 = ~(P2_U2535 & P2_INSTQUEUE_REG_11__3__SCAN_IN); 
assign P2_U7307 = ~(P2_U2534 & P2_INSTQUEUE_REG_12__3__SCAN_IN); 
assign P2_U7308 = ~(P2_U2533 & P2_INSTQUEUE_REG_13__3__SCAN_IN); 
assign P2_U7309 = ~(P2_U2531 & P2_INSTQUEUE_REG_14__3__SCAN_IN); 
assign P2_U7310 = ~(P2_U2530 & P2_INSTQUEUE_REG_15__3__SCAN_IN); 
assign P2_U7337 = ~(P2_U2538 & P2_INSTQUEUE_REG_8__2__SCAN_IN); 
assign P2_U7338 = ~(P2_U2537 & P2_INSTQUEUE_REG_9__2__SCAN_IN); 
assign P2_U7339 = ~(P2_U2536 & P2_INSTQUEUE_REG_10__2__SCAN_IN); 
assign P2_U7340 = ~(P2_U2535 & P2_INSTQUEUE_REG_11__2__SCAN_IN); 
assign P2_U7341 = ~(P2_U2534 & P2_INSTQUEUE_REG_12__2__SCAN_IN); 
assign P2_U7342 = ~(P2_U2533 & P2_INSTQUEUE_REG_13__2__SCAN_IN); 
assign P2_U7343 = ~(P2_U2531 & P2_INSTQUEUE_REG_14__2__SCAN_IN); 
assign P2_U7344 = ~(P2_U2530 & P2_INSTQUEUE_REG_15__2__SCAN_IN); 
assign P2_U7371 = ~(P2_U2538 & P2_INSTQUEUE_REG_8__1__SCAN_IN); 
assign P2_U7372 = ~(P2_U2537 & P2_INSTQUEUE_REG_9__1__SCAN_IN); 
assign P2_U7373 = ~(P2_U2536 & P2_INSTQUEUE_REG_10__1__SCAN_IN); 
assign P2_U7374 = ~(P2_U2535 & P2_INSTQUEUE_REG_11__1__SCAN_IN); 
assign P2_U7375 = ~(P2_U2534 & P2_INSTQUEUE_REG_12__1__SCAN_IN); 
assign P2_U7376 = ~(P2_U2533 & P2_INSTQUEUE_REG_13__1__SCAN_IN); 
assign P2_U7377 = ~(P2_U2531 & P2_INSTQUEUE_REG_14__1__SCAN_IN); 
assign P2_U7378 = ~(P2_U2530 & P2_INSTQUEUE_REG_15__1__SCAN_IN); 
assign P2_U7405 = ~(P2_U2538 & P2_INSTQUEUE_REG_8__0__SCAN_IN); 
assign P2_U7406 = ~(P2_U2537 & P2_INSTQUEUE_REG_9__0__SCAN_IN); 
assign P2_U7407 = ~(P2_U2536 & P2_INSTQUEUE_REG_10__0__SCAN_IN); 
assign P2_U7408 = ~(P2_U2535 & P2_INSTQUEUE_REG_11__0__SCAN_IN); 
assign P2_U7409 = ~(P2_U2534 & P2_INSTQUEUE_REG_12__0__SCAN_IN); 
assign P2_U7410 = ~(P2_U2533 & P2_INSTQUEUE_REG_13__0__SCAN_IN); 
assign P2_U7411 = ~(P2_U2531 & P2_INSTQUEUE_REG_14__0__SCAN_IN); 
assign P2_U7412 = ~(P2_U2530 & P2_INSTQUEUE_REG_15__0__SCAN_IN); 
assign P2_U7859 = ~P2_U3280; 
assign P2_U7861 = ~P2_U3279; 
assign P2_U7863 = ~P2_U3278; 
assign P2_U7865 = ~P2_U3521; 
assign P2_U7867 = ~P2_U3255; 
assign P2_U7869 = ~P2_U2617; 
assign P2_U7871 = ~P2_U3253; 
assign P2_U7873 = ~P2_U2616; 
assign P2_U7914 = ~(P2_U4584 & P2_U3244); 
assign P2_U7918 = ~(P2_U7917 & P2_DATAWIDTH_REG_0__SCAN_IN); 
assign P2_U7921 = ~(P2_U7917 & P2_DATAWIDTH_REG_1__SCAN_IN); 
assign P2_U8116 = ~(P2_U2359 & P2_U3280 & P2_U2616); 
assign P2_U8135 = ~(P2_U7917 & P2_STATEBS16_REG_SCAN_IN); 
assign P2_U8369 = ~(P2_R2337_U65 & P2_U3284); 
assign P2_U8431 = ~(P2_R2238_U22 & P2_U3269); 
assign P1_U2452 = P1_U4400 & P1_U3277 & P1_U3391 & P1_U4173; 
assign P1_U2523 = P1_U2522 & P1_U2521; 
assign P1_U2525 = P1_U2522 & P1_U2524; 
assign P1_U2527 = P1_U2522 & P1_U2526; 
assign P1_U2529 = P1_U2522 & P1_U2528; 
assign P1_U2531 = P1_U2530 & P1_U2521; 
assign P1_U2532 = P1_U2530 & P1_U2524; 
assign P1_U2533 = P1_U2530 & P1_U2526; 
assign P1_U2534 = P1_U2530 & P1_U2528; 
assign P1_U2545 = P1_U5480 & P1_U7720; 
assign P1_U2550 = P1_U5480 & P1_U3456; 
assign P1_U2556 = P1_U2555 & P1_U2454; 
assign P1_U2557 = P1_U2555 & P1_U3498; 
assign P1_U2558 = P1_U2555 & P1_U4378; 
assign P1_U2559 = P1_U2555 & P1_U2456; 
assign P1_U2561 = P1_U2560 & P1_U2454; 
assign P1_U2562 = P1_U2560 & P1_U3498; 
assign P1_U2563 = P1_U2560 & P1_U4378; 
assign P1_U2564 = P1_U2560 & P1_U2456; 
assign P1_U2583 = P1_U7790 & P1_U4184; 
assign P1_U2588 = P1_U7790 & P1_U3452; 
assign P1_U2594 = P1_U2593 & P1_U2524; 
assign P1_U2595 = P1_U2593 & P1_U2521; 
assign P1_U2596 = P1_U2593 & P1_U2528; 
assign P1_U2597 = P1_U2593 & P1_U2526; 
assign P1_U2599 = P1_U2598 & P1_U2524; 
assign P1_U2600 = P1_U2598 & P1_U2521; 
assign P1_U2601 = P1_U2598 & P1_U2528; 
assign P1_U2602 = P1_U2598 & P1_U2526; 
assign P1_U2802 = ~(P1_U7650 & P1_U6613); 
assign P1_U3164 = P1_U7650 & P1_DATAWIDTH_REG_31__SCAN_IN; 
assign P1_U3165 = P1_U7650 & P1_DATAWIDTH_REG_30__SCAN_IN; 
assign P1_U3166 = P1_U7650 & P1_DATAWIDTH_REG_29__SCAN_IN; 
assign P1_U3167 = P1_U7650 & P1_DATAWIDTH_REG_28__SCAN_IN; 
assign P1_U3168 = P1_U7650 & P1_DATAWIDTH_REG_27__SCAN_IN; 
assign P1_U3169 = P1_U7650 & P1_DATAWIDTH_REG_26__SCAN_IN; 
assign P1_U3170 = P1_U7650 & P1_DATAWIDTH_REG_25__SCAN_IN; 
assign P1_U3171 = P1_U7650 & P1_DATAWIDTH_REG_24__SCAN_IN; 
assign P1_U3172 = P1_U7650 & P1_DATAWIDTH_REG_23__SCAN_IN; 
assign P1_U3173 = P1_U7650 & P1_DATAWIDTH_REG_22__SCAN_IN; 
assign P1_U3174 = P1_U7650 & P1_DATAWIDTH_REG_21__SCAN_IN; 
assign P1_U3175 = P1_U7650 & P1_DATAWIDTH_REG_20__SCAN_IN; 
assign P1_U3176 = P1_U7650 & P1_DATAWIDTH_REG_19__SCAN_IN; 
assign P1_U3177 = P1_U7650 & P1_DATAWIDTH_REG_18__SCAN_IN; 
assign P1_U3178 = P1_U7650 & P1_DATAWIDTH_REG_17__SCAN_IN; 
assign P1_U3179 = P1_U7650 & P1_DATAWIDTH_REG_16__SCAN_IN; 
assign P1_U3180 = P1_U7650 & P1_DATAWIDTH_REG_15__SCAN_IN; 
assign P1_U3181 = P1_U7650 & P1_DATAWIDTH_REG_14__SCAN_IN; 
assign P1_U3182 = P1_U7650 & P1_DATAWIDTH_REG_13__SCAN_IN; 
assign P1_U3183 = P1_U7650 & P1_DATAWIDTH_REG_12__SCAN_IN; 
assign P1_U3184 = P1_U7650 & P1_DATAWIDTH_REG_11__SCAN_IN; 
assign P1_U3185 = P1_U7650 & P1_DATAWIDTH_REG_10__SCAN_IN; 
assign P1_U3186 = P1_U7650 & P1_DATAWIDTH_REG_9__SCAN_IN; 
assign P1_U3187 = P1_U7650 & P1_DATAWIDTH_REG_8__SCAN_IN; 
assign P1_U3188 = P1_U7650 & P1_DATAWIDTH_REG_7__SCAN_IN; 
assign P1_U3189 = P1_U7650 & P1_DATAWIDTH_REG_6__SCAN_IN; 
assign P1_U3190 = P1_U7650 & P1_DATAWIDTH_REG_5__SCAN_IN; 
assign P1_U3191 = P1_U7650 & P1_DATAWIDTH_REG_4__SCAN_IN; 
assign P1_U3192 = P1_U7650 & P1_DATAWIDTH_REG_3__SCAN_IN; 
assign P1_U3193 = P1_U7650 & P1_DATAWIDTH_REG_2__SCAN_IN; 
assign P1_U3195 = ~(P1_U7645 & P1_U7644 & P1_U3495); 
assign P1_U3197 = ~(P1_U4355 & P1_U4354 & P1_U4356); 
assign P1_U3198 = ~(P1_U4352 & P1_U4351 & P1_U4353); 
assign P1_U3199 = ~(P1_U4349 & P1_U4348 & P1_U4350); 
assign P1_U3200 = ~(P1_U4346 & P1_U4345 & P1_U4347); 
assign P1_U3201 = ~(P1_U4343 & P1_U4342 & P1_U4344); 
assign P1_U3202 = ~(P1_U4340 & P1_U4339 & P1_U4341); 
assign P1_U3203 = ~(P1_U4337 & P1_U4336 & P1_U4338); 
assign P1_U3204 = ~(P1_U4334 & P1_U4333 & P1_U4335); 
assign P1_U3205 = ~(P1_U4331 & P1_U4330 & P1_U4332); 
assign P1_U3206 = ~(P1_U4328 & P1_U4327 & P1_U4329); 
assign P1_U3207 = ~(P1_U4325 & P1_U4324 & P1_U4326); 
assign P1_U3208 = ~(P1_U4322 & P1_U4321 & P1_U4323); 
assign P1_U3209 = ~(P1_U4319 & P1_U4318 & P1_U4320); 
assign P1_U3210 = ~(P1_U4316 & P1_U4315 & P1_U4317); 
assign P1_U3211 = ~(P1_U4313 & P1_U4312 & P1_U4314); 
assign P1_U3212 = ~(P1_U4310 & P1_U4309 & P1_U4311); 
assign P1_U3213 = ~(P1_U4307 & P1_U4306 & P1_U4308); 
assign P1_U3214 = ~(P1_U4304 & P1_U4303 & P1_U4305); 
assign P1_U3215 = ~(P1_U4301 & P1_U4300 & P1_U4302); 
assign P1_U3216 = ~(P1_U4298 & P1_U4297 & P1_U4299); 
assign P1_U3217 = ~(P1_U4295 & P1_U4294 & P1_U4296); 
assign P1_U3218 = ~(P1_U4292 & P1_U4291 & P1_U4293); 
assign P1_U3219 = ~(P1_U4289 & P1_U4288 & P1_U4290); 
assign P1_U3220 = ~(P1_U4286 & P1_U4285 & P1_U4287); 
assign P1_U3221 = ~(P1_U4283 & P1_U4282 & P1_U4284); 
assign P1_U3222 = ~(P1_U4280 & P1_U4279 & P1_U4281); 
assign P1_U3223 = ~(P1_U4277 & P1_U4276 & P1_U4278); 
assign P1_U3224 = ~(P1_U4274 & P1_U4273 & P1_U4275); 
assign P1_U3225 = ~(P1_U4271 & P1_U4270 & P1_U4272); 
assign P1_U3226 = ~(P1_U4268 & P1_U4267 & P1_U4269); 
assign P1_U3238 = ~(P1_U2434 & P1_U3235); 
assign P1_U3239 = ~(P1_U2434 & P1_U4543); 
assign P1_U3240 = ~(P1_U2433 & P1_U3235); 
assign P1_U3241 = ~(P1_U2433 & P1_U4543); 
assign P1_U3242 = ~(P1_U2435 & P1_U3235); 
assign P1_U3243 = ~(P1_U2435 & P1_U4543); 
assign P1_U3290 = ~(P1_U3271 & P1_U3283); 
assign P1_U3322 = ~(P1_U3306 & P1_U4544); 
assign P1_U3336 = ~(P1_U3330 & P1_U4663); 
assign P1_U3389 = ~(P1_U3284 & P1_U3278); 
assign P1_U3390 = ~(P1_U3284 & P1_U3271); 
assign P1_U3394 = ~(P1_U2605 & P1_U3277); 
assign P1_U3405 = ~(P1_U3278 & P1_U3284 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U3407 = ~(P1_U3277 & P1_U3391); 
assign P1_U3412 = ~(P1_U3271 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U3481 = ~(P1_U7755 & P1_U7754); 
assign P1_U3865 = P1_U2368 & P1_U3284; 
assign P1_U3884 = P1_U2605 & P1_U3391; 
assign P1_U4063 = P1_U7069 & P1_U7068 & P1_U7067 & P1_U7066; 
assign P1_U4066 = P1_U7081 & P1_U7080 & P1_U7079 & P1_U7078; 
assign P1_U4072 = P1_U4400 & P1_U3391; 
assign P1_U4073 = P1_U3284 & P1_STATE2_REG_0__SCAN_IN; 
assign P1_U4079 = P1_U7101 & P1_U7100 & P1_U7099 & P1_U7098; 
assign P1_U4082 = P1_U7113 & P1_U7112 & P1_U7111 & P1_U7110; 
assign P1_U4083 = P1_U7118 & P1_U7117 & P1_U7116 & P1_U7115; 
assign P1_U4086 = P1_U7130 & P1_U7129 & P1_U7128 & P1_U7127; 
assign P1_U4087 = P1_U7135 & P1_U7134 & P1_U7133 & P1_U7132; 
assign P1_U4090 = P1_U7145 & P1_U7144; 
assign P1_U4092 = P1_U7150 & P1_U7149 & P1_U7148 & P1_U7147; 
assign P1_U4095 = P1_U7162 & P1_U7161 & P1_U7160 & P1_U7159; 
assign P1_U4096 = P1_U7167 & P1_U7166 & P1_U7165 & P1_U7164; 
assign P1_U4099 = P1_U7179 & P1_U7178 & P1_U7177 & P1_U7176; 
assign P1_U4100 = P1_U7184 & P1_U7183 & P1_U7182 & P1_U7181; 
assign P1_U4103 = P1_U7196 & P1_U7195 & P1_U7194 & P1_U7193; 
assign P1_U4104 = P1_U7201 & P1_U7200 & P1_U7199 & P1_U7198; 
assign P1_U4107 = P1_U7213 & P1_U7212 & P1_U7211 & P1_U7210; 
assign P1_U4154 = P1_U3283 & P1_U3391; 
assign P1_U4159 = P1_U3271 & P1_U4173; 
assign P1_U4168 = P1_U7462 & P1_U7461; 
assign P1_U4251 = ~P1_U3415; 
assign P1_U4265 = ~P1_U3453; 
assign P1_U4369 = ~(P1_U4363 & P1_STATE_REG_2__SCAN_IN); 
assign P1_U4399 = ~P1_U3283; 
assign P1_U4432 = ~P1_U4171; 
assign P1_U4449 = ~P1_U3391; 
assign P1_U4460 = ~P1_U3277; 
assign P1_U4477 = ~P1_U3271; 
assign P1_U4494 = ~P1_U3284; 
assign P1_U4605 = ~P1_U3236; 
assign P1_U4611 = ~(P1_U3236 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U4721 = ~P1_U3237; 
assign P1_U4727 = ~(P1_U3237 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U4778 = ~(P1_U2434 & P1_U2436); 
assign P1_U4893 = ~(P1_U2434 & P1_U2437); 
assign P1_U5007 = ~(P1_U2433 & P1_U2436); 
assign P1_U5121 = ~(P1_U2433 & P1_U2437); 
assign P1_U5236 = ~(P1_U2435 & P1_U2436); 
assign P1_U5351 = ~(P1_U2435 & P1_U2437); 
assign P1_U5526 = ~(P1_U7712 & P1_U2446); 
assign P1_U6618 = ~(P1_U2544 & P1_INSTQUEUE_REG_15__7__SCAN_IN); 
assign P1_U6619 = ~(P1_U2543 & P1_INSTQUEUE_REG_14__7__SCAN_IN); 
assign P1_U6620 = ~(P1_U2542 & P1_INSTQUEUE_REG_13__7__SCAN_IN); 
assign P1_U6621 = ~(P1_U2541 & P1_INSTQUEUE_REG_12__7__SCAN_IN); 
assign P1_U6622 = ~(P1_U2539 & P1_INSTQUEUE_REG_11__7__SCAN_IN); 
assign P1_U6623 = ~(P1_U2538 & P1_INSTQUEUE_REG_10__7__SCAN_IN); 
assign P1_U6624 = ~(P1_U2537 & P1_INSTQUEUE_REG_9__7__SCAN_IN); 
assign P1_U6625 = ~(P1_U2536 & P1_INSTQUEUE_REG_8__7__SCAN_IN); 
assign P1_U6634 = ~(P1_U2544 & P1_INSTQUEUE_REG_15__6__SCAN_IN); 
assign P1_U6635 = ~(P1_U2543 & P1_INSTQUEUE_REG_14__6__SCAN_IN); 
assign P1_U6636 = ~(P1_U2542 & P1_INSTQUEUE_REG_13__6__SCAN_IN); 
assign P1_U6637 = ~(P1_U2541 & P1_INSTQUEUE_REG_12__6__SCAN_IN); 
assign P1_U6638 = ~(P1_U2539 & P1_INSTQUEUE_REG_11__6__SCAN_IN); 
assign P1_U6639 = ~(P1_U2538 & P1_INSTQUEUE_REG_10__6__SCAN_IN); 
assign P1_U6640 = ~(P1_U2537 & P1_INSTQUEUE_REG_9__6__SCAN_IN); 
assign P1_U6641 = ~(P1_U2536 & P1_INSTQUEUE_REG_8__6__SCAN_IN); 
assign P1_U6650 = ~(P1_U2544 & P1_INSTQUEUE_REG_15__5__SCAN_IN); 
assign P1_U6651 = ~(P1_U2543 & P1_INSTQUEUE_REG_14__5__SCAN_IN); 
assign P1_U6652 = ~(P1_U2542 & P1_INSTQUEUE_REG_13__5__SCAN_IN); 
assign P1_U6653 = ~(P1_U2541 & P1_INSTQUEUE_REG_12__5__SCAN_IN); 
assign P1_U6654 = ~(P1_U2539 & P1_INSTQUEUE_REG_11__5__SCAN_IN); 
assign P1_U6655 = ~(P1_U2538 & P1_INSTQUEUE_REG_10__5__SCAN_IN); 
assign P1_U6656 = ~(P1_U2537 & P1_INSTQUEUE_REG_9__5__SCAN_IN); 
assign P1_U6657 = ~(P1_U2536 & P1_INSTQUEUE_REG_8__5__SCAN_IN); 
assign P1_U6666 = ~(P1_U2544 & P1_INSTQUEUE_REG_15__4__SCAN_IN); 
assign P1_U6667 = ~(P1_U2543 & P1_INSTQUEUE_REG_14__4__SCAN_IN); 
assign P1_U6668 = ~(P1_U2542 & P1_INSTQUEUE_REG_13__4__SCAN_IN); 
assign P1_U6669 = ~(P1_U2541 & P1_INSTQUEUE_REG_12__4__SCAN_IN); 
assign P1_U6670 = ~(P1_U2539 & P1_INSTQUEUE_REG_11__4__SCAN_IN); 
assign P1_U6671 = ~(P1_U2538 & P1_INSTQUEUE_REG_10__4__SCAN_IN); 
assign P1_U6672 = ~(P1_U2537 & P1_INSTQUEUE_REG_9__4__SCAN_IN); 
assign P1_U6673 = ~(P1_U2536 & P1_INSTQUEUE_REG_8__4__SCAN_IN); 
assign P1_U6681 = ~(P1_U2544 & P1_INSTQUEUE_REG_15__3__SCAN_IN); 
assign P1_U6682 = ~(P1_U2543 & P1_INSTQUEUE_REG_14__3__SCAN_IN); 
assign P1_U6683 = ~(P1_U2542 & P1_INSTQUEUE_REG_13__3__SCAN_IN); 
assign P1_U6684 = ~(P1_U2541 & P1_INSTQUEUE_REG_12__3__SCAN_IN); 
assign P1_U6685 = ~(P1_U2539 & P1_INSTQUEUE_REG_11__3__SCAN_IN); 
assign P1_U6686 = ~(P1_U2538 & P1_INSTQUEUE_REG_10__3__SCAN_IN); 
assign P1_U6687 = ~(P1_U2537 & P1_INSTQUEUE_REG_9__3__SCAN_IN); 
assign P1_U6688 = ~(P1_U2536 & P1_INSTQUEUE_REG_8__3__SCAN_IN); 
assign P1_U6697 = ~(P1_U2544 & P1_INSTQUEUE_REG_15__2__SCAN_IN); 
assign P1_U6698 = ~(P1_U2543 & P1_INSTQUEUE_REG_14__2__SCAN_IN); 
assign P1_U6699 = ~(P1_U2542 & P1_INSTQUEUE_REG_13__2__SCAN_IN); 
assign P1_U6700 = ~(P1_U2541 & P1_INSTQUEUE_REG_12__2__SCAN_IN); 
assign P1_U6701 = ~(P1_U2539 & P1_INSTQUEUE_REG_11__2__SCAN_IN); 
assign P1_U6702 = ~(P1_U2538 & P1_INSTQUEUE_REG_10__2__SCAN_IN); 
assign P1_U6703 = ~(P1_U2537 & P1_INSTQUEUE_REG_9__2__SCAN_IN); 
assign P1_U6704 = ~(P1_U2536 & P1_INSTQUEUE_REG_8__2__SCAN_IN); 
assign P1_U6713 = ~(P1_U2544 & P1_INSTQUEUE_REG_15__1__SCAN_IN); 
assign P1_U6714 = ~(P1_U2543 & P1_INSTQUEUE_REG_14__1__SCAN_IN); 
assign P1_U6715 = ~(P1_U2542 & P1_INSTQUEUE_REG_13__1__SCAN_IN); 
assign P1_U6716 = ~(P1_U2541 & P1_INSTQUEUE_REG_12__1__SCAN_IN); 
assign P1_U6717 = ~(P1_U2539 & P1_INSTQUEUE_REG_11__1__SCAN_IN); 
assign P1_U6718 = ~(P1_U2538 & P1_INSTQUEUE_REG_10__1__SCAN_IN); 
assign P1_U6719 = ~(P1_U2537 & P1_INSTQUEUE_REG_9__1__SCAN_IN); 
assign P1_U6720 = ~(P1_U2536 & P1_INSTQUEUE_REG_8__1__SCAN_IN); 
assign P1_U6729 = ~(P1_U2544 & P1_INSTQUEUE_REG_15__0__SCAN_IN); 
assign P1_U6730 = ~(P1_U2543 & P1_INSTQUEUE_REG_14__0__SCAN_IN); 
assign P1_U6731 = ~(P1_U2542 & P1_INSTQUEUE_REG_13__0__SCAN_IN); 
assign P1_U6732 = ~(P1_U2541 & P1_INSTQUEUE_REG_12__0__SCAN_IN); 
assign P1_U6733 = ~(P1_U2539 & P1_INSTQUEUE_REG_11__0__SCAN_IN); 
assign P1_U6734 = ~(P1_U2538 & P1_INSTQUEUE_REG_10__0__SCAN_IN); 
assign P1_U6735 = ~(P1_U2537 & P1_INSTQUEUE_REG_9__0__SCAN_IN); 
assign P1_U6736 = ~(P1_U2536 & P1_INSTQUEUE_REG_8__0__SCAN_IN); 
assign P1_U6766 = ~(P1_R2337_U67 & P1_U2352); 
assign P1_U6888 = ~(P1_U2605 & P1_U3284); 
assign P1_U7074 = ~(P1_U2573 & P1_INSTQUEUE_REG_0__7__SCAN_IN); 
assign P1_U7075 = ~(P1_U2572 & P1_INSTQUEUE_REG_1__7__SCAN_IN); 
assign P1_U7076 = ~(P1_U2571 & P1_INSTQUEUE_REG_2__7__SCAN_IN); 
assign P1_U7077 = ~(P1_U2570 & P1_INSTQUEUE_REG_3__7__SCAN_IN); 
assign P1_U7106 = ~(P1_U2573 & P1_INSTQUEUE_REG_0__6__SCAN_IN); 
assign P1_U7107 = ~(P1_U2572 & P1_INSTQUEUE_REG_1__6__SCAN_IN); 
assign P1_U7108 = ~(P1_U2571 & P1_INSTQUEUE_REG_2__6__SCAN_IN); 
assign P1_U7109 = ~(P1_U2570 & P1_INSTQUEUE_REG_3__6__SCAN_IN); 
assign P1_U7123 = ~(P1_U2573 & P1_INSTQUEUE_REG_0__5__SCAN_IN); 
assign P1_U7124 = ~(P1_U2572 & P1_INSTQUEUE_REG_1__5__SCAN_IN); 
assign P1_U7125 = ~(P1_U2571 & P1_INSTQUEUE_REG_2__5__SCAN_IN); 
assign P1_U7126 = ~(P1_U2570 & P1_INSTQUEUE_REG_3__5__SCAN_IN); 
assign P1_U7140 = ~(P1_U2572 & P1_INSTQUEUE_REG_1__4__SCAN_IN); 
assign P1_U7141 = ~(P1_U2571 & P1_INSTQUEUE_REG_2__4__SCAN_IN); 
assign P1_U7142 = ~(P1_U2570 & P1_INSTQUEUE_REG_3__4__SCAN_IN); 
assign P1_U7155 = ~(P1_U2573 & P1_INSTQUEUE_REG_0__3__SCAN_IN); 
assign P1_U7156 = ~(P1_U2572 & P1_INSTQUEUE_REG_1__3__SCAN_IN); 
assign P1_U7157 = ~(P1_U2571 & P1_INSTQUEUE_REG_2__3__SCAN_IN); 
assign P1_U7158 = ~(P1_U2570 & P1_INSTQUEUE_REG_3__3__SCAN_IN); 
assign P1_U7172 = ~(P1_U2573 & P1_INSTQUEUE_REG_0__2__SCAN_IN); 
assign P1_U7173 = ~(P1_U2572 & P1_INSTQUEUE_REG_1__2__SCAN_IN); 
assign P1_U7174 = ~(P1_U2571 & P1_INSTQUEUE_REG_2__2__SCAN_IN); 
assign P1_U7175 = ~(P1_U2570 & P1_INSTQUEUE_REG_3__2__SCAN_IN); 
assign P1_U7189 = ~(P1_U2573 & P1_INSTQUEUE_REG_0__1__SCAN_IN); 
assign P1_U7190 = ~(P1_U2572 & P1_INSTQUEUE_REG_1__1__SCAN_IN); 
assign P1_U7191 = ~(P1_U2571 & P1_INSTQUEUE_REG_2__1__SCAN_IN); 
assign P1_U7192 = ~(P1_U2570 & P1_INSTQUEUE_REG_3__1__SCAN_IN); 
assign P1_U7206 = ~(P1_U2573 & P1_INSTQUEUE_REG_0__0__SCAN_IN); 
assign P1_U7207 = ~(P1_U2572 & P1_INSTQUEUE_REG_1__0__SCAN_IN); 
assign P1_U7208 = ~(P1_U2571 & P1_INSTQUEUE_REG_2__0__SCAN_IN); 
assign P1_U7209 = ~(P1_U2570 & P1_INSTQUEUE_REG_3__0__SCAN_IN); 
assign P1_U7384 = ~(P1_U2450 & P1_U3271); 
assign P1_U7464 = ~(P1_U2446 & P1_U7712 & P1_FLUSH_REG_SCAN_IN); 
assign P1_U7494 = ~P1_U3276; 
assign P1_U7617 = ~(P1_U2573 & P1_INSTQUEUE_REG_0__4__SCAN_IN); 
assign P1_U7647 = ~(P1_U4371 & P1_U3251); 
assign P1_U7651 = ~(P1_U7650 & P1_DATAWIDTH_REG_0__SCAN_IN); 
assign P1_U7654 = ~(P1_U7650 & P1_DATAWIDTH_REG_1__SCAN_IN); 
assign P1_U7704 = ~(P1_U4415 & P1_U3277); 
assign P1_U7705 = ~(P1_U3271 & P1_U3415); 
assign P1_U7764 = ~(P1_U7650 & P1_STATEBS16_REG_SCAN_IN); 
assign P1_U7784 = ~(P1_U2605 & P1_U3277); 
assign P1_U7791 = ~(P1_U3276 & P1_U3284); 
assign P3_ADD_526_U17 = ~(P3_ADD_526_U84 & P3_ADD_526_U118); 
assign P3_ADD_526_U95 = ~(P3_ADD_526_U118 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_526_U145 = ~(P3_ADD_526_U118 & P3_ADD_526_U15); 
assign P3_ADD_526_U148 = ~(P3_ADD_526_U126 & P3_ADD_526_U11); 
assign P3_ADD_552_U17 = ~(P3_ADD_552_U84 & P3_ADD_552_U118); 
assign P3_ADD_552_U95 = ~(P3_ADD_552_U118 & P3_EBX_REG_7__SCAN_IN); 
assign P3_ADD_552_U145 = ~(P3_ADD_552_U118 & P3_ADD_552_U15); 
assign P3_ADD_552_U148 = ~(P3_ADD_552_U126 & P3_ADD_552_U11); 
assign P3_ADD_546_U17 = ~(P3_ADD_546_U84 & P3_ADD_546_U118); 
assign P3_ADD_546_U95 = ~(P3_ADD_546_U118 & P3_EAX_REG_7__SCAN_IN); 
assign P3_ADD_546_U145 = ~(P3_ADD_546_U118 & P3_ADD_546_U15); 
assign P3_ADD_546_U148 = ~(P3_ADD_546_U126 & P3_ADD_546_U11); 
assign P3_GTE_401_U9 = P3_SUB_401_U7 | P3_SUB_401_U22; 
assign P3_ADD_476_U12 = ~(P3_ADD_476_U96 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_476_U132 = ~(P3_ADD_476_U96 & P3_ADD_476_U11); 
assign P3_GTE_390_U9 = P3_SUB_390_U7 | P3_SUB_390_U22; 
assign P3_ADD_531_U13 = ~(P3_ADD_531_U100 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_531_U139 = ~(P3_ADD_531_U100 & P3_ADD_531_U12); 
assign P3_SUB_320_U27 = ~P3_ADD_318_U67; 
assign P3_SUB_320_U59 = P3_SUB_320_U135 & P3_SUB_320_U134; 
assign P3_SUB_320_U92 = ~(P3_ADD_318_U67 & P3_SUB_320_U91); 
assign P3_ADD_505_U6 = P3_ADD_505_U20 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P3_ADD_505_U22 = ~(P3_ADD_505_U20 & P3_ADD_505_U13); 
assign P3_ADD_318_U12 = ~(P3_ADD_318_U96 & P3_PHYADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_318_U132 = ~(P3_ADD_318_U96 & P3_ADD_318_U11); 
assign P3_SUB_370_U34 = ~P3_SUB_370_U28; 
assign P3_SUB_370_U36 = ~(P3_SUB_370_U35 & P3_SUB_370_U28); 
assign P3_SUB_370_U61 = ~(P3_SUB_370_U25 & P3_SUB_370_U28); 
assign P3_ADD_315_U12 = ~(P3_ADD_315_U93 & P3_PHYADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_315_U126 = ~(P3_ADD_315_U93 & P3_ADD_315_U11); 
assign P3_GTE_355_U7 = P3_SUB_355_U7 & P3_SUB_355_U22; 
assign P3_SUB_589_U7 = ~P3_U3302; 
assign P3_ADD_467_U12 = ~(P3_ADD_467_U96 & P3_REIP_REG_5__SCAN_IN); 
assign P3_ADD_467_U132 = ~(P3_ADD_467_U96 & P3_ADD_467_U11); 
assign P3_ADD_430_U12 = ~(P3_ADD_430_U96 & P3_REIP_REG_5__SCAN_IN); 
assign P3_ADD_430_U132 = ~(P3_ADD_430_U96 & P3_ADD_430_U11); 
assign P3_ADD_380_U13 = ~(P3_ADD_380_U100 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_380_U139 = ~(P3_ADD_380_U100 & P3_ADD_380_U12); 
assign P3_GTE_370_U9 = P3_SUB_370_U7 | P3_SUB_370_U22; 
assign P3_ADD_344_U13 = ~(P3_ADD_344_U100 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_344_U139 = ~(P3_ADD_344_U100 & P3_ADD_344_U12); 
assign P3_ADD_339_U12 = ~(P3_ADD_339_U96 & P3_PHYADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_339_U132 = ~(P3_ADD_339_U96 & P3_ADD_339_U11); 
assign P3_ADD_541_U12 = ~(P3_ADD_541_U96 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_541_U132 = ~(P3_ADD_541_U96 & P3_ADD_541_U11); 
assign P3_SUB_355_U34 = ~P3_SUB_355_U28; 
assign P3_SUB_355_U36 = ~(P3_SUB_355_U35 & P3_SUB_355_U28); 
assign P3_SUB_355_U61 = ~(P3_SUB_355_U25 & P3_SUB_355_U28); 
assign P3_SUB_450_U32 = ~P3_SUB_450_U25; 
assign P3_SUB_450_U34 = ~(P3_SUB_450_U33 & P3_SUB_450_U25); 
assign P3_SUB_450_U58 = ~(P3_SUB_450_U22 & P3_SUB_450_U25); 
assign P3_ADD_486_U6 = P3_ADD_486_U20 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P3_ADD_486_U22 = ~(P3_ADD_486_U20 & P3_ADD_486_U13); 
assign P3_SUB_485_U32 = ~P3_SUB_485_U25; 
assign P3_SUB_485_U34 = ~(P3_SUB_485_U33 & P3_SUB_485_U25); 
assign P3_SUB_485_U58 = ~(P3_SUB_485_U22 & P3_SUB_485_U25); 
assign P3_ADD_515_U12 = ~(P3_ADD_515_U96 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_515_U132 = ~(P3_ADD_515_U96 & P3_ADD_515_U11); 
assign P3_ADD_394_U12 = ~(P3_ADD_394_U99 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_394_U136 = ~(P3_ADD_394_U99 & P3_ADD_394_U11); 
assign P3_SUB_414_U19 = P3_SUB_414_U90 & P3_SUB_414_U23; 
assign P3_SUB_414_U24 = ~(P3_SUB_414_U25 & P3_SUB_414_U54 & P3_SUB_414_U85); 
assign P3_SUB_414_U87 = ~(P3_SUB_414_U85 & P3_SUB_414_U54); 
assign P3_SUB_414_U131 = ~(P3_SUB_414_U85 & P3_SUB_414_U54); 
assign P3_ADD_441_U12 = ~(P3_ADD_441_U96 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_441_U132 = ~(P3_ADD_441_U96 & P3_ADD_441_U11); 
assign P3_ADD_349_U13 = ~(P3_ADD_349_U100 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_349_U139 = ~(P3_ADD_349_U100 & P3_ADD_349_U12); 
assign P3_ADD_405_U12 = ~(P3_ADD_405_U99 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_405_U136 = ~(P3_ADD_405_U99 & P3_ADD_405_U11); 
assign P3_ADD_553_U13 = ~(P3_ADD_553_U100 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_553_U139 = ~(P3_ADD_553_U100 & P3_ADD_553_U12); 
assign P3_ADD_558_U13 = ~(P3_ADD_558_U100 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_558_U139 = ~(P3_ADD_558_U100 & P3_ADD_558_U12); 
assign P3_ADD_385_U13 = ~(P3_ADD_385_U100 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_385_U139 = ~(P3_ADD_385_U100 & P3_ADD_385_U12); 
assign P3_ADD_547_U13 = ~(P3_ADD_547_U100 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_547_U139 = ~(P3_ADD_547_U100 & P3_ADD_547_U12); 
assign P3_SUB_412_U32 = ~P3_SUB_412_U25; 
assign P3_SUB_412_U34 = ~(P3_SUB_412_U33 & P3_SUB_412_U25); 
assign P3_SUB_412_U58 = ~(P3_SUB_412_U22 & P3_SUB_412_U25); 
assign P3_SUB_504_U32 = ~P3_SUB_504_U25; 
assign P3_SUB_504_U34 = ~(P3_SUB_504_U33 & P3_SUB_504_U25); 
assign P3_SUB_504_U58 = ~(P3_SUB_504_U22 & P3_SUB_504_U25); 
assign P3_SUB_401_U34 = ~P3_SUB_401_U28; 
assign P3_SUB_401_U36 = ~(P3_SUB_401_U35 & P3_SUB_401_U28); 
assign P3_SUB_401_U61 = ~(P3_SUB_401_U25 & P3_SUB_401_U28); 
assign P3_SUB_390_U34 = ~P3_SUB_390_U28; 
assign P3_SUB_390_U36 = ~(P3_SUB_390_U35 & P3_SUB_390_U28); 
assign P3_SUB_390_U61 = ~(P3_SUB_390_U25 & P3_SUB_390_U28); 
assign P3_ADD_494_U12 = ~(P3_ADD_494_U96 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_494_U132 = ~(P3_ADD_494_U96 & P3_ADD_494_U11); 
assign P3_ADD_536_U12 = ~(P3_ADD_536_U96 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_536_U132 = ~(P3_ADD_536_U96 & P3_ADD_536_U11); 
assign P2_R2027_U13 = ~(P2_R2027_U100 & P2_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P2_R2027_U139 = ~(P2_R2027_U100 & P2_R2027_U12); 
assign P2_R2337_U13 = ~(P2_R2337_U97 & P2_PHYADDRPOINTER_REG_6__SCAN_IN); 
assign P2_R2337_U130 = ~(P2_R2337_U97 & P2_R2337_U12); 
assign P2_R2238_U34 = ~P2_R2238_U28; 
assign P2_R2238_U36 = ~(P2_R2238_U35 & P2_R2238_U28); 
assign P2_R2238_U61 = ~(P2_R2238_U25 & P2_R2238_U28); 
assign P2_R1957_U17 = P2_R1957_U105 & P2_R1957_U21; 
assign P2_R1957_U51 = ~(P2_U3660 | P2_U3658); 
assign P2_R1957_U58 = ~P2_U3660; 
assign P2_R1957_U83 = ~P2_R1957_U21; 
assign P2_R1957_U134 = ~(P2_U3660 & P2_R1957_U21); 
assign P2_SUB_450_U32 = ~P2_SUB_450_U26; 
assign P2_SUB_450_U34 = ~(P2_SUB_450_U33 & P2_SUB_450_U26); 
assign P2_SUB_450_U58 = ~(P2_SUB_450_U23 & P2_SUB_450_U26); 
assign P2_ADD_394_U13 = ~(P2_ADD_394_U99 & P2_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P2_ADD_394_U160 = ~(P2_ADD_394_U99 & P2_ADD_394_U11); 
assign P2_R2267_U42 = ~P2_U2617; 
assign P2_ADD_371_1212_U12 = P2_ADD_371_1212_U8 & P2_ADD_371_1212_U92; 
assign P2_ADD_371_1212_U93 = P2_ADD_371_1212_U8 & P2_ADD_371_1212_U94; 
assign P2_ADD_371_1212_U108 = P2_ADD_371_1212_U8 & P2_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P1_R2027_U17 = ~(P1_R2027_U84 & P1_R2027_U118); 
assign P1_R2027_U95 = ~(P1_R2027_U118 & P1_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P1_R2027_U145 = ~(P1_R2027_U118 & P1_R2027_U15); 
assign P1_R2027_U148 = ~(P1_R2027_U126 & P1_R2027_U11); 
assign P1_R2337_U12 = ~(P1_R2337_U96 & P1_PHYADDRPOINTER_REG_5__SCAN_IN); 
assign P1_R2337_U132 = ~(P1_R2337_U96 & P1_R2337_U11); 
assign P1_R2096_U12 = ~(P1_R2096_U96 & P1_REIP_REG_5__SCAN_IN); 
assign P1_R2096_U132 = ~(P1_R2096_U96 & P1_R2096_U11); 
assign P1_R2238_U34 = ~P1_R2238_U28; 
assign P1_R2238_U36 = ~(P1_R2238_U35 & P1_R2238_U28); 
assign P1_R2238_U61 = ~(P1_R2238_U25 & P1_R2238_U28); 
assign P1_SUB_450_U34 = ~P1_SUB_450_U28; 
assign P1_SUB_450_U36 = ~(P1_SUB_450_U35 & P1_SUB_450_U28); 
assign P1_SUB_450_U61 = ~(P1_SUB_450_U25 & P1_SUB_450_U28); 
assign P1_ADD_405_U13 = ~(P1_ADD_405_U99 & P1_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P1_ADD_405_U160 = ~(P1_ADD_405_U99 & P1_ADD_405_U11); 
assign P1_ADD_515_U13 = ~(P1_ADD_515_U96 & P1_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P1_ADD_515_U158 = ~(P1_ADD_515_U96 & P1_ADD_515_U11); 
assign U389 = ~(U207 & P2_DATAO_REG_0__SCAN_IN); 
assign U391 = ~(U388 & BUF1_REG_0__SCAN_IN); 
assign U392 = ~(U207 & P2_DATAO_REG_1__SCAN_IN); 
assign U394 = ~(U388 & BUF1_REG_1__SCAN_IN); 
assign U395 = ~(U207 & P2_DATAO_REG_2__SCAN_IN); 
assign U397 = ~(U388 & BUF1_REG_2__SCAN_IN); 
assign U398 = ~(U207 & P2_DATAO_REG_3__SCAN_IN); 
assign U400 = ~(U388 & BUF1_REG_3__SCAN_IN); 
assign U401 = ~(U207 & P2_DATAO_REG_4__SCAN_IN); 
assign U403 = ~(U388 & BUF1_REG_4__SCAN_IN); 
assign U404 = ~(U207 & P2_DATAO_REG_5__SCAN_IN); 
assign U406 = ~(U388 & BUF1_REG_5__SCAN_IN); 
assign U407 = ~(U207 & P2_DATAO_REG_6__SCAN_IN); 
assign U409 = ~(U388 & BUF1_REG_6__SCAN_IN); 
assign U410 = ~(U207 & P2_DATAO_REG_7__SCAN_IN); 
assign U412 = ~(U388 & BUF1_REG_7__SCAN_IN); 
assign U413 = ~(U207 & P2_DATAO_REG_8__SCAN_IN); 
assign U415 = ~(U388 & BUF1_REG_8__SCAN_IN); 
assign U416 = ~(U207 & P2_DATAO_REG_9__SCAN_IN); 
assign U418 = ~(U388 & BUF1_REG_9__SCAN_IN); 
assign U419 = ~(U207 & P2_DATAO_REG_10__SCAN_IN); 
assign U421 = ~(U388 & BUF1_REG_10__SCAN_IN); 
assign U422 = ~(U207 & P2_DATAO_REG_11__SCAN_IN); 
assign U424 = ~(U388 & BUF1_REG_11__SCAN_IN); 
assign U425 = ~(U207 & P2_DATAO_REG_12__SCAN_IN); 
assign U427 = ~(U388 & BUF1_REG_12__SCAN_IN); 
assign U428 = ~(U207 & P2_DATAO_REG_13__SCAN_IN); 
assign U430 = ~(U388 & BUF1_REG_13__SCAN_IN); 
assign U431 = ~(U207 & P2_DATAO_REG_14__SCAN_IN); 
assign U433 = ~(U388 & BUF1_REG_14__SCAN_IN); 
assign U434 = ~(U207 & P2_DATAO_REG_15__SCAN_IN); 
assign U436 = ~(U388 & BUF1_REG_15__SCAN_IN); 
assign U437 = ~(U207 & P2_DATAO_REG_16__SCAN_IN); 
assign U439 = ~(U388 & BUF1_REG_16__SCAN_IN); 
assign U440 = ~(U207 & P2_DATAO_REG_17__SCAN_IN); 
assign U442 = ~(U388 & BUF1_REG_17__SCAN_IN); 
assign U443 = ~(U207 & P2_DATAO_REG_18__SCAN_IN); 
assign U445 = ~(U388 & BUF1_REG_18__SCAN_IN); 
assign U446 = ~(U207 & P2_DATAO_REG_19__SCAN_IN); 
assign U448 = ~(U388 & BUF1_REG_19__SCAN_IN); 
assign U449 = ~(U207 & P2_DATAO_REG_20__SCAN_IN); 
assign U451 = ~(U388 & BUF1_REG_20__SCAN_IN); 
assign U452 = ~(U207 & P2_DATAO_REG_21__SCAN_IN); 
assign U454 = ~(U388 & BUF1_REG_21__SCAN_IN); 
assign U455 = ~(U207 & P2_DATAO_REG_22__SCAN_IN); 
assign U457 = ~(U388 & BUF1_REG_22__SCAN_IN); 
assign U458 = ~(U207 & P2_DATAO_REG_23__SCAN_IN); 
assign U460 = ~(U388 & BUF1_REG_23__SCAN_IN); 
assign U461 = ~(U207 & P2_DATAO_REG_24__SCAN_IN); 
assign U463 = ~(U388 & BUF1_REG_24__SCAN_IN); 
assign U464 = ~(U207 & P2_DATAO_REG_25__SCAN_IN); 
assign U466 = ~(U388 & BUF1_REG_25__SCAN_IN); 
assign U467 = ~(U207 & P2_DATAO_REG_26__SCAN_IN); 
assign U469 = ~(U388 & BUF1_REG_26__SCAN_IN); 
assign U470 = ~(U207 & P2_DATAO_REG_27__SCAN_IN); 
assign U472 = ~(U388 & BUF1_REG_27__SCAN_IN); 
assign U473 = ~(U207 & P2_DATAO_REG_28__SCAN_IN); 
assign U475 = ~(U388 & BUF1_REG_28__SCAN_IN); 
assign U476 = ~(U207 & P2_DATAO_REG_29__SCAN_IN); 
assign U478 = ~(U388 & BUF1_REG_29__SCAN_IN); 
assign U479 = ~(U207 & P2_DATAO_REG_30__SCAN_IN); 
assign U481 = ~(U388 & BUF1_REG_30__SCAN_IN); 
assign U482 = ~(U207 & P2_DATAO_REG_31__SCAN_IN); 
assign U484 = ~(U388 & BUF1_REG_31__SCAN_IN); 
assign P3_U2458 = P3_U4652 & P3_U3269; 
assign P3_U2460 = P3_U7962 & P3_U4652; 
assign P3_U2496 = P3_U4643 & P3_U3128; 
assign P3_U2521 = P3_U2520 & P3_U2519; 
assign P3_U2523 = P3_U2520 & P3_U2522; 
assign P3_U2525 = P3_U2520 & P3_U2524; 
assign P3_U2527 = P3_U2520 & P3_U2526; 
assign P3_U2529 = P3_U2528 & P3_U2519; 
assign P3_U2530 = P3_U2528 & P3_U2522; 
assign P3_U2531 = P3_U2528 & P3_U2524; 
assign P3_U2532 = P3_U2528 & P3_U2526; 
assign P3_U2554 = P3_U2553 & P3_U2468; 
assign P3_U2555 = P3_U2553 & P3_U4467; 
assign P3_U2556 = P3_U2553 & P3_U4332; 
assign P3_U2557 = P3_U2553 & P3_U2466; 
assign P3_U2559 = P3_U2558 & P3_U2468; 
assign P3_U2560 = P3_U2558 & P3_U4467; 
assign P3_U2561 = P3_U2558 & P3_U4332; 
assign P3_U2562 = P3_U2558 & P3_U2466; 
assign P3_U2564 = P3_U2563 & P3_U2522; 
assign P3_U2565 = P3_U2563 & P3_U2519; 
assign P3_U2566 = P3_U2563 & P3_U2526; 
assign P3_U2567 = P3_U2563 & P3_U2524; 
assign P3_U2569 = P3_U2568 & P3_U2522; 
assign P3_U2570 = P3_U2568 & P3_U2519; 
assign P3_U2571 = P3_U2568 & P3_U2526; 
assign P3_U2572 = P3_U2568 & P3_U2524; 
assign P3_U2636 = ~(P3_U8021 & P3_U8020 & P3_U4335); 
assign P3_U3029 = ~(P3_U7934 & P3_U7933 & P3_U4463); 
assign P3_U3031 = ~(P3_U3310 & P3_U4457); 
assign P3_U3070 = ~(P3_U2457 & P3_U4642); 
assign P3_U3071 = ~(P3_U2459 & P3_U4642); 
assign P3_U3074 = ~(P3_U3346 & P3_U3345 & P3_U3347 & P3_U3344 & P3_U3343); 
assign P3_U3101 = ~(P3_U3341 & P3_U3340 & P3_U3342 & P3_U3339 & P3_U3338); 
assign P3_U3102 = ~(P3_U3326 & P3_U3325 & P3_U3327 & P3_U3324 & P3_U3323); 
assign P3_U3104 = ~(P3_U3321 & P3_U3320 & P3_U3322 & P3_U3319 & P3_U3318); 
assign P3_U3107 = ~(P3_U3331 & P3_U3330 & P3_U3332 & P3_U3329 & P3_U3328); 
assign P3_U3108 = ~(P3_U3316 & P3_U3315 & P3_U3317 & P3_U3314 & P3_U3313); 
assign P3_U3110 = ~(P3_U3351 & P3_U3350 & P3_U3352 & P3_U3349 & P3_U3348); 
assign P3_U3155 = ~(P3_U4643 & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P3_U3218 = ~(P3_U3336 & P3_U3335 & P3_U3337 & P3_U3334 & P3_U3333); 
assign P3_U3280 = ~(P3_U7939 & P3_U7938); 
assign P3_U3281 = ~(P3_U7941 & P3_U7940); 
assign P3_U3301 = ~(P3_U8041 & P3_U8040); 
assign P3_U3683 = P3_U5568 & P3_U5567; 
assign P3_U4250 = P3_U7787 & P3_U7786 & P3_U7785 & P3_U7784; 
assign P3_U4254 = P3_U7803 & P3_U7802 & P3_U7801 & P3_U7800; 
assign P3_U4258 = P3_U7819 & P3_U7818 & P3_U7817 & P3_U7816; 
assign P3_U4262 = P3_U7835 & P3_U7834 & P3_U7833 & P3_U7832; 
assign P3_U4266 = P3_U7851 & P3_U7850 & P3_U7849 & P3_U7848; 
assign P3_U4270 = P3_U7867 & P3_U7866 & P3_U7865 & P3_U7864; 
assign P3_U4274 = P3_U7883 & P3_U7882 & P3_U7881 & P3_U7880; 
assign P3_U4278 = P3_U7899 & P3_U7898 & P3_U7897 & P3_U7896; 
assign P3_U4644 = ~P3_U3148; 
assign P3_U4657 = ~P3_U3140; 
assign P3_U4663 = ~(P3_U2457 & P3_U4653); 
assign P3_U4717 = ~(P3_U4342 & P3_U2457); 
assign P3_U4769 = ~(P3_U4343 & P3_U2457); 
assign P3_U4872 = ~(P3_U2459 & P3_U4653); 
assign P3_U4924 = ~(P3_U2459 & P3_U4342); 
assign P3_U4976 = ~(P3_U2459 & P3_U4343); 
assign P3_U5594 = ~(P3_U3270 & P3_U5582); 
assign P3_U7387 = ~(P3_U2542 & P3_INSTQUEUE_REG_15__7__SCAN_IN); 
assign P3_U7388 = ~(P3_U2541 & P3_INSTQUEUE_REG_14__7__SCAN_IN); 
assign P3_U7389 = ~(P3_U2540 & P3_INSTQUEUE_REG_13__7__SCAN_IN); 
assign P3_U7390 = ~(P3_U2539 & P3_INSTQUEUE_REG_12__7__SCAN_IN); 
assign P3_U7391 = ~(P3_U2537 & P3_INSTQUEUE_REG_11__7__SCAN_IN); 
assign P3_U7392 = ~(P3_U2536 & P3_INSTQUEUE_REG_10__7__SCAN_IN); 
assign P3_U7393 = ~(P3_U2535 & P3_INSTQUEUE_REG_9__7__SCAN_IN); 
assign P3_U7394 = ~(P3_U2534 & P3_INSTQUEUE_REG_8__7__SCAN_IN); 
assign P3_U7403 = ~(P3_U2542 & P3_INSTQUEUE_REG_15__6__SCAN_IN); 
assign P3_U7404 = ~(P3_U2541 & P3_INSTQUEUE_REG_14__6__SCAN_IN); 
assign P3_U7405 = ~(P3_U2540 & P3_INSTQUEUE_REG_13__6__SCAN_IN); 
assign P3_U7406 = ~(P3_U2539 & P3_INSTQUEUE_REG_12__6__SCAN_IN); 
assign P3_U7407 = ~(P3_U2537 & P3_INSTQUEUE_REG_11__6__SCAN_IN); 
assign P3_U7408 = ~(P3_U2536 & P3_INSTQUEUE_REG_10__6__SCAN_IN); 
assign P3_U7409 = ~(P3_U2535 & P3_INSTQUEUE_REG_9__6__SCAN_IN); 
assign P3_U7410 = ~(P3_U2534 & P3_INSTQUEUE_REG_8__6__SCAN_IN); 
assign P3_U7419 = ~(P3_U2542 & P3_INSTQUEUE_REG_15__5__SCAN_IN); 
assign P3_U7420 = ~(P3_U2541 & P3_INSTQUEUE_REG_14__5__SCAN_IN); 
assign P3_U7421 = ~(P3_U2540 & P3_INSTQUEUE_REG_13__5__SCAN_IN); 
assign P3_U7422 = ~(P3_U2539 & P3_INSTQUEUE_REG_12__5__SCAN_IN); 
assign P3_U7423 = ~(P3_U2537 & P3_INSTQUEUE_REG_11__5__SCAN_IN); 
assign P3_U7424 = ~(P3_U2536 & P3_INSTQUEUE_REG_10__5__SCAN_IN); 
assign P3_U7425 = ~(P3_U2535 & P3_INSTQUEUE_REG_9__5__SCAN_IN); 
assign P3_U7426 = ~(P3_U2534 & P3_INSTQUEUE_REG_8__5__SCAN_IN); 
assign P3_U7435 = ~(P3_U2542 & P3_INSTQUEUE_REG_15__4__SCAN_IN); 
assign P3_U7436 = ~(P3_U2541 & P3_INSTQUEUE_REG_14__4__SCAN_IN); 
assign P3_U7437 = ~(P3_U2540 & P3_INSTQUEUE_REG_13__4__SCAN_IN); 
assign P3_U7438 = ~(P3_U2539 & P3_INSTQUEUE_REG_12__4__SCAN_IN); 
assign P3_U7439 = ~(P3_U2537 & P3_INSTQUEUE_REG_11__4__SCAN_IN); 
assign P3_U7440 = ~(P3_U2536 & P3_INSTQUEUE_REG_10__4__SCAN_IN); 
assign P3_U7441 = ~(P3_U2535 & P3_INSTQUEUE_REG_9__4__SCAN_IN); 
assign P3_U7442 = ~(P3_U2534 & P3_INSTQUEUE_REG_8__4__SCAN_IN); 
assign P3_U7451 = ~(P3_U2542 & P3_INSTQUEUE_REG_15__3__SCAN_IN); 
assign P3_U7452 = ~(P3_U2541 & P3_INSTQUEUE_REG_14__3__SCAN_IN); 
assign P3_U7453 = ~(P3_U2540 & P3_INSTQUEUE_REG_13__3__SCAN_IN); 
assign P3_U7454 = ~(P3_U2539 & P3_INSTQUEUE_REG_12__3__SCAN_IN); 
assign P3_U7455 = ~(P3_U2537 & P3_INSTQUEUE_REG_11__3__SCAN_IN); 
assign P3_U7456 = ~(P3_U2536 & P3_INSTQUEUE_REG_10__3__SCAN_IN); 
assign P3_U7457 = ~(P3_U2535 & P3_INSTQUEUE_REG_9__3__SCAN_IN); 
assign P3_U7458 = ~(P3_U2534 & P3_INSTQUEUE_REG_8__3__SCAN_IN); 
assign P3_U7467 = ~(P3_U2542 & P3_INSTQUEUE_REG_15__2__SCAN_IN); 
assign P3_U7468 = ~(P3_U2541 & P3_INSTQUEUE_REG_14__2__SCAN_IN); 
assign P3_U7469 = ~(P3_U2540 & P3_INSTQUEUE_REG_13__2__SCAN_IN); 
assign P3_U7470 = ~(P3_U2539 & P3_INSTQUEUE_REG_12__2__SCAN_IN); 
assign P3_U7471 = ~(P3_U2537 & P3_INSTQUEUE_REG_11__2__SCAN_IN); 
assign P3_U7472 = ~(P3_U2536 & P3_INSTQUEUE_REG_10__2__SCAN_IN); 
assign P3_U7473 = ~(P3_U2535 & P3_INSTQUEUE_REG_9__2__SCAN_IN); 
assign P3_U7474 = ~(P3_U2534 & P3_INSTQUEUE_REG_8__2__SCAN_IN); 
assign P3_U7483 = ~(P3_U2542 & P3_INSTQUEUE_REG_15__1__SCAN_IN); 
assign P3_U7484 = ~(P3_U2541 & P3_INSTQUEUE_REG_14__1__SCAN_IN); 
assign P3_U7485 = ~(P3_U2540 & P3_INSTQUEUE_REG_13__1__SCAN_IN); 
assign P3_U7486 = ~(P3_U2539 & P3_INSTQUEUE_REG_12__1__SCAN_IN); 
assign P3_U7487 = ~(P3_U2537 & P3_INSTQUEUE_REG_11__1__SCAN_IN); 
assign P3_U7488 = ~(P3_U2536 & P3_INSTQUEUE_REG_10__1__SCAN_IN); 
assign P3_U7489 = ~(P3_U2535 & P3_INSTQUEUE_REG_9__1__SCAN_IN); 
assign P3_U7490 = ~(P3_U2534 & P3_INSTQUEUE_REG_8__1__SCAN_IN); 
assign P3_U7499 = ~(P3_U2542 & P3_INSTQUEUE_REG_15__0__SCAN_IN); 
assign P3_U7500 = ~(P3_U2541 & P3_INSTQUEUE_REG_14__0__SCAN_IN); 
assign P3_U7501 = ~(P3_U2540 & P3_INSTQUEUE_REG_13__0__SCAN_IN); 
assign P3_U7502 = ~(P3_U2539 & P3_INSTQUEUE_REG_12__0__SCAN_IN); 
assign P3_U7503 = ~(P3_U2537 & P3_INSTQUEUE_REG_11__0__SCAN_IN); 
assign P3_U7504 = ~(P3_U2536 & P3_INSTQUEUE_REG_10__0__SCAN_IN); 
assign P3_U7505 = ~(P3_U2535 & P3_INSTQUEUE_REG_9__0__SCAN_IN); 
assign P3_U7506 = ~(P3_U2534 & P3_INSTQUEUE_REG_8__0__SCAN_IN); 
assign P3_U7525 = ~(P3_U2552 & P3_INSTQUEUE_REG_8__7__SCAN_IN); 
assign P3_U7526 = ~(P3_U2551 & P3_INSTQUEUE_REG_9__7__SCAN_IN); 
assign P3_U7527 = ~(P3_U2550 & P3_INSTQUEUE_REG_10__7__SCAN_IN); 
assign P3_U7528 = ~(P3_U2549 & P3_INSTQUEUE_REG_11__7__SCAN_IN); 
assign P3_U7529 = ~(P3_U2547 & P3_INSTQUEUE_REG_12__7__SCAN_IN); 
assign P3_U7530 = ~(P3_U2546 & P3_INSTQUEUE_REG_13__7__SCAN_IN); 
assign P3_U7531 = ~(P3_U2545 & P3_INSTQUEUE_REG_14__7__SCAN_IN); 
assign P3_U7532 = ~(P3_U2544 & P3_INSTQUEUE_REG_15__7__SCAN_IN); 
assign P3_U7541 = ~(P3_U2552 & P3_INSTQUEUE_REG_8__6__SCAN_IN); 
assign P3_U7542 = ~(P3_U2551 & P3_INSTQUEUE_REG_9__6__SCAN_IN); 
assign P3_U7543 = ~(P3_U2550 & P3_INSTQUEUE_REG_10__6__SCAN_IN); 
assign P3_U7544 = ~(P3_U2549 & P3_INSTQUEUE_REG_11__6__SCAN_IN); 
assign P3_U7545 = ~(P3_U2547 & P3_INSTQUEUE_REG_12__6__SCAN_IN); 
assign P3_U7546 = ~(P3_U2546 & P3_INSTQUEUE_REG_13__6__SCAN_IN); 
assign P3_U7547 = ~(P3_U2545 & P3_INSTQUEUE_REG_14__6__SCAN_IN); 
assign P3_U7548 = ~(P3_U2544 & P3_INSTQUEUE_REG_15__6__SCAN_IN); 
assign P3_U7557 = ~(P3_U2552 & P3_INSTQUEUE_REG_8__5__SCAN_IN); 
assign P3_U7558 = ~(P3_U2551 & P3_INSTQUEUE_REG_9__5__SCAN_IN); 
assign P3_U7559 = ~(P3_U2550 & P3_INSTQUEUE_REG_10__5__SCAN_IN); 
assign P3_U7560 = ~(P3_U2549 & P3_INSTQUEUE_REG_11__5__SCAN_IN); 
assign P3_U7561 = ~(P3_U2547 & P3_INSTQUEUE_REG_12__5__SCAN_IN); 
assign P3_U7562 = ~(P3_U2546 & P3_INSTQUEUE_REG_13__5__SCAN_IN); 
assign P3_U7563 = ~(P3_U2545 & P3_INSTQUEUE_REG_14__5__SCAN_IN); 
assign P3_U7564 = ~(P3_U2544 & P3_INSTQUEUE_REG_15__5__SCAN_IN); 
assign P3_U7573 = ~(P3_U2552 & P3_INSTQUEUE_REG_8__4__SCAN_IN); 
assign P3_U7574 = ~(P3_U2551 & P3_INSTQUEUE_REG_9__4__SCAN_IN); 
assign P3_U7575 = ~(P3_U2550 & P3_INSTQUEUE_REG_10__4__SCAN_IN); 
assign P3_U7576 = ~(P3_U2549 & P3_INSTQUEUE_REG_11__4__SCAN_IN); 
assign P3_U7577 = ~(P3_U2547 & P3_INSTQUEUE_REG_12__4__SCAN_IN); 
assign P3_U7578 = ~(P3_U2546 & P3_INSTQUEUE_REG_13__4__SCAN_IN); 
assign P3_U7579 = ~(P3_U2545 & P3_INSTQUEUE_REG_14__4__SCAN_IN); 
assign P3_U7580 = ~(P3_U2544 & P3_INSTQUEUE_REG_15__4__SCAN_IN); 
assign P3_U7589 = ~(P3_U2552 & P3_INSTQUEUE_REG_8__3__SCAN_IN); 
assign P3_U7590 = ~(P3_U2551 & P3_INSTQUEUE_REG_9__3__SCAN_IN); 
assign P3_U7591 = ~(P3_U2550 & P3_INSTQUEUE_REG_10__3__SCAN_IN); 
assign P3_U7592 = ~(P3_U2549 & P3_INSTQUEUE_REG_11__3__SCAN_IN); 
assign P3_U7593 = ~(P3_U2547 & P3_INSTQUEUE_REG_12__3__SCAN_IN); 
assign P3_U7594 = ~(P3_U2546 & P3_INSTQUEUE_REG_13__3__SCAN_IN); 
assign P3_U7595 = ~(P3_U2545 & P3_INSTQUEUE_REG_14__3__SCAN_IN); 
assign P3_U7596 = ~(P3_U2544 & P3_INSTQUEUE_REG_15__3__SCAN_IN); 
assign P3_U7605 = ~(P3_U2552 & P3_INSTQUEUE_REG_8__2__SCAN_IN); 
assign P3_U7606 = ~(P3_U2551 & P3_INSTQUEUE_REG_9__2__SCAN_IN); 
assign P3_U7607 = ~(P3_U2550 & P3_INSTQUEUE_REG_10__2__SCAN_IN); 
assign P3_U7608 = ~(P3_U2549 & P3_INSTQUEUE_REG_11__2__SCAN_IN); 
assign P3_U7609 = ~(P3_U2547 & P3_INSTQUEUE_REG_12__2__SCAN_IN); 
assign P3_U7610 = ~(P3_U2546 & P3_INSTQUEUE_REG_13__2__SCAN_IN); 
assign P3_U7611 = ~(P3_U2545 & P3_INSTQUEUE_REG_14__2__SCAN_IN); 
assign P3_U7612 = ~(P3_U2544 & P3_INSTQUEUE_REG_15__2__SCAN_IN); 
assign P3_U7621 = ~(P3_U2552 & P3_INSTQUEUE_REG_8__1__SCAN_IN); 
assign P3_U7622 = ~(P3_U2551 & P3_INSTQUEUE_REG_9__1__SCAN_IN); 
assign P3_U7623 = ~(P3_U2550 & P3_INSTQUEUE_REG_10__1__SCAN_IN); 
assign P3_U7624 = ~(P3_U2549 & P3_INSTQUEUE_REG_11__1__SCAN_IN); 
assign P3_U7625 = ~(P3_U2547 & P3_INSTQUEUE_REG_12__1__SCAN_IN); 
assign P3_U7626 = ~(P3_U2546 & P3_INSTQUEUE_REG_13__1__SCAN_IN); 
assign P3_U7627 = ~(P3_U2545 & P3_INSTQUEUE_REG_14__1__SCAN_IN); 
assign P3_U7628 = ~(P3_U2544 & P3_INSTQUEUE_REG_15__1__SCAN_IN); 
assign P3_U7637 = ~(P3_U2552 & P3_INSTQUEUE_REG_8__0__SCAN_IN); 
assign P3_U7638 = ~(P3_U2551 & P3_INSTQUEUE_REG_9__0__SCAN_IN); 
assign P3_U7639 = ~(P3_U2550 & P3_INSTQUEUE_REG_10__0__SCAN_IN); 
assign P3_U7640 = ~(P3_U2549 & P3_INSTQUEUE_REG_11__0__SCAN_IN); 
assign P3_U7641 = ~(P3_U2547 & P3_INSTQUEUE_REG_12__0__SCAN_IN); 
assign P3_U7642 = ~(P3_U2546 & P3_INSTQUEUE_REG_13__0__SCAN_IN); 
assign P3_U7643 = ~(P3_U2545 & P3_INSTQUEUE_REG_14__0__SCAN_IN); 
assign P3_U7644 = ~(P3_U2544 & P3_INSTQUEUE_REG_15__0__SCAN_IN); 
assign P3_U7646 = ~(P3_U2582 & P3_INSTQUEUE_REG_8__7__SCAN_IN); 
assign P3_U7647 = ~(P3_U2581 & P3_INSTQUEUE_REG_9__7__SCAN_IN); 
assign P3_U7648 = ~(P3_U2580 & P3_INSTQUEUE_REG_10__7__SCAN_IN); 
assign P3_U7649 = ~(P3_U2579 & P3_INSTQUEUE_REG_11__7__SCAN_IN); 
assign P3_U7650 = ~(P3_U2577 & P3_INSTQUEUE_REG_12__7__SCAN_IN); 
assign P3_U7651 = ~(P3_U2576 & P3_INSTQUEUE_REG_13__7__SCAN_IN); 
assign P3_U7652 = ~(P3_U2575 & P3_INSTQUEUE_REG_14__7__SCAN_IN); 
assign P3_U7653 = ~(P3_U2574 & P3_INSTQUEUE_REG_15__7__SCAN_IN); 
assign P3_U7662 = ~(P3_U2582 & P3_INSTQUEUE_REG_8__6__SCAN_IN); 
assign P3_U7663 = ~(P3_U2581 & P3_INSTQUEUE_REG_9__6__SCAN_IN); 
assign P3_U7664 = ~(P3_U2580 & P3_INSTQUEUE_REG_10__6__SCAN_IN); 
assign P3_U7665 = ~(P3_U2579 & P3_INSTQUEUE_REG_11__6__SCAN_IN); 
assign P3_U7666 = ~(P3_U2577 & P3_INSTQUEUE_REG_12__6__SCAN_IN); 
assign P3_U7667 = ~(P3_U2576 & P3_INSTQUEUE_REG_13__6__SCAN_IN); 
assign P3_U7668 = ~(P3_U2575 & P3_INSTQUEUE_REG_14__6__SCAN_IN); 
assign P3_U7669 = ~(P3_U2574 & P3_INSTQUEUE_REG_15__6__SCAN_IN); 
assign P3_U7678 = ~(P3_U2582 & P3_INSTQUEUE_REG_8__5__SCAN_IN); 
assign P3_U7679 = ~(P3_U2581 & P3_INSTQUEUE_REG_9__5__SCAN_IN); 
assign P3_U7680 = ~(P3_U2580 & P3_INSTQUEUE_REG_10__5__SCAN_IN); 
assign P3_U7681 = ~(P3_U2579 & P3_INSTQUEUE_REG_11__5__SCAN_IN); 
assign P3_U7682 = ~(P3_U2577 & P3_INSTQUEUE_REG_12__5__SCAN_IN); 
assign P3_U7683 = ~(P3_U2576 & P3_INSTQUEUE_REG_13__5__SCAN_IN); 
assign P3_U7684 = ~(P3_U2575 & P3_INSTQUEUE_REG_14__5__SCAN_IN); 
assign P3_U7685 = ~(P3_U2574 & P3_INSTQUEUE_REG_15__5__SCAN_IN); 
assign P3_U7694 = ~(P3_U2582 & P3_INSTQUEUE_REG_8__4__SCAN_IN); 
assign P3_U7695 = ~(P3_U2581 & P3_INSTQUEUE_REG_9__4__SCAN_IN); 
assign P3_U7696 = ~(P3_U2580 & P3_INSTQUEUE_REG_10__4__SCAN_IN); 
assign P3_U7697 = ~(P3_U2579 & P3_INSTQUEUE_REG_11__4__SCAN_IN); 
assign P3_U7698 = ~(P3_U2577 & P3_INSTQUEUE_REG_12__4__SCAN_IN); 
assign P3_U7699 = ~(P3_U2576 & P3_INSTQUEUE_REG_13__4__SCAN_IN); 
assign P3_U7700 = ~(P3_U2575 & P3_INSTQUEUE_REG_14__4__SCAN_IN); 
assign P3_U7701 = ~(P3_U2574 & P3_INSTQUEUE_REG_15__4__SCAN_IN); 
assign P3_U7710 = ~(P3_U2582 & P3_INSTQUEUE_REG_8__3__SCAN_IN); 
assign P3_U7711 = ~(P3_U2581 & P3_INSTQUEUE_REG_9__3__SCAN_IN); 
assign P3_U7712 = ~(P3_U2580 & P3_INSTQUEUE_REG_10__3__SCAN_IN); 
assign P3_U7713 = ~(P3_U2579 & P3_INSTQUEUE_REG_11__3__SCAN_IN); 
assign P3_U7714 = ~(P3_U2577 & P3_INSTQUEUE_REG_12__3__SCAN_IN); 
assign P3_U7715 = ~(P3_U2576 & P3_INSTQUEUE_REG_13__3__SCAN_IN); 
assign P3_U7716 = ~(P3_U2575 & P3_INSTQUEUE_REG_14__3__SCAN_IN); 
assign P3_U7717 = ~(P3_U2574 & P3_INSTQUEUE_REG_15__3__SCAN_IN); 
assign P3_U7726 = ~(P3_U2582 & P3_INSTQUEUE_REG_8__2__SCAN_IN); 
assign P3_U7727 = ~(P3_U2581 & P3_INSTQUEUE_REG_9__2__SCAN_IN); 
assign P3_U7728 = ~(P3_U2580 & P3_INSTQUEUE_REG_10__2__SCAN_IN); 
assign P3_U7729 = ~(P3_U2579 & P3_INSTQUEUE_REG_11__2__SCAN_IN); 
assign P3_U7730 = ~(P3_U2577 & P3_INSTQUEUE_REG_12__2__SCAN_IN); 
assign P3_U7731 = ~(P3_U2576 & P3_INSTQUEUE_REG_13__2__SCAN_IN); 
assign P3_U7732 = ~(P3_U2575 & P3_INSTQUEUE_REG_14__2__SCAN_IN); 
assign P3_U7733 = ~(P3_U2574 & P3_INSTQUEUE_REG_15__2__SCAN_IN); 
assign P3_U7742 = ~(P3_U2582 & P3_INSTQUEUE_REG_8__1__SCAN_IN); 
assign P3_U7743 = ~(P3_U2581 & P3_INSTQUEUE_REG_9__1__SCAN_IN); 
assign P3_U7744 = ~(P3_U2580 & P3_INSTQUEUE_REG_10__1__SCAN_IN); 
assign P3_U7745 = ~(P3_U2579 & P3_INSTQUEUE_REG_11__1__SCAN_IN); 
assign P3_U7746 = ~(P3_U2577 & P3_INSTQUEUE_REG_12__1__SCAN_IN); 
assign P3_U7747 = ~(P3_U2576 & P3_INSTQUEUE_REG_13__1__SCAN_IN); 
assign P3_U7748 = ~(P3_U2575 & P3_INSTQUEUE_REG_14__1__SCAN_IN); 
assign P3_U7749 = ~(P3_U2574 & P3_INSTQUEUE_REG_15__1__SCAN_IN); 
assign P3_U7758 = ~(P3_U2582 & P3_INSTQUEUE_REG_8__0__SCAN_IN); 
assign P3_U7759 = ~(P3_U2581 & P3_INSTQUEUE_REG_9__0__SCAN_IN); 
assign P3_U7760 = ~(P3_U2580 & P3_INSTQUEUE_REG_10__0__SCAN_IN); 
assign P3_U7761 = ~(P3_U2579 & P3_INSTQUEUE_REG_11__0__SCAN_IN); 
assign P3_U7762 = ~(P3_U2577 & P3_INSTQUEUE_REG_12__0__SCAN_IN); 
assign P3_U7763 = ~(P3_U2576 & P3_INSTQUEUE_REG_13__0__SCAN_IN); 
assign P3_U7764 = ~(P3_U2575 & P3_INSTQUEUE_REG_14__0__SCAN_IN); 
assign P3_U7765 = ~(P3_U2574 & P3_INSTQUEUE_REG_15__0__SCAN_IN); 
assign P3_U7965 = ~P3_U3270; 
assign P3_U7967 = ~(P3_U3270 & P3_U3140); 
assign P2_U2352 = P2_U2617 & P2_U3300 & P2_U7873; 
assign P2_U2354 = P2_U7861 & P2_U7873 & P2_STATE2_REG_0__SCAN_IN; 
assign P2_U2355 = P2_U2447 & P2_U7861; 
assign P2_U2436 = P2_U7859 & P2_U7867; 
assign P2_U2438 = P2_U7859 & P2_U3278; 
assign P2_U2458 = P2_U2617 & P2_U3279 & P2_U7863; 
assign P2_U2578 = P2_U2577 & P2_U2563; 
assign P2_U2579 = P2_U2577 & P2_U2566; 
assign P2_U2580 = P2_U2577 & P2_U2568; 
assign P2_U2581 = P2_U2577 & P2_U2570; 
assign P2_U2583 = P2_U2563 & P2_U2582; 
assign P2_U2584 = P2_U2566 & P2_U2582; 
assign P2_U2585 = P2_U2568 & P2_U2582; 
assign P2_U2586 = P2_U2570 & P2_U2582; 
assign P2_U2591 = ~(P2_U4274 & P2_U4273); 
assign P2_U2592 = ~(P2_U4272 & P2_U4271); 
assign P2_U2593 = ~(P2_U4270 & P2_U4269); 
assign P2_U2594 = ~(P2_U4268 & P2_U4267); 
assign P2_U2595 = ~(P2_U4266 & P2_U4265); 
assign P2_U2596 = ~(P2_U4264 & P2_U4263); 
assign P2_U2597 = ~(P2_U4262 & P2_U4261); 
assign P2_U2598 = ~(P2_U4260 & P2_U4259); 
assign P2_U2715 = ~(P2_U2356 & P2_U2616); 
assign P2_U2752 = P2_U3280 & P2_U7873 & P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P2_U2818 = ~(P2_U8136 & P2_U8135 & P2_U4463); 
assign P2_U2822 = ~(P2_U4398 & P2_U6836); 
assign P2_U3209 = ~(P2_U7914 & P2_U7913 & P2_U4588); 
assign P2_U3211 = ~(P2_U3690 & P2_U4579); 
assign P2_U3281 = ~(P2_U7861 & P2_U7863 & P2_U7859); 
assign P2_U3283 = ~(P2_U3253 & P2_U7873); 
assign P2_U3289 = ~(P2_U2616 & P2_U7871); 
assign P2_U3294 = ~(P2_U7871 & P2_U7873); 
assign P2_U3295 = ~(P2_U7861 & P2_U2617); 
assign P2_U3380 = ~(P2_U3377 & P2_U4885); 
assign P2_U3403 = ~(P2_U3401 & P2_U5000); 
assign P2_U3429 = ~(P2_U3424 & P2_U5114); 
assign P2_U3452 = ~(P2_U3450 & P2_U5228); 
assign P2_U3475 = ~(P2_U3473 & P2_U5343); 
assign P2_U3498 = ~(P2_U3496 & P2_U5458); 
assign P2_U3525 = ~(P2_U7865 & P2_U7863 & P2_U3279 & P2_U7869); 
assign P2_U3536 = ~(P2_U7873 & P2_STATE2_REG_0__SCAN_IN); 
assign P2_U3571 = ~(P2_U7865 & P2_U3300); 
assign P2_U3591 = ~(P2_U7919 & P2_U7918); 
assign P2_U3592 = ~(P2_U7921 & P2_U7920); 
assign P2_U3657 = ~(P2_U8370 & P2_U8369); 
assign P2_U3712 = P2_U3521 & P2_U7867; 
assign P2_U3873 = P2_U3521 & P2_U7869; 
assign P2_U3874 = P2_U7861 & P2_U3278; 
assign P2_U3878 = P2_U7863 & P2_U3521; 
assign P2_U3887 = P2_U3582 & P2_U7859; 
assign P2_U3889 = P2_U7859 & P2_U3272; 
assign P2_U4055 = P2_U4468 & P2_U6133 & P2_U2356; 
assign P2_U4056 = P2_U3280 & P2_U7871 & P2_STATE2_REG_0__SCAN_IN; 
assign P2_U4184 = P2_U6844 & P2_U7873; 
assign P2_U4191 = P2_U6865 & P2_U6864 & P2_U6863 & P2_U6862; 
assign P2_U4192 = P2_U6869 & P2_U6868 & P2_U6867 & P2_U6866; 
assign P2_U4195 = P2_U6881 & P2_U6880 & P2_U6879 & P2_U6878; 
assign P2_U4196 = P2_U6885 & P2_U6884 & P2_U6883 & P2_U6882; 
assign P2_U4199 = P2_U6897 & P2_U6896 & P2_U6895 & P2_U6894; 
assign P2_U4200 = P2_U6901 & P2_U6900 & P2_U6899 & P2_U6898; 
assign P2_U4203 = P2_U6913 & P2_U6912 & P2_U6911 & P2_U6910; 
assign P2_U4204 = P2_U6917 & P2_U6916 & P2_U6915 & P2_U6914; 
assign P2_U4207 = P2_U6929 & P2_U6928 & P2_U6927 & P2_U6926; 
assign P2_U4208 = P2_U6933 & P2_U6932 & P2_U6931 & P2_U6930; 
assign P2_U4211 = P2_U6945 & P2_U6944 & P2_U6943 & P2_U6942; 
assign P2_U4212 = P2_U6949 & P2_U6948 & P2_U6947 & P2_U6946; 
assign P2_U4215 = P2_U6961 & P2_U6960 & P2_U6959 & P2_U6958; 
assign P2_U4216 = P2_U6965 & P2_U6964 & P2_U6963 & P2_U6962; 
assign P2_U4219 = P2_U6977 & P2_U6976 & P2_U6975 & P2_U6974; 
assign P2_U4220 = P2_U6981 & P2_U6980 & P2_U6979 & P2_U6978; 
assign P2_U4223 = P2_U6993 & P2_U6992 & P2_U6991 & P2_U6990; 
assign P2_U4224 = P2_U6997 & P2_U6996 & P2_U6995 & P2_U6994; 
assign P2_U4275 = P2_U7861 & P2_U4276; 
assign P2_U4285 = P2_U7204 & P2_U7203 & P2_U7202 & P2_U7201; 
assign P2_U4286 = P2_U7208 & P2_U7207 & P2_U7206 & P2_U7205; 
assign P2_U4293 = P2_U7238 & P2_U7237 & P2_U7236 & P2_U7235; 
assign P2_U4294 = P2_U7242 & P2_U7241 & P2_U7240 & P2_U7239; 
assign P2_U4301 = P2_U7272 & P2_U7271 & P2_U7270 & P2_U7269; 
assign P2_U4302 = P2_U7276 & P2_U7275 & P2_U7274 & P2_U7273; 
assign P2_U4309 = P2_U7306 & P2_U7305 & P2_U7304 & P2_U7303; 
assign P2_U4310 = P2_U7310 & P2_U7309 & P2_U7308 & P2_U7307; 
assign P2_U4317 = P2_U7340 & P2_U7339 & P2_U7338 & P2_U7337; 
assign P2_U4318 = P2_U7344 & P2_U7343 & P2_U7342 & P2_U7341; 
assign P2_U4325 = P2_U7374 & P2_U7373 & P2_U7372 & P2_U7371; 
assign P2_U4326 = P2_U7378 & P2_U7377 & P2_U7376 & P2_U7375; 
assign P2_U4333 = P2_U7408 & P2_U7407 & P2_U7406 & P2_U7405; 
assign P2_U4334 = P2_U7412 & P2_U7411 & P2_U7410 & P2_U7409; 
assign P2_U4343 = P2_U7869 & P2_U7873; 
assign P2_U4377 = P2_U7863 & P2_U3255; 
assign P2_U4378 = P2_U2356 & P2_U7873; 
assign P2_U4381 = P2_U2356 & P2_U4595; 
assign P2_U4414 = ~(P2_U2616 & P2_U3300 & P2_U7869); 
assign P2_U4415 = ~(P2_U2447 & P2_U3279); 
assign P2_U4428 = ~P2_U3286; 
assign P2_U4457 = ~(P2_U2356 & P2_U3280); 
assign P2_U4652 = ~P2_U3325; 
assign P2_U4771 = ~P2_U3355; 
assign P2_U4943 = ~P2_U3247; 
assign P2_U5058 = ~P2_U3248; 
assign P2_U5171 = ~P2_U3249; 
assign P2_U5286 = ~P2_U3250; 
assign P2_U5401 = ~P2_U3251; 
assign P2_U5516 = ~P2_U3252; 
assign P2_U5571 = ~(P2_U3279 & P2_U7869); 
assign P2_U5573 = ~(P2_U7863 & P2_U2617 & P2_U7861); 
assign P2_U5588 = ~(P2_U7865 & P2_U3278); 
assign P2_U5597 = ~(P2_U3279 & P2_U7871); 
assign P2_U6870 = ~(P2_U2528 & P2_INSTQUEUE_REG_7__7__SCAN_IN); 
assign P2_U6871 = ~(P2_U2527 & P2_INSTQUEUE_REG_6__7__SCAN_IN); 
assign P2_U6872 = ~(P2_U2526 & P2_INSTQUEUE_REG_5__7__SCAN_IN); 
assign P2_U6873 = ~(P2_U2524 & P2_INSTQUEUE_REG_4__7__SCAN_IN); 
assign P2_U6874 = ~(P2_U2522 & P2_INSTQUEUE_REG_3__7__SCAN_IN); 
assign P2_U6875 = ~(P2_U2521 & P2_INSTQUEUE_REG_2__7__SCAN_IN); 
assign P2_U6876 = ~(P2_U2519 & P2_INSTQUEUE_REG_1__7__SCAN_IN); 
assign P2_U6877 = ~(P2_U2517 & P2_INSTQUEUE_REG_0__7__SCAN_IN); 
assign P2_U6886 = ~(P2_U2552 & P2_INSTQUEUE_REG_7__7__SCAN_IN); 
assign P2_U6887 = ~(P2_U2551 & P2_INSTQUEUE_REG_6__7__SCAN_IN); 
assign P2_U6890 = ~(P2_U2546 & P2_INSTQUEUE_REG_3__7__SCAN_IN); 
assign P2_U6891 = ~(P2_U2545 & P2_INSTQUEUE_REG_2__7__SCAN_IN); 
assign P2_U6902 = ~(P2_U2552 & P2_INSTQUEUE_REG_7__6__SCAN_IN); 
assign P2_U6903 = ~(P2_U2551 & P2_INSTQUEUE_REG_6__6__SCAN_IN); 
assign P2_U6906 = ~(P2_U2546 & P2_INSTQUEUE_REG_3__6__SCAN_IN); 
assign P2_U6907 = ~(P2_U2545 & P2_INSTQUEUE_REG_2__6__SCAN_IN); 
assign P2_U6918 = ~(P2_U2552 & P2_INSTQUEUE_REG_7__5__SCAN_IN); 
assign P2_U6919 = ~(P2_U2551 & P2_INSTQUEUE_REG_6__5__SCAN_IN); 
assign P2_U6922 = ~(P2_U2546 & P2_INSTQUEUE_REG_3__5__SCAN_IN); 
assign P2_U6923 = ~(P2_U2545 & P2_INSTQUEUE_REG_2__5__SCAN_IN); 
assign P2_U6934 = ~(P2_U2552 & P2_INSTQUEUE_REG_7__4__SCAN_IN); 
assign P2_U6935 = ~(P2_U2551 & P2_INSTQUEUE_REG_6__4__SCAN_IN); 
assign P2_U6938 = ~(P2_U2546 & P2_INSTQUEUE_REG_3__4__SCAN_IN); 
assign P2_U6939 = ~(P2_U2545 & P2_INSTQUEUE_REG_2__4__SCAN_IN); 
assign P2_U6950 = ~(P2_U2552 & P2_INSTQUEUE_REG_7__3__SCAN_IN); 
assign P2_U6951 = ~(P2_U2551 & P2_INSTQUEUE_REG_6__3__SCAN_IN); 
assign P2_U6954 = ~(P2_U2546 & P2_INSTQUEUE_REG_3__3__SCAN_IN); 
assign P2_U6955 = ~(P2_U2545 & P2_INSTQUEUE_REG_2__3__SCAN_IN); 
assign P2_U6966 = ~(P2_U2552 & P2_INSTQUEUE_REG_7__2__SCAN_IN); 
assign P2_U6967 = ~(P2_U2551 & P2_INSTQUEUE_REG_6__2__SCAN_IN); 
assign P2_U6970 = ~(P2_U2546 & P2_INSTQUEUE_REG_3__2__SCAN_IN); 
assign P2_U6971 = ~(P2_U2545 & P2_INSTQUEUE_REG_2__2__SCAN_IN); 
assign P2_U6982 = ~(P2_U2552 & P2_INSTQUEUE_REG_7__1__SCAN_IN); 
assign P2_U6983 = ~(P2_U2551 & P2_INSTQUEUE_REG_6__1__SCAN_IN); 
assign P2_U6986 = ~(P2_U2546 & P2_INSTQUEUE_REG_3__1__SCAN_IN); 
assign P2_U6987 = ~(P2_U2545 & P2_INSTQUEUE_REG_2__1__SCAN_IN); 
assign P2_U6998 = ~(P2_U2552 & P2_INSTQUEUE_REG_7__0__SCAN_IN); 
assign P2_U6999 = ~(P2_U2551 & P2_INSTQUEUE_REG_6__0__SCAN_IN); 
assign P2_U7002 = ~(P2_U2546 & P2_INSTQUEUE_REG_3__0__SCAN_IN); 
assign P2_U7003 = ~(P2_U2545 & P2_INSTQUEUE_REG_2__0__SCAN_IN); 
assign P2_U7016 = ~(P2_U2576 & P2_INSTQUEUE_REG_8__7__SCAN_IN); 
assign P2_U7017 = ~(P2_U2575 & P2_INSTQUEUE_REG_9__7__SCAN_IN); 
assign P2_U7018 = ~(P2_U2574 & P2_INSTQUEUE_REG_10__7__SCAN_IN); 
assign P2_U7019 = ~(P2_U2573 & P2_INSTQUEUE_REG_11__7__SCAN_IN); 
assign P2_U7020 = ~(P2_U2571 & P2_INSTQUEUE_REG_12__7__SCAN_IN); 
assign P2_U7021 = ~(P2_U2569 & P2_INSTQUEUE_REG_13__7__SCAN_IN); 
assign P2_U7022 = ~(P2_U2567 & P2_INSTQUEUE_REG_14__7__SCAN_IN); 
assign P2_U7023 = ~(P2_U2565 & P2_INSTQUEUE_REG_15__7__SCAN_IN); 
assign P2_U7032 = ~(P2_U2576 & P2_INSTQUEUE_REG_8__6__SCAN_IN); 
assign P2_U7033 = ~(P2_U2575 & P2_INSTQUEUE_REG_9__6__SCAN_IN); 
assign P2_U7034 = ~(P2_U2574 & P2_INSTQUEUE_REG_10__6__SCAN_IN); 
assign P2_U7035 = ~(P2_U2573 & P2_INSTQUEUE_REG_11__6__SCAN_IN); 
assign P2_U7036 = ~(P2_U2571 & P2_INSTQUEUE_REG_12__6__SCAN_IN); 
assign P2_U7037 = ~(P2_U2569 & P2_INSTQUEUE_REG_13__6__SCAN_IN); 
assign P2_U7038 = ~(P2_U2567 & P2_INSTQUEUE_REG_14__6__SCAN_IN); 
assign P2_U7039 = ~(P2_U2565 & P2_INSTQUEUE_REG_15__6__SCAN_IN); 
assign P2_U7048 = ~(P2_U2576 & P2_INSTQUEUE_REG_8__5__SCAN_IN); 
assign P2_U7049 = ~(P2_U2575 & P2_INSTQUEUE_REG_9__5__SCAN_IN); 
assign P2_U7050 = ~(P2_U2574 & P2_INSTQUEUE_REG_10__5__SCAN_IN); 
assign P2_U7051 = ~(P2_U2573 & P2_INSTQUEUE_REG_11__5__SCAN_IN); 
assign P2_U7052 = ~(P2_U2571 & P2_INSTQUEUE_REG_12__5__SCAN_IN); 
assign P2_U7053 = ~(P2_U2569 & P2_INSTQUEUE_REG_13__5__SCAN_IN); 
assign P2_U7054 = ~(P2_U2567 & P2_INSTQUEUE_REG_14__5__SCAN_IN); 
assign P2_U7055 = ~(P2_U2565 & P2_INSTQUEUE_REG_15__5__SCAN_IN); 
assign P2_U7064 = ~(P2_U2576 & P2_INSTQUEUE_REG_8__4__SCAN_IN); 
assign P2_U7065 = ~(P2_U2575 & P2_INSTQUEUE_REG_9__4__SCAN_IN); 
assign P2_U7066 = ~(P2_U2574 & P2_INSTQUEUE_REG_10__4__SCAN_IN); 
assign P2_U7067 = ~(P2_U2573 & P2_INSTQUEUE_REG_11__4__SCAN_IN); 
assign P2_U7068 = ~(P2_U2571 & P2_INSTQUEUE_REG_12__4__SCAN_IN); 
assign P2_U7069 = ~(P2_U2569 & P2_INSTQUEUE_REG_13__4__SCAN_IN); 
assign P2_U7070 = ~(P2_U2567 & P2_INSTQUEUE_REG_14__4__SCAN_IN); 
assign P2_U7071 = ~(P2_U2565 & P2_INSTQUEUE_REG_15__4__SCAN_IN); 
assign P2_U7080 = ~(P2_U2576 & P2_INSTQUEUE_REG_8__3__SCAN_IN); 
assign P2_U7081 = ~(P2_U2575 & P2_INSTQUEUE_REG_9__3__SCAN_IN); 
assign P2_U7082 = ~(P2_U2574 & P2_INSTQUEUE_REG_10__3__SCAN_IN); 
assign P2_U7083 = ~(P2_U2573 & P2_INSTQUEUE_REG_11__3__SCAN_IN); 
assign P2_U7084 = ~(P2_U2571 & P2_INSTQUEUE_REG_12__3__SCAN_IN); 
assign P2_U7085 = ~(P2_U2569 & P2_INSTQUEUE_REG_13__3__SCAN_IN); 
assign P2_U7086 = ~(P2_U2567 & P2_INSTQUEUE_REG_14__3__SCAN_IN); 
assign P2_U7087 = ~(P2_U2565 & P2_INSTQUEUE_REG_15__3__SCAN_IN); 
assign P2_U7096 = ~(P2_U2576 & P2_INSTQUEUE_REG_8__2__SCAN_IN); 
assign P2_U7097 = ~(P2_U2575 & P2_INSTQUEUE_REG_9__2__SCAN_IN); 
assign P2_U7098 = ~(P2_U2574 & P2_INSTQUEUE_REG_10__2__SCAN_IN); 
assign P2_U7099 = ~(P2_U2573 & P2_INSTQUEUE_REG_11__2__SCAN_IN); 
assign P2_U7100 = ~(P2_U2571 & P2_INSTQUEUE_REG_12__2__SCAN_IN); 
assign P2_U7101 = ~(P2_U2569 & P2_INSTQUEUE_REG_13__2__SCAN_IN); 
assign P2_U7102 = ~(P2_U2567 & P2_INSTQUEUE_REG_14__2__SCAN_IN); 
assign P2_U7103 = ~(P2_U2565 & P2_INSTQUEUE_REG_15__2__SCAN_IN); 
assign P2_U7112 = ~(P2_U2576 & P2_INSTQUEUE_REG_8__1__SCAN_IN); 
assign P2_U7113 = ~(P2_U2575 & P2_INSTQUEUE_REG_9__1__SCAN_IN); 
assign P2_U7114 = ~(P2_U2574 & P2_INSTQUEUE_REG_10__1__SCAN_IN); 
assign P2_U7115 = ~(P2_U2573 & P2_INSTQUEUE_REG_11__1__SCAN_IN); 
assign P2_U7116 = ~(P2_U2571 & P2_INSTQUEUE_REG_12__1__SCAN_IN); 
assign P2_U7117 = ~(P2_U2569 & P2_INSTQUEUE_REG_13__1__SCAN_IN); 
assign P2_U7118 = ~(P2_U2567 & P2_INSTQUEUE_REG_14__1__SCAN_IN); 
assign P2_U7119 = ~(P2_U2565 & P2_INSTQUEUE_REG_15__1__SCAN_IN); 
assign P2_U7128 = ~(P2_U2576 & P2_INSTQUEUE_REG_8__0__SCAN_IN); 
assign P2_U7129 = ~(P2_U2575 & P2_INSTQUEUE_REG_9__0__SCAN_IN); 
assign P2_U7130 = ~(P2_U2574 & P2_INSTQUEUE_REG_10__0__SCAN_IN); 
assign P2_U7131 = ~(P2_U2573 & P2_INSTQUEUE_REG_11__0__SCAN_IN); 
assign P2_U7132 = ~(P2_U2571 & P2_INSTQUEUE_REG_12__0__SCAN_IN); 
assign P2_U7133 = ~(P2_U2569 & P2_INSTQUEUE_REG_13__0__SCAN_IN); 
assign P2_U7134 = ~(P2_U2567 & P2_INSTQUEUE_REG_14__0__SCAN_IN); 
assign P2_U7135 = ~(P2_U2565 & P2_INSTQUEUE_REG_15__0__SCAN_IN); 
assign P2_U7209 = ~(P2_U2528 & P2_INSTQUEUE_REG_7__6__SCAN_IN); 
assign P2_U7210 = ~(P2_U2527 & P2_INSTQUEUE_REG_6__6__SCAN_IN); 
assign P2_U7211 = ~(P2_U2526 & P2_INSTQUEUE_REG_5__6__SCAN_IN); 
assign P2_U7212 = ~(P2_U2524 & P2_INSTQUEUE_REG_4__6__SCAN_IN); 
assign P2_U7213 = ~(P2_U2522 & P2_INSTQUEUE_REG_3__6__SCAN_IN); 
assign P2_U7214 = ~(P2_U2521 & P2_INSTQUEUE_REG_2__6__SCAN_IN); 
assign P2_U7215 = ~(P2_U2519 & P2_INSTQUEUE_REG_1__6__SCAN_IN); 
assign P2_U7216 = ~(P2_U2517 & P2_INSTQUEUE_REG_0__6__SCAN_IN); 
assign P2_U7243 = ~(P2_U2528 & P2_INSTQUEUE_REG_7__5__SCAN_IN); 
assign P2_U7244 = ~(P2_U2527 & P2_INSTQUEUE_REG_6__5__SCAN_IN); 
assign P2_U7245 = ~(P2_U2526 & P2_INSTQUEUE_REG_5__5__SCAN_IN); 
assign P2_U7246 = ~(P2_U2524 & P2_INSTQUEUE_REG_4__5__SCAN_IN); 
assign P2_U7247 = ~(P2_U2522 & P2_INSTQUEUE_REG_3__5__SCAN_IN); 
assign P2_U7248 = ~(P2_U2521 & P2_INSTQUEUE_REG_2__5__SCAN_IN); 
assign P2_U7249 = ~(P2_U2519 & P2_INSTQUEUE_REG_1__5__SCAN_IN); 
assign P2_U7250 = ~(P2_U2517 & P2_INSTQUEUE_REG_0__5__SCAN_IN); 
assign P2_U7277 = ~(P2_U2528 & P2_INSTQUEUE_REG_7__4__SCAN_IN); 
assign P2_U7278 = ~(P2_U2527 & P2_INSTQUEUE_REG_6__4__SCAN_IN); 
assign P2_U7279 = ~(P2_U2526 & P2_INSTQUEUE_REG_5__4__SCAN_IN); 
assign P2_U7280 = ~(P2_U2524 & P2_INSTQUEUE_REG_4__4__SCAN_IN); 
assign P2_U7281 = ~(P2_U2522 & P2_INSTQUEUE_REG_3__4__SCAN_IN); 
assign P2_U7282 = ~(P2_U2521 & P2_INSTQUEUE_REG_2__4__SCAN_IN); 
assign P2_U7283 = ~(P2_U2519 & P2_INSTQUEUE_REG_1__4__SCAN_IN); 
assign P2_U7284 = ~(P2_U2517 & P2_INSTQUEUE_REG_0__4__SCAN_IN); 
assign P2_U7311 = ~(P2_U2528 & P2_INSTQUEUE_REG_7__3__SCAN_IN); 
assign P2_U7312 = ~(P2_U2527 & P2_INSTQUEUE_REG_6__3__SCAN_IN); 
assign P2_U7313 = ~(P2_U2526 & P2_INSTQUEUE_REG_5__3__SCAN_IN); 
assign P2_U7314 = ~(P2_U2524 & P2_INSTQUEUE_REG_4__3__SCAN_IN); 
assign P2_U7315 = ~(P2_U2522 & P2_INSTQUEUE_REG_3__3__SCAN_IN); 
assign P2_U7316 = ~(P2_U2521 & P2_INSTQUEUE_REG_2__3__SCAN_IN); 
assign P2_U7317 = ~(P2_U2519 & P2_INSTQUEUE_REG_1__3__SCAN_IN); 
assign P2_U7318 = ~(P2_U2517 & P2_INSTQUEUE_REG_0__3__SCAN_IN); 
assign P2_U7345 = ~(P2_U2528 & P2_INSTQUEUE_REG_7__2__SCAN_IN); 
assign P2_U7346 = ~(P2_U2527 & P2_INSTQUEUE_REG_6__2__SCAN_IN); 
assign P2_U7347 = ~(P2_U2526 & P2_INSTQUEUE_REG_5__2__SCAN_IN); 
assign P2_U7348 = ~(P2_U2524 & P2_INSTQUEUE_REG_4__2__SCAN_IN); 
assign P2_U7349 = ~(P2_U2522 & P2_INSTQUEUE_REG_3__2__SCAN_IN); 
assign P2_U7350 = ~(P2_U2521 & P2_INSTQUEUE_REG_2__2__SCAN_IN); 
assign P2_U7351 = ~(P2_U2519 & P2_INSTQUEUE_REG_1__2__SCAN_IN); 
assign P2_U7352 = ~(P2_U2517 & P2_INSTQUEUE_REG_0__2__SCAN_IN); 
assign P2_U7379 = ~(P2_U2528 & P2_INSTQUEUE_REG_7__1__SCAN_IN); 
assign P2_U7380 = ~(P2_U2527 & P2_INSTQUEUE_REG_6__1__SCAN_IN); 
assign P2_U7381 = ~(P2_U2526 & P2_INSTQUEUE_REG_5__1__SCAN_IN); 
assign P2_U7382 = ~(P2_U2524 & P2_INSTQUEUE_REG_4__1__SCAN_IN); 
assign P2_U7383 = ~(P2_U2522 & P2_INSTQUEUE_REG_3__1__SCAN_IN); 
assign P2_U7384 = ~(P2_U2521 & P2_INSTQUEUE_REG_2__1__SCAN_IN); 
assign P2_U7385 = ~(P2_U2519 & P2_INSTQUEUE_REG_1__1__SCAN_IN); 
assign P2_U7386 = ~(P2_U2517 & P2_INSTQUEUE_REG_0__1__SCAN_IN); 
assign P2_U7413 = ~(P2_U2528 & P2_INSTQUEUE_REG_7__0__SCAN_IN); 
assign P2_U7414 = ~(P2_U2527 & P2_INSTQUEUE_REG_6__0__SCAN_IN); 
assign P2_U7415 = ~(P2_U2526 & P2_INSTQUEUE_REG_5__0__SCAN_IN); 
assign P2_U7416 = ~(P2_U2524 & P2_INSTQUEUE_REG_4__0__SCAN_IN); 
assign P2_U7417 = ~(P2_U2522 & P2_INSTQUEUE_REG_3__0__SCAN_IN); 
assign P2_U7418 = ~(P2_U2521 & P2_INSTQUEUE_REG_2__0__SCAN_IN); 
assign P2_U7419 = ~(P2_U2519 & P2_INSTQUEUE_REG_1__0__SCAN_IN); 
assign P2_U7420 = ~(P2_U2517 & P2_INSTQUEUE_REG_0__0__SCAN_IN); 
assign P2_U7431 = ~(P2_U2439 & P2_U3279); 
assign P2_U7537 = ~(P2_U7869 & P2_EBX_REG_9__SCAN_IN); 
assign P2_U7538 = ~(P2_U7869 & P2_EBX_REG_8__SCAN_IN); 
assign P2_U7539 = ~(P2_U7869 & P2_EBX_REG_31__SCAN_IN); 
assign P2_U7540 = ~(P2_U7869 & P2_EBX_REG_30__SCAN_IN); 
assign P2_U7541 = ~(P2_U7869 & P2_EBX_REG_29__SCAN_IN); 
assign P2_U7542 = ~(P2_U7869 & P2_EBX_REG_28__SCAN_IN); 
assign P2_U7543 = ~(P2_U7869 & P2_EBX_REG_27__SCAN_IN); 
assign P2_U7544 = ~(P2_U7869 & P2_EBX_REG_26__SCAN_IN); 
assign P2_U7545 = ~(P2_U7869 & P2_EBX_REG_25__SCAN_IN); 
assign P2_U7546 = ~(P2_U7869 & P2_EBX_REG_24__SCAN_IN); 
assign P2_U7547 = ~(P2_U7869 & P2_EBX_REG_23__SCAN_IN); 
assign P2_U7548 = ~(P2_U7869 & P2_EBX_REG_22__SCAN_IN); 
assign P2_U7549 = ~(P2_U7869 & P2_EBX_REG_21__SCAN_IN); 
assign P2_U7550 = ~(P2_U7869 & P2_EBX_REG_20__SCAN_IN); 
assign P2_U7551 = ~(P2_U7869 & P2_EBX_REG_19__SCAN_IN); 
assign P2_U7552 = ~(P2_U7869 & P2_EBX_REG_18__SCAN_IN); 
assign P2_U7553 = ~(P2_U7869 & P2_EBX_REG_17__SCAN_IN); 
assign P2_U7554 = ~(P2_U7869 & P2_EBX_REG_16__SCAN_IN); 
assign P2_U7555 = ~(P2_U7869 & P2_EBX_REG_15__SCAN_IN); 
assign P2_U7556 = ~(P2_U7869 & P2_EBX_REG_14__SCAN_IN); 
assign P2_U7557 = ~(P2_U7869 & P2_EBX_REG_13__SCAN_IN); 
assign P2_U7558 = ~(P2_U7869 & P2_EBX_REG_12__SCAN_IN); 
assign P2_U7559 = ~(P2_U7869 & P2_EBX_REG_11__SCAN_IN); 
assign P2_U7560 = ~(P2_U7869 & P2_EBX_REG_10__SCAN_IN); 
assign P2_U7732 = ~(P2_R2238_U22 & P2_U2356); 
assign P2_U7734 = ~(P2_R2238_U7 & P2_U2356); 
assign P2_U7738 = ~(P2_U7861 & P2_U2617); 
assign P2_U7745 = ~(P2_U7861 & P2_U2617); 
assign P2_U7895 = ~(P2_U7863 & P2_U7871); 
assign P2_U8075 = ~(P2_U2617 & P2_U3279 & P2_U7859); 
assign P2_U8121 = ~(P2_U7859 & P2_U7873); 
assign P2_U8332 = ~(P2_U7869 & P2_EBX_REG_7__SCAN_IN); 
assign P2_U8334 = ~(P2_U7869 & P2_EBX_REG_6__SCAN_IN); 
assign P2_U8336 = ~(P2_U7869 & P2_EBX_REG_5__SCAN_IN); 
assign P2_U8338 = ~(P2_U7869 & P2_EBX_REG_4__SCAN_IN); 
assign P2_U8340 = ~(P2_U7869 & P2_EBX_REG_3__SCAN_IN); 
assign P2_U8342 = ~(P2_U7869 & P2_EBX_REG_2__SCAN_IN); 
assign P2_U8344 = ~(P2_U7869 & P2_EBX_REG_1__SCAN_IN); 
assign P2_U8346 = ~(P2_U7869 & P2_EBX_REG_0__SCAN_IN); 
assign P1_U2354 = P1_U4265 & P1_U4477; 
assign P1_U2389 = P1_U2452 & P1_U7494; 
assign P1_U2449 = P1_U4494 & P1_U3271; 
assign P1_U2451 = P1_U4251 & P1_STATE2_REG_0__SCAN_IN; 
assign P1_U2546 = P1_U2545 & P1_U2454; 
assign P1_U2547 = P1_U2545 & P1_U3498; 
assign P1_U2548 = P1_U2545 & P1_U4378; 
assign P1_U2549 = P1_U2545 & P1_U2456; 
assign P1_U2551 = P1_U2550 & P1_U2454; 
assign P1_U2552 = P1_U2550 & P1_U3498; 
assign P1_U2553 = P1_U2550 & P1_U4378; 
assign P1_U2554 = P1_U2550 & P1_U2456; 
assign P1_U2584 = P1_U2583 & P1_U2524; 
assign P1_U2585 = P1_U2583 & P1_U2521; 
assign P1_U2586 = P1_U2583 & P1_U2528; 
assign P1_U2587 = P1_U2583 & P1_U2526; 
assign P1_U2589 = P1_U2588 & P1_U2524; 
assign P1_U2590 = P1_U2588 & P1_U2521; 
assign P1_U2591 = P1_U2588 & P1_U2528; 
assign P1_U2592 = P1_U2588 & P1_U2526; 
assign P1_U2603 = P1_U3389 & P1_STATE2_REG_0__SCAN_IN; 
assign P1_U2805 = ~(P1_U7765 & P1_U7764 & P1_U4243); 
assign P1_U3194 = ~(P1_U7647 & P1_U7646 & P1_U4375); 
assign P1_U3196 = ~(P1_U3494 & P1_U4369); 
assign P1_U3282 = ~(P1_U4477 & P1_U3284); 
assign P1_U3287 = ~(P1_U4494 & P1_U4477); 
assign P1_U3289 = ~(P1_U4460 & P1_U3391 & P1_U4173 & P1_U3278); 
assign P1_U3345 = ~(P1_U3341 & P1_U4778); 
assign P1_U3352 = ~(P1_U3349 & P1_U4893); 
assign P1_U3362 = ~(P1_U3356 & P1_U5007); 
assign P1_U3369 = ~(P1_U3366 & P1_U5121); 
assign P1_U3376 = ~(P1_U3373 & P1_U5236); 
assign P1_U3383 = ~(P1_U3380 & P1_U5351); 
assign P1_U3393 = ~(P1_U4399 & P1_U3284); 
assign P1_U3395 = ~(P1_U4399 & P1_U7494 & P1_U4494); 
assign P1_U3397 = ~(P1_U7494 & P1_U4477 & P1_U2605 & P1_U4494 & P1_U4399); 
assign P1_U3398 = ~(P1_U2605 & P1_U4460 & P1_U4171 & P1_U4449 & P1_U4400); 
assign P1_U3409 = ~(P1_U4460 & P1_U3391); 
assign P1_U3418 = ~(P1_U4494 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U3419 = ~(P1_U4399 & P1_U7494); 
assign P1_U3439 = ~(P1_U4449 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U3449 = ~(P1_U4477 & P1_U4496); 
assign P1_U3464 = ~(P1_U7652 & P1_U7651); 
assign P1_U3465 = ~(P1_U7654 & P1_U7653); 
assign P1_U3558 = P1_U3391 & P1_U3283 & P1_U7494; 
assign P1_U3559 = P1_U4460 & P1_U2605 & P1_U4400; 
assign P1_U3577 = P1_U4399 & P1_U4171; 
assign P1_U3579 = P1_U3284 & P1_U3283 & P1_U4400 & P1_U7494; 
assign P1_U3732 = P1_U4494 & P1_U4399; 
assign P1_U3741 = P1_U4449 & P1_U4400; 
assign P1_U3755 = P1_U3284 & P1_U3407; 
assign P1_U3862 = P1_U3283 & P1_U3262 & P1_U7494; 
assign P1_U3885 = P1_U3271 & P1_U7494 & P1_STATE2_REG_0__SCAN_IN; 
assign P1_U3886 = P1_U4399 & P1_U4171; 
assign P1_U3970 = P1_U6621 & P1_U6620 & P1_U6619 & P1_U6618; 
assign P1_U3971 = P1_U6625 & P1_U6624 & P1_U6623 & P1_U6622; 
assign P1_U3974 = P1_U6637 & P1_U6636 & P1_U6635 & P1_U6634; 
assign P1_U3975 = P1_U6641 & P1_U6640 & P1_U6639 & P1_U6638; 
assign P1_U3978 = P1_U6653 & P1_U6652 & P1_U6651 & P1_U6650; 
assign P1_U3979 = P1_U6657 & P1_U6656 & P1_U6655 & P1_U6654; 
assign P1_U3982 = P1_U6669 & P1_U6668 & P1_U6667 & P1_U6666; 
assign P1_U3983 = P1_U6673 & P1_U6672 & P1_U6671 & P1_U6670; 
assign P1_U3986 = P1_U6684 & P1_U6683 & P1_U6682 & P1_U6681; 
assign P1_U3987 = P1_U6688 & P1_U6687 & P1_U6686 & P1_U6685; 
assign P1_U3990 = P1_U6700 & P1_U6699 & P1_U6698 & P1_U6697; 
assign P1_U3991 = P1_U6704 & P1_U6703 & P1_U6702 & P1_U6701; 
assign P1_U3994 = P1_U6716 & P1_U6715 & P1_U6714 & P1_U6713; 
assign P1_U3995 = P1_U6720 & P1_U6719 & P1_U6718 & P1_U6717; 
assign P1_U3998 = P1_U6732 & P1_U6731 & P1_U6730 & P1_U6729; 
assign P1_U3999 = P1_U6736 & P1_U6735 & P1_U6734 & P1_U6733; 
assign P1_U4028 = P1_U7494 & P1_U6888 & P1_U3283; 
assign P1_U4065 = P1_U7077 & P1_U7076 & P1_U7075 & P1_U7074; 
assign P1_U4081 = P1_U7109 & P1_U7108 & P1_U7107 & P1_U7106; 
assign P1_U4085 = P1_U7126 & P1_U7125 & P1_U7124 & P1_U7123; 
assign P1_U4089 = P1_U7143 & P1_U7142 & P1_U7141 & P1_U7140; 
assign P1_U4091 = P1_U7617 & P1_U7146 & P1_U4090; 
assign P1_U4094 = P1_U7158 & P1_U7157 & P1_U7156 & P1_U7155; 
assign P1_U4098 = P1_U7175 & P1_U7174 & P1_U7173 & P1_U7172; 
assign P1_U4102 = P1_U7192 & P1_U7191 & P1_U7190 & P1_U7189; 
assign P1_U4106 = P1_U7209 & P1_U7208 & P1_U7207 & P1_U7206; 
assign P1_U4166 = P1_U3453 & P1_U7384; 
assign P1_U4169 = P1_U7465 & P1_U7464; 
assign P1_U4186 = ~P1_U3412; 
assign P1_U4190 = ~P1_U3290; 
assign P1_U4192 = ~P1_U3405; 
assign P1_U4195 = ~(P1_U4265 & P1_U3271); 
assign P1_U4196 = ~(P1_U4460 & P1_U2605); 
assign P1_U4210 = ~P1_U3390; 
assign P1_U4219 = ~(P1_U4449 & P1_U3271); 
assign P1_U4231 = ~P1_U3407; 
assign P1_U4247 = ~P1_U3394; 
assign P1_U4257 = ~P1_U3389; 
assign P1_U4503 = ~(P1_U4460 & P1_U4173); 
assign P1_U4545 = ~P1_U3322; 
assign P1_U4558 = ~(P1_U3322 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U4616 = ~(P1_U4605 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U4664 = ~P1_U3336; 
assign P1_U4675 = ~(P1_U3336 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U4732 = ~(P1_U4721 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U4836 = ~P1_U3238; 
assign P1_U4842 = ~(P1_U3238 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U4951 = ~P1_U3239; 
assign P1_U4957 = ~(P1_U3239 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U5064 = ~P1_U3240; 
assign P1_U5070 = ~(P1_U3240 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U5179 = ~P1_U3241; 
assign P1_U5185 = ~(P1_U3241 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U5294 = ~P1_U3242; 
assign P1_U5300 = ~(P1_U3242 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U5409 = ~P1_U3243; 
assign P1_U5415 = ~(P1_U3243 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U5463 = ~(P1_U4400 & P1_U4173 & P1_U4460); 
assign P1_U5487 = ~(P1_U4494 & P1_U3290); 
assign P1_U5490 = ~(P1_U4449 & P1_U5488); 
assign P1_U5494 = ~(P1_U4460 & P1_U4171); 
assign P1_U5558 = ~(P1_U4477 & P1_U3272); 
assign P1_U6626 = ~(P1_U2534 & P1_INSTQUEUE_REG_7__7__SCAN_IN); 
assign P1_U6627 = ~(P1_U2533 & P1_INSTQUEUE_REG_6__7__SCAN_IN); 
assign P1_U6628 = ~(P1_U2532 & P1_INSTQUEUE_REG_5__7__SCAN_IN); 
assign P1_U6629 = ~(P1_U2531 & P1_INSTQUEUE_REG_4__7__SCAN_IN); 
assign P1_U6630 = ~(P1_U2529 & P1_INSTQUEUE_REG_3__7__SCAN_IN); 
assign P1_U6631 = ~(P1_U2527 & P1_INSTQUEUE_REG_2__7__SCAN_IN); 
assign P1_U6632 = ~(P1_U2525 & P1_INSTQUEUE_REG_1__7__SCAN_IN); 
assign P1_U6633 = ~(P1_U2523 & P1_INSTQUEUE_REG_0__7__SCAN_IN); 
assign P1_U6642 = ~(P1_U2534 & P1_INSTQUEUE_REG_7__6__SCAN_IN); 
assign P1_U6643 = ~(P1_U2533 & P1_INSTQUEUE_REG_6__6__SCAN_IN); 
assign P1_U6644 = ~(P1_U2532 & P1_INSTQUEUE_REG_5__6__SCAN_IN); 
assign P1_U6645 = ~(P1_U2531 & P1_INSTQUEUE_REG_4__6__SCAN_IN); 
assign P1_U6646 = ~(P1_U2529 & P1_INSTQUEUE_REG_3__6__SCAN_IN); 
assign P1_U6647 = ~(P1_U2527 & P1_INSTQUEUE_REG_2__6__SCAN_IN); 
assign P1_U6648 = ~(P1_U2525 & P1_INSTQUEUE_REG_1__6__SCAN_IN); 
assign P1_U6649 = ~(P1_U2523 & P1_INSTQUEUE_REG_0__6__SCAN_IN); 
assign P1_U6658 = ~(P1_U2534 & P1_INSTQUEUE_REG_7__5__SCAN_IN); 
assign P1_U6659 = ~(P1_U2533 & P1_INSTQUEUE_REG_6__5__SCAN_IN); 
assign P1_U6660 = ~(P1_U2532 & P1_INSTQUEUE_REG_5__5__SCAN_IN); 
assign P1_U6661 = ~(P1_U2531 & P1_INSTQUEUE_REG_4__5__SCAN_IN); 
assign P1_U6662 = ~(P1_U2529 & P1_INSTQUEUE_REG_3__5__SCAN_IN); 
assign P1_U6663 = ~(P1_U2527 & P1_INSTQUEUE_REG_2__5__SCAN_IN); 
assign P1_U6664 = ~(P1_U2525 & P1_INSTQUEUE_REG_1__5__SCAN_IN); 
assign P1_U6665 = ~(P1_U2523 & P1_INSTQUEUE_REG_0__5__SCAN_IN); 
assign P1_U6674 = ~(P1_U2534 & P1_INSTQUEUE_REG_7__4__SCAN_IN); 
assign P1_U6675 = ~(P1_U2533 & P1_INSTQUEUE_REG_6__4__SCAN_IN); 
assign P1_U6676 = ~(P1_U2532 & P1_INSTQUEUE_REG_5__4__SCAN_IN); 
assign P1_U6677 = ~(P1_U2531 & P1_INSTQUEUE_REG_4__4__SCAN_IN); 
assign P1_U6678 = ~(P1_U2529 & P1_INSTQUEUE_REG_3__4__SCAN_IN); 
assign P1_U6679 = ~(P1_U2527 & P1_INSTQUEUE_REG_2__4__SCAN_IN); 
assign P1_U6680 = ~(P1_U2525 & P1_INSTQUEUE_REG_1__4__SCAN_IN); 
assign P1_U6689 = ~(P1_U2534 & P1_INSTQUEUE_REG_7__3__SCAN_IN); 
assign P1_U6690 = ~(P1_U2533 & P1_INSTQUEUE_REG_6__3__SCAN_IN); 
assign P1_U6691 = ~(P1_U2532 & P1_INSTQUEUE_REG_5__3__SCAN_IN); 
assign P1_U6692 = ~(P1_U2531 & P1_INSTQUEUE_REG_4__3__SCAN_IN); 
assign P1_U6693 = ~(P1_U2529 & P1_INSTQUEUE_REG_3__3__SCAN_IN); 
assign P1_U6694 = ~(P1_U2527 & P1_INSTQUEUE_REG_2__3__SCAN_IN); 
assign P1_U6695 = ~(P1_U2525 & P1_INSTQUEUE_REG_1__3__SCAN_IN); 
assign P1_U6696 = ~(P1_U2523 & P1_INSTQUEUE_REG_0__3__SCAN_IN); 
assign P1_U6705 = ~(P1_U2534 & P1_INSTQUEUE_REG_7__2__SCAN_IN); 
assign P1_U6706 = ~(P1_U2533 & P1_INSTQUEUE_REG_6__2__SCAN_IN); 
assign P1_U6707 = ~(P1_U2532 & P1_INSTQUEUE_REG_5__2__SCAN_IN); 
assign P1_U6708 = ~(P1_U2531 & P1_INSTQUEUE_REG_4__2__SCAN_IN); 
assign P1_U6709 = ~(P1_U2529 & P1_INSTQUEUE_REG_3__2__SCAN_IN); 
assign P1_U6710 = ~(P1_U2527 & P1_INSTQUEUE_REG_2__2__SCAN_IN); 
assign P1_U6711 = ~(P1_U2525 & P1_INSTQUEUE_REG_1__2__SCAN_IN); 
assign P1_U6712 = ~(P1_U2523 & P1_INSTQUEUE_REG_0__2__SCAN_IN); 
assign P1_U6721 = ~(P1_U2534 & P1_INSTQUEUE_REG_7__1__SCAN_IN); 
assign P1_U6722 = ~(P1_U2533 & P1_INSTQUEUE_REG_6__1__SCAN_IN); 
assign P1_U6723 = ~(P1_U2532 & P1_INSTQUEUE_REG_5__1__SCAN_IN); 
assign P1_U6724 = ~(P1_U2531 & P1_INSTQUEUE_REG_4__1__SCAN_IN); 
assign P1_U6725 = ~(P1_U2529 & P1_INSTQUEUE_REG_3__1__SCAN_IN); 
assign P1_U6726 = ~(P1_U2527 & P1_INSTQUEUE_REG_2__1__SCAN_IN); 
assign P1_U6727 = ~(P1_U2525 & P1_INSTQUEUE_REG_1__1__SCAN_IN); 
assign P1_U6728 = ~(P1_U2523 & P1_INSTQUEUE_REG_0__1__SCAN_IN); 
assign P1_U6737 = ~(P1_U2534 & P1_INSTQUEUE_REG_7__0__SCAN_IN); 
assign P1_U6738 = ~(P1_U2533 & P1_INSTQUEUE_REG_6__0__SCAN_IN); 
assign P1_U6739 = ~(P1_U2532 & P1_INSTQUEUE_REG_5__0__SCAN_IN); 
assign P1_U6740 = ~(P1_U2531 & P1_INSTQUEUE_REG_4__0__SCAN_IN); 
assign P1_U6741 = ~(P1_U2529 & P1_INSTQUEUE_REG_3__0__SCAN_IN); 
assign P1_U6742 = ~(P1_U2527 & P1_INSTQUEUE_REG_2__0__SCAN_IN); 
assign P1_U6743 = ~(P1_U2525 & P1_INSTQUEUE_REG_1__0__SCAN_IN); 
assign P1_U6744 = ~(P1_U2523 & P1_INSTQUEUE_REG_0__0__SCAN_IN); 
assign P1_U6745 = ~(P1_U4460 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U6885 = ~(P1_U4494 & P1_U3283); 
assign P1_U6891 = ~(P1_U4494 & P1_U3283); 
assign P1_U6892 = ~(P1_U2564 & P1_INSTQUEUE_REG_15__1__SCAN_IN); 
assign P1_U6893 = ~(P1_U2563 & P1_INSTQUEUE_REG_14__1__SCAN_IN); 
assign P1_U6894 = ~(P1_U2562 & P1_INSTQUEUE_REG_13__1__SCAN_IN); 
assign P1_U6895 = ~(P1_U2561 & P1_INSTQUEUE_REG_12__1__SCAN_IN); 
assign P1_U6896 = ~(P1_U2559 & P1_INSTQUEUE_REG_11__1__SCAN_IN); 
assign P1_U6897 = ~(P1_U2558 & P1_INSTQUEUE_REG_10__1__SCAN_IN); 
assign P1_U6898 = ~(P1_U2557 & P1_INSTQUEUE_REG_9__1__SCAN_IN); 
assign P1_U6899 = ~(P1_U2556 & P1_INSTQUEUE_REG_8__1__SCAN_IN); 
assign P1_U6910 = ~(P1_U2564 & P1_INSTQUEUE_REG_15__0__SCAN_IN); 
assign P1_U6911 = ~(P1_U2563 & P1_INSTQUEUE_REG_14__0__SCAN_IN); 
assign P1_U6912 = ~(P1_U2562 & P1_INSTQUEUE_REG_13__0__SCAN_IN); 
assign P1_U6913 = ~(P1_U2561 & P1_INSTQUEUE_REG_12__0__SCAN_IN); 
assign P1_U6914 = ~(P1_U2559 & P1_INSTQUEUE_REG_11__0__SCAN_IN); 
assign P1_U6915 = ~(P1_U2558 & P1_INSTQUEUE_REG_10__0__SCAN_IN); 
assign P1_U6916 = ~(P1_U2557 & P1_INSTQUEUE_REG_9__0__SCAN_IN); 
assign P1_U6917 = ~(P1_U2556 & P1_INSTQUEUE_REG_8__0__SCAN_IN); 
assign P1_U6941 = ~(P1_U2564 & P1_INSTQUEUE_REG_15__7__SCAN_IN); 
assign P1_U6942 = ~(P1_U2563 & P1_INSTQUEUE_REG_14__7__SCAN_IN); 
assign P1_U6943 = ~(P1_U2562 & P1_INSTQUEUE_REG_13__7__SCAN_IN); 
assign P1_U6944 = ~(P1_U2561 & P1_INSTQUEUE_REG_12__7__SCAN_IN); 
assign P1_U6945 = ~(P1_U2559 & P1_INSTQUEUE_REG_11__7__SCAN_IN); 
assign P1_U6946 = ~(P1_U2558 & P1_INSTQUEUE_REG_10__7__SCAN_IN); 
assign P1_U6947 = ~(P1_U2557 & P1_INSTQUEUE_REG_9__7__SCAN_IN); 
assign P1_U6948 = ~(P1_U2556 & P1_INSTQUEUE_REG_8__7__SCAN_IN); 
assign P1_U6958 = ~(P1_U2564 & P1_INSTQUEUE_REG_15__6__SCAN_IN); 
assign P1_U6959 = ~(P1_U2563 & P1_INSTQUEUE_REG_14__6__SCAN_IN); 
assign P1_U6960 = ~(P1_U2562 & P1_INSTQUEUE_REG_13__6__SCAN_IN); 
assign P1_U6961 = ~(P1_U2561 & P1_INSTQUEUE_REG_12__6__SCAN_IN); 
assign P1_U6962 = ~(P1_U2559 & P1_INSTQUEUE_REG_11__6__SCAN_IN); 
assign P1_U6963 = ~(P1_U2558 & P1_INSTQUEUE_REG_10__6__SCAN_IN); 
assign P1_U6964 = ~(P1_U2557 & P1_INSTQUEUE_REG_9__6__SCAN_IN); 
assign P1_U6965 = ~(P1_U2556 & P1_INSTQUEUE_REG_8__6__SCAN_IN); 
assign P1_U6975 = ~(P1_U2564 & P1_INSTQUEUE_REG_15__5__SCAN_IN); 
assign P1_U6976 = ~(P1_U2563 & P1_INSTQUEUE_REG_14__5__SCAN_IN); 
assign P1_U6977 = ~(P1_U2562 & P1_INSTQUEUE_REG_13__5__SCAN_IN); 
assign P1_U6978 = ~(P1_U2561 & P1_INSTQUEUE_REG_12__5__SCAN_IN); 
assign P1_U6979 = ~(P1_U2559 & P1_INSTQUEUE_REG_11__5__SCAN_IN); 
assign P1_U6980 = ~(P1_U2558 & P1_INSTQUEUE_REG_10__5__SCAN_IN); 
assign P1_U6981 = ~(P1_U2557 & P1_INSTQUEUE_REG_9__5__SCAN_IN); 
assign P1_U6982 = ~(P1_U2556 & P1_INSTQUEUE_REG_8__5__SCAN_IN); 
assign P1_U6992 = ~(P1_U2564 & P1_INSTQUEUE_REG_15__4__SCAN_IN); 
assign P1_U6993 = ~(P1_U2563 & P1_INSTQUEUE_REG_14__4__SCAN_IN); 
assign P1_U6994 = ~(P1_U2562 & P1_INSTQUEUE_REG_13__4__SCAN_IN); 
assign P1_U6995 = ~(P1_U2561 & P1_INSTQUEUE_REG_12__4__SCAN_IN); 
assign P1_U6996 = ~(P1_U2559 & P1_INSTQUEUE_REG_11__4__SCAN_IN); 
assign P1_U6997 = ~(P1_U2558 & P1_INSTQUEUE_REG_10__4__SCAN_IN); 
assign P1_U6998 = ~(P1_U2557 & P1_INSTQUEUE_REG_9__4__SCAN_IN); 
assign P1_U6999 = ~(P1_U2556 & P1_INSTQUEUE_REG_8__4__SCAN_IN); 
assign P1_U7007 = ~(P1_U2564 & P1_INSTQUEUE_REG_15__3__SCAN_IN); 
assign P1_U7008 = ~(P1_U2563 & P1_INSTQUEUE_REG_14__3__SCAN_IN); 
assign P1_U7009 = ~(P1_U2562 & P1_INSTQUEUE_REG_13__3__SCAN_IN); 
assign P1_U7010 = ~(P1_U2561 & P1_INSTQUEUE_REG_12__3__SCAN_IN); 
assign P1_U7011 = ~(P1_U2559 & P1_INSTQUEUE_REG_11__3__SCAN_IN); 
assign P1_U7012 = ~(P1_U2558 & P1_INSTQUEUE_REG_10__3__SCAN_IN); 
assign P1_U7013 = ~(P1_U2557 & P1_INSTQUEUE_REG_9__3__SCAN_IN); 
assign P1_U7014 = ~(P1_U2556 & P1_INSTQUEUE_REG_8__3__SCAN_IN); 
assign P1_U7024 = ~(P1_U2564 & P1_INSTQUEUE_REG_15__2__SCAN_IN); 
assign P1_U7025 = ~(P1_U2563 & P1_INSTQUEUE_REG_14__2__SCAN_IN); 
assign P1_U7026 = ~(P1_U2562 & P1_INSTQUEUE_REG_13__2__SCAN_IN); 
assign P1_U7027 = ~(P1_U2561 & P1_INSTQUEUE_REG_12__2__SCAN_IN); 
assign P1_U7028 = ~(P1_U2559 & P1_INSTQUEUE_REG_11__2__SCAN_IN); 
assign P1_U7029 = ~(P1_U2558 & P1_INSTQUEUE_REG_10__2__SCAN_IN); 
assign P1_U7030 = ~(P1_U2557 & P1_INSTQUEUE_REG_9__2__SCAN_IN); 
assign P1_U7031 = ~(P1_U2556 & P1_INSTQUEUE_REG_8__2__SCAN_IN); 
assign P1_U7220 = ~(P1_U2602 & P1_INSTQUEUE_REG_8__7__SCAN_IN); 
assign P1_U7221 = ~(P1_U2601 & P1_INSTQUEUE_REG_9__7__SCAN_IN); 
assign P1_U7222 = ~(P1_U2600 & P1_INSTQUEUE_REG_10__7__SCAN_IN); 
assign P1_U7223 = ~(P1_U2599 & P1_INSTQUEUE_REG_11__7__SCAN_IN); 
assign P1_U7224 = ~(P1_U2597 & P1_INSTQUEUE_REG_12__7__SCAN_IN); 
assign P1_U7225 = ~(P1_U2596 & P1_INSTQUEUE_REG_13__7__SCAN_IN); 
assign P1_U7226 = ~(P1_U2595 & P1_INSTQUEUE_REG_14__7__SCAN_IN); 
assign P1_U7227 = ~(P1_U2594 & P1_INSTQUEUE_REG_15__7__SCAN_IN); 
assign P1_U7237 = ~(P1_U2602 & P1_INSTQUEUE_REG_8__6__SCAN_IN); 
assign P1_U7238 = ~(P1_U2601 & P1_INSTQUEUE_REG_9__6__SCAN_IN); 
assign P1_U7239 = ~(P1_U2600 & P1_INSTQUEUE_REG_10__6__SCAN_IN); 
assign P1_U7240 = ~(P1_U2599 & P1_INSTQUEUE_REG_11__6__SCAN_IN); 
assign P1_U7241 = ~(P1_U2597 & P1_INSTQUEUE_REG_12__6__SCAN_IN); 
assign P1_U7242 = ~(P1_U2596 & P1_INSTQUEUE_REG_13__6__SCAN_IN); 
assign P1_U7243 = ~(P1_U2595 & P1_INSTQUEUE_REG_14__6__SCAN_IN); 
assign P1_U7244 = ~(P1_U2594 & P1_INSTQUEUE_REG_15__6__SCAN_IN); 
assign P1_U7254 = ~(P1_U2602 & P1_INSTQUEUE_REG_8__5__SCAN_IN); 
assign P1_U7255 = ~(P1_U2601 & P1_INSTQUEUE_REG_9__5__SCAN_IN); 
assign P1_U7256 = ~(P1_U2600 & P1_INSTQUEUE_REG_10__5__SCAN_IN); 
assign P1_U7257 = ~(P1_U2599 & P1_INSTQUEUE_REG_11__5__SCAN_IN); 
assign P1_U7258 = ~(P1_U2597 & P1_INSTQUEUE_REG_12__5__SCAN_IN); 
assign P1_U7259 = ~(P1_U2596 & P1_INSTQUEUE_REG_13__5__SCAN_IN); 
assign P1_U7260 = ~(P1_U2595 & P1_INSTQUEUE_REG_14__5__SCAN_IN); 
assign P1_U7261 = ~(P1_U2594 & P1_INSTQUEUE_REG_15__5__SCAN_IN); 
assign P1_U7271 = ~(P1_U2602 & P1_INSTQUEUE_REG_8__4__SCAN_IN); 
assign P1_U7272 = ~(P1_U2601 & P1_INSTQUEUE_REG_9__4__SCAN_IN); 
assign P1_U7273 = ~(P1_U2600 & P1_INSTQUEUE_REG_10__4__SCAN_IN); 
assign P1_U7274 = ~(P1_U2599 & P1_INSTQUEUE_REG_11__4__SCAN_IN); 
assign P1_U7275 = ~(P1_U2597 & P1_INSTQUEUE_REG_12__4__SCAN_IN); 
assign P1_U7276 = ~(P1_U2596 & P1_INSTQUEUE_REG_13__4__SCAN_IN); 
assign P1_U7277 = ~(P1_U2595 & P1_INSTQUEUE_REG_14__4__SCAN_IN); 
assign P1_U7278 = ~(P1_U2594 & P1_INSTQUEUE_REG_15__4__SCAN_IN); 
assign P1_U7286 = ~(P1_U2602 & P1_INSTQUEUE_REG_8__3__SCAN_IN); 
assign P1_U7287 = ~(P1_U2601 & P1_INSTQUEUE_REG_9__3__SCAN_IN); 
assign P1_U7288 = ~(P1_U2600 & P1_INSTQUEUE_REG_10__3__SCAN_IN); 
assign P1_U7289 = ~(P1_U2599 & P1_INSTQUEUE_REG_11__3__SCAN_IN); 
assign P1_U7290 = ~(P1_U2597 & P1_INSTQUEUE_REG_12__3__SCAN_IN); 
assign P1_U7291 = ~(P1_U2596 & P1_INSTQUEUE_REG_13__3__SCAN_IN); 
assign P1_U7292 = ~(P1_U2595 & P1_INSTQUEUE_REG_14__3__SCAN_IN); 
assign P1_U7293 = ~(P1_U2594 & P1_INSTQUEUE_REG_15__3__SCAN_IN); 
assign P1_U7303 = ~(P1_U2602 & P1_INSTQUEUE_REG_8__2__SCAN_IN); 
assign P1_U7304 = ~(P1_U2601 & P1_INSTQUEUE_REG_9__2__SCAN_IN); 
assign P1_U7305 = ~(P1_U2600 & P1_INSTQUEUE_REG_10__2__SCAN_IN); 
assign P1_U7306 = ~(P1_U2599 & P1_INSTQUEUE_REG_11__2__SCAN_IN); 
assign P1_U7307 = ~(P1_U2597 & P1_INSTQUEUE_REG_12__2__SCAN_IN); 
assign P1_U7308 = ~(P1_U2596 & P1_INSTQUEUE_REG_13__2__SCAN_IN); 
assign P1_U7309 = ~(P1_U2595 & P1_INSTQUEUE_REG_14__2__SCAN_IN); 
assign P1_U7310 = ~(P1_U2594 & P1_INSTQUEUE_REG_15__2__SCAN_IN); 
assign P1_U7320 = ~(P1_U2602 & P1_INSTQUEUE_REG_8__1__SCAN_IN); 
assign P1_U7321 = ~(P1_U2601 & P1_INSTQUEUE_REG_9__1__SCAN_IN); 
assign P1_U7322 = ~(P1_U2600 & P1_INSTQUEUE_REG_10__1__SCAN_IN); 
assign P1_U7323 = ~(P1_U2599 & P1_INSTQUEUE_REG_11__1__SCAN_IN); 
assign P1_U7324 = ~(P1_U2597 & P1_INSTQUEUE_REG_12__1__SCAN_IN); 
assign P1_U7325 = ~(P1_U2596 & P1_INSTQUEUE_REG_13__1__SCAN_IN); 
assign P1_U7326 = ~(P1_U2595 & P1_INSTQUEUE_REG_14__1__SCAN_IN); 
assign P1_U7327 = ~(P1_U2594 & P1_INSTQUEUE_REG_15__1__SCAN_IN); 
assign P1_U7337 = ~(P1_U2602 & P1_INSTQUEUE_REG_8__0__SCAN_IN); 
assign P1_U7338 = ~(P1_U2601 & P1_INSTQUEUE_REG_9__0__SCAN_IN); 
assign P1_U7339 = ~(P1_U2600 & P1_INSTQUEUE_REG_10__0__SCAN_IN); 
assign P1_U7340 = ~(P1_U2599 & P1_INSTQUEUE_REG_11__0__SCAN_IN); 
assign P1_U7341 = ~(P1_U2597 & P1_INSTQUEUE_REG_12__0__SCAN_IN); 
assign P1_U7342 = ~(P1_U2596 & P1_INSTQUEUE_REG_13__0__SCAN_IN); 
assign P1_U7343 = ~(P1_U2595 & P1_INSTQUEUE_REG_14__0__SCAN_IN); 
assign P1_U7344 = ~(P1_U2594 & P1_INSTQUEUE_REG_15__0__SCAN_IN); 
assign P1_U7456 = ~(P1_U4477 & P1_U4496); 
assign P1_U7613 = ~(P1_U2523 & P1_INSTQUEUE_REG_0__4__SCAN_IN); 
assign P1_U7703 = ~(P1_U4460 & P1_U3278); 
assign P1_U7785 = ~(P1_U4460 & P1_U7495); 
assign P3_ADD_526_U53 = ~(P3_ADD_526_U146 & P3_ADD_526_U145); 
assign P3_ADD_526_U54 = ~(P3_ADD_526_U148 & P3_ADD_526_U147); 
assign P3_ADD_526_U120 = ~P3_ADD_526_U17; 
assign P3_ADD_526_U125 = ~P3_ADD_526_U95; 
assign P3_ADD_526_U142 = ~(P3_ADD_526_U17 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_526_U143 = ~(P3_ADD_526_U95 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_552_U53 = ~(P3_ADD_552_U146 & P3_ADD_552_U145); 
assign P3_ADD_552_U54 = ~(P3_ADD_552_U148 & P3_ADD_552_U147); 
assign P3_ADD_552_U120 = ~P3_ADD_552_U17; 
assign P3_ADD_552_U125 = ~P3_ADD_552_U95; 
assign P3_ADD_552_U142 = ~(P3_ADD_552_U17 & P3_EBX_REG_9__SCAN_IN); 
assign P3_ADD_552_U143 = ~(P3_ADD_552_U95 & P3_EBX_REG_8__SCAN_IN); 
assign P3_ADD_546_U53 = ~(P3_ADD_546_U146 & P3_ADD_546_U145); 
assign P3_ADD_546_U54 = ~(P3_ADD_546_U148 & P3_ADD_546_U147); 
assign P3_ADD_546_U120 = ~P3_ADD_546_U17; 
assign P3_ADD_546_U125 = ~P3_ADD_546_U95; 
assign P3_ADD_546_U142 = ~(P3_ADD_546_U17 & P3_EAX_REG_9__SCAN_IN); 
assign P3_ADD_546_U143 = ~(P3_ADD_546_U95 & P3_EAX_REG_8__SCAN_IN); 
assign P3_ADD_476_U66 = ~(P3_ADD_476_U132 & P3_ADD_476_U131); 
assign P3_ADD_476_U97 = ~P3_ADD_476_U12; 
assign P3_ADD_476_U129 = ~(P3_ADD_476_U12 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_531_U70 = ~(P3_ADD_531_U139 & P3_ADD_531_U138); 
assign P3_ADD_531_U101 = ~P3_ADD_531_U13; 
assign P3_ADD_531_U136 = ~(P3_ADD_531_U13 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_SUB_320_U22 = ~(P3_SUB_320_U27 & P3_SUB_320_U58 & P3_SUB_320_U83); 
assign P3_ADD_505_U14 = ~(P3_ADD_505_U22 & P3_ADD_505_U21); 
assign P3_ADD_318_U66 = ~(P3_ADD_318_U132 & P3_ADD_318_U131); 
assign P3_ADD_318_U97 = ~P3_ADD_318_U12; 
assign P3_ADD_318_U129 = ~(P3_ADD_318_U12 & P3_PHYADDRPOINTER_REG_6__SCAN_IN); 
assign P3_SUB_370_U27 = ~(P3_SUB_370_U37 & P3_SUB_370_U36); 
assign P3_SUB_370_U60 = ~(P3_SUB_370_U34 & P3_SUB_370_U59); 
assign P3_ADD_315_U63 = ~(P3_ADD_315_U126 & P3_ADD_315_U125); 
assign P3_ADD_315_U94 = ~P3_ADD_315_U12; 
assign P3_ADD_315_U123 = ~(P3_ADD_315_U12 & P3_PHYADDRPOINTER_REG_7__SCAN_IN); 
assign P3_SUB_589_U9 = ~P3_U3300; 
assign P3_ADD_467_U66 = ~(P3_ADD_467_U132 & P3_ADD_467_U131); 
assign P3_ADD_467_U97 = ~P3_ADD_467_U12; 
assign P3_ADD_467_U129 = ~(P3_ADD_467_U12 & P3_REIP_REG_6__SCAN_IN); 
assign P3_ADD_430_U66 = ~(P3_ADD_430_U132 & P3_ADD_430_U131); 
assign P3_ADD_430_U97 = ~P3_ADD_430_U12; 
assign P3_ADD_430_U129 = ~(P3_ADD_430_U12 & P3_REIP_REG_6__SCAN_IN); 
assign P3_ADD_380_U70 = ~(P3_ADD_380_U139 & P3_ADD_380_U138); 
assign P3_ADD_380_U101 = ~P3_ADD_380_U13; 
assign P3_ADD_380_U136 = ~(P3_ADD_380_U13 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_344_U70 = ~(P3_ADD_344_U139 & P3_ADD_344_U138); 
assign P3_ADD_344_U101 = ~P3_ADD_344_U13; 
assign P3_ADD_344_U136 = ~(P3_ADD_344_U13 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_339_U66 = ~(P3_ADD_339_U132 & P3_ADD_339_U131); 
assign P3_ADD_339_U97 = ~P3_ADD_339_U12; 
assign P3_ADD_339_U129 = ~(P3_ADD_339_U12 & P3_PHYADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_541_U66 = ~(P3_ADD_541_U132 & P3_ADD_541_U131); 
assign P3_ADD_541_U97 = ~P3_ADD_541_U12; 
assign P3_ADD_541_U129 = ~(P3_ADD_541_U12 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_SUB_355_U27 = ~(P3_SUB_355_U37 & P3_SUB_355_U36); 
assign P3_SUB_355_U60 = ~(P3_SUB_355_U34 & P3_SUB_355_U59); 
assign P3_SUB_450_U24 = ~(P3_SUB_450_U35 & P3_SUB_450_U34); 
assign P3_SUB_450_U57 = ~(P3_SUB_450_U32 & P3_SUB_450_U56); 
assign P3_ADD_486_U14 = ~(P3_ADD_486_U22 & P3_ADD_486_U21); 
assign P3_SUB_485_U24 = ~(P3_SUB_485_U35 & P3_SUB_485_U34); 
assign P3_SUB_485_U57 = ~(P3_SUB_485_U32 & P3_SUB_485_U56); 
assign P3_ADD_515_U66 = ~(P3_ADD_515_U132 & P3_ADD_515_U131); 
assign P3_ADD_515_U97 = ~P3_ADD_515_U12; 
assign P3_ADD_515_U129 = ~(P3_ADD_515_U12 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_394_U67 = ~(P3_ADD_394_U136 & P3_ADD_394_U135); 
assign P3_ADD_394_U100 = ~P3_ADD_394_U12; 
assign P3_ADD_394_U133 = ~(P3_ADD_394_U12 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_SUB_414_U55 = P3_SUB_414_U131 & P3_SUB_414_U130; 
assign P3_SUB_414_U86 = ~P3_SUB_414_U24; 
assign P3_SUB_414_U88 = ~(P3_SUB_414_U87 & P3_EBX_REG_8__SCAN_IN); 
assign P3_SUB_414_U128 = ~(P3_SUB_414_U24 & P3_EBX_REG_9__SCAN_IN); 
assign P3_ADD_441_U66 = ~(P3_ADD_441_U132 & P3_ADD_441_U131); 
assign P3_ADD_441_U97 = ~P3_ADD_441_U12; 
assign P3_ADD_441_U129 = ~(P3_ADD_441_U12 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_349_U70 = ~(P3_ADD_349_U139 & P3_ADD_349_U138); 
assign P3_ADD_349_U101 = ~P3_ADD_349_U13; 
assign P3_ADD_349_U136 = ~(P3_ADD_349_U13 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_405_U67 = ~(P3_ADD_405_U136 & P3_ADD_405_U135); 
assign P3_ADD_405_U100 = ~P3_ADD_405_U12; 
assign P3_ADD_405_U133 = ~(P3_ADD_405_U12 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_553_U70 = ~(P3_ADD_553_U139 & P3_ADD_553_U138); 
assign P3_ADD_553_U101 = ~P3_ADD_553_U13; 
assign P3_ADD_553_U136 = ~(P3_ADD_553_U13 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_558_U70 = ~(P3_ADD_558_U139 & P3_ADD_558_U138); 
assign P3_ADD_558_U101 = ~P3_ADD_558_U13; 
assign P3_ADD_558_U136 = ~(P3_ADD_558_U13 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_385_U70 = ~(P3_ADD_385_U139 & P3_ADD_385_U138); 
assign P3_ADD_385_U101 = ~P3_ADD_385_U13; 
assign P3_ADD_385_U136 = ~(P3_ADD_385_U13 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_547_U70 = ~(P3_ADD_547_U139 & P3_ADD_547_U138); 
assign P3_ADD_547_U101 = ~P3_ADD_547_U13; 
assign P3_ADD_547_U136 = ~(P3_ADD_547_U13 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_SUB_412_U24 = ~(P3_SUB_412_U35 & P3_SUB_412_U34); 
assign P3_SUB_412_U57 = ~(P3_SUB_412_U32 & P3_SUB_412_U56); 
assign P3_SUB_504_U24 = ~(P3_SUB_504_U35 & P3_SUB_504_U34); 
assign P3_SUB_504_U57 = ~(P3_SUB_504_U32 & P3_SUB_504_U56); 
assign P3_SUB_401_U27 = ~(P3_SUB_401_U37 & P3_SUB_401_U36); 
assign P3_SUB_401_U60 = ~(P3_SUB_401_U34 & P3_SUB_401_U59); 
assign P3_SUB_390_U27 = ~(P3_SUB_390_U37 & P3_SUB_390_U36); 
assign P3_SUB_390_U60 = ~(P3_SUB_390_U34 & P3_SUB_390_U59); 
assign P3_ADD_494_U66 = ~(P3_ADD_494_U132 & P3_ADD_494_U131); 
assign P3_ADD_494_U97 = ~P3_ADD_494_U12; 
assign P3_ADD_494_U129 = ~(P3_ADD_494_U12 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_536_U66 = ~(P3_ADD_536_U132 & P3_ADD_536_U131); 
assign P3_ADD_536_U97 = ~P3_ADD_536_U12; 
assign P3_ADD_536_U129 = ~(P3_ADD_536_U12 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P2_R2027_U70 = ~(P2_R2027_U139 & P2_R2027_U138); 
assign P2_R2027_U101 = ~P2_R2027_U13; 
assign P2_R2027_U136 = ~(P2_R2027_U13 & P2_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P2_R2337_U64 = ~(P2_R2337_U130 & P2_R2337_U129); 
assign P2_R2337_U98 = ~P2_R2337_U13; 
assign P2_R2337_U127 = ~(P2_R2337_U13 & P2_PHYADDRPOINTER_REG_7__SCAN_IN); 
assign P2_R2238_U27 = ~(P2_R2238_U37 & P2_R2238_U36); 
assign P2_R2238_U60 = ~(P2_R2238_U34 & P2_R2238_U59); 
assign P2_R1957_U22 = ~(P2_R1957_U51 & P2_R1957_U83); 
assign P2_R1957_U91 = ~(P2_R1957_U83 & P2_R1957_U58); 
assign P2_R1957_U135 = ~(P2_R1957_U83 & P2_R1957_U58); 
assign P2_SUB_450_U25 = ~(P2_SUB_450_U35 & P2_SUB_450_U34); 
assign P2_SUB_450_U57 = ~(P2_SUB_450_U32 & P2_SUB_450_U56); 
assign P2_ADD_394_U79 = ~(P2_ADD_394_U160 & P2_ADD_394_U159); 
assign P2_ADD_394_U100 = ~P2_ADD_394_U13; 
assign P2_ADD_394_U127 = ~(P2_ADD_394_U13 & P2_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P2_ADD_371_1212_U106 = P2_ADD_371_1212_U12 & P2_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P2_ADD_371_1212_U107 = P2_ADD_371_1212_U12 & P2_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P1_R2027_U53 = ~(P1_R2027_U146 & P1_R2027_U145); 
assign P1_R2027_U54 = ~(P1_R2027_U148 & P1_R2027_U147); 
assign P1_R2027_U120 = ~P1_R2027_U17; 
assign P1_R2027_U125 = ~P1_R2027_U95; 
assign P1_R2027_U142 = ~(P1_R2027_U17 & P1_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P1_R2027_U143 = ~(P1_R2027_U95 & P1_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P1_R2337_U66 = ~(P1_R2337_U132 & P1_R2337_U131); 
assign P1_R2337_U97 = ~P1_R2337_U12; 
assign P1_R2337_U129 = ~(P1_R2337_U12 & P1_PHYADDRPOINTER_REG_6__SCAN_IN); 
assign P1_R2096_U66 = ~(P1_R2096_U132 & P1_R2096_U131); 
assign P1_R2096_U97 = ~P1_R2096_U12; 
assign P1_R2096_U129 = ~(P1_R2096_U12 & P1_REIP_REG_6__SCAN_IN); 
assign P1_R2238_U27 = ~(P1_R2238_U37 & P1_R2238_U36); 
assign P1_R2238_U60 = ~(P1_R2238_U34 & P1_R2238_U59); 
assign P1_SUB_450_U27 = ~(P1_SUB_450_U37 & P1_SUB_450_U36); 
assign P1_SUB_450_U60 = ~(P1_SUB_450_U34 & P1_SUB_450_U59); 
assign P1_ADD_405_U79 = ~(P1_ADD_405_U160 & P1_ADD_405_U159); 
assign P1_ADD_405_U100 = ~P1_ADD_405_U13; 
assign P1_ADD_405_U127 = ~(P1_ADD_405_U13 & P1_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P1_ADD_515_U79 = ~(P1_ADD_515_U158 & P1_ADD_515_U157); 
assign P1_ADD_515_U97 = ~P1_ADD_515_U13; 
assign P1_ADD_515_U123 = ~(P1_ADD_515_U13 & P1_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign U216 = ~(U483 & U484 & U482); 
assign U217 = ~(U480 & U481 & U479); 
assign U218 = ~(U477 & U478 & U476); 
assign U219 = ~(U474 & U475 & U473); 
assign U220 = ~(U471 & U472 & U470); 
assign U221 = ~(U468 & U469 & U467); 
assign U222 = ~(U465 & U466 & U464); 
assign U223 = ~(U462 & U463 & U461); 
assign U224 = ~(U459 & U460 & U458); 
assign U225 = ~(U456 & U457 & U455); 
assign U226 = ~(U453 & U454 & U452); 
assign U227 = ~(U450 & U451 & U449); 
assign U228 = ~(U447 & U448 & U446); 
assign U229 = ~(U444 & U445 & U443); 
assign U230 = ~(U441 & U442 & U440); 
assign U231 = ~(U438 & U439 & U437); 
assign U232 = ~(U435 & U436 & U434); 
assign U233 = ~(U432 & U433 & U431); 
assign U234 = ~(U429 & U430 & U428); 
assign U235 = ~(U426 & U427 & U425); 
assign U236 = ~(U423 & U424 & U422); 
assign U237 = ~(U420 & U421 & U419); 
assign U238 = ~(U417 & U418 & U416); 
assign U239 = ~(U414 & U415 & U413); 
assign U240 = ~(U411 & U412 & U410); 
assign U241 = ~(U408 & U409 & U407); 
assign U242 = ~(U405 & U406 & U404); 
assign U243 = ~(U402 & U403 & U401); 
assign U244 = ~(U399 & U400 & U398); 
assign U245 = ~(U396 & U397 & U395); 
assign U246 = ~(U393 & U394 & U392); 
assign U247 = ~(U390 & U391 & U389); 
assign P3_U2437 = P3_U2381 & P3_U3108; 
assign P3_U2438 = P3_U2381 & P3_U3104; 
assign P3_U2439 = P3_U2381 & P3_U3101; 
assign P3_U2440 = P3_U2381 & P3_U3107; 
assign P3_U2441 = P3_U2381 & P3_U3102; 
assign P3_U2442 = P3_U2381 & P3_U3110; 
assign P3_U2443 = P3_U2381 & P3_U3074; 
assign P3_U2445 = P3_U2381 & P3_U3218; 
assign P3_U2613 = ~(P3_U4279 & P3_U4278 & P3_U4277 & P3_U4276); 
assign P3_U2614 = ~(P3_U4275 & P3_U4274 & P3_U4273 & P3_U4272); 
assign P3_U2615 = ~(P3_U4271 & P3_U4270 & P3_U4269 & P3_U4268); 
assign P3_U2616 = ~(P3_U4267 & P3_U4266 & P3_U4265 & P3_U4264); 
assign P3_U2617 = ~(P3_U4263 & P3_U4262 & P3_U4261 & P3_U4260); 
assign P3_U2618 = ~(P3_U4259 & P3_U4258 & P3_U4257 & P3_U4256); 
assign P3_U2619 = ~(P3_U4255 & P3_U4254 & P3_U4253 & P3_U4252); 
assign P3_U2620 = ~(P3_U4251 & P3_U4250 & P3_U4249 & P3_U4248); 
assign P3_U3072 = ~(P3_U2458 & P3_U4642); 
assign P3_U3073 = ~(P3_U2460 & P3_U4642); 
assign P3_U3103 = ~(P3_U3074 & P3_U3110); 
assign P3_U3111 = ~(P3_U3104 & P3_U3108); 
assign P3_U3146 = ~(P3_U3134 & P3_U4663); 
assign P3_U3152 = ~(P3_U3147 & P3_U4717); 
assign P3_U3156 = ~(P3_U3148 & P3_U3155); 
assign P3_U3160 = ~(P3_U3154 & P3_U4769); 
assign P3_U3168 = ~(P3_U3164 & P3_U4872); 
assign P3_U3172 = ~(P3_U3169 & P3_U4924); 
assign P3_U3176 = ~(P3_U3173 & P3_U4976); 
assign P3_U3235 = ~(P3_U3101 & P3_U3104 & P3_U4294); 
assign P3_U3360 = P3_U3107 & P3_U3108 & P3_U3218; 
assign P3_U3686 = P3_U5594 & P3_U5592; 
assign P3_U3951 = P3_U3104 & P3_STATE2_REG_0__SCAN_IN; 
assign P3_U4152 = P3_U7390 & P3_U7389 & P3_U7388 & P3_U7387; 
assign P3_U4153 = P3_U7394 & P3_U7393 & P3_U7392 & P3_U7391; 
assign P3_U4156 = P3_U7406 & P3_U7405 & P3_U7404 & P3_U7403; 
assign P3_U4157 = P3_U7410 & P3_U7409 & P3_U7408 & P3_U7407; 
assign P3_U4160 = P3_U7422 & P3_U7421 & P3_U7420 & P3_U7419; 
assign P3_U4161 = P3_U7426 & P3_U7425 & P3_U7424 & P3_U7423; 
assign P3_U4164 = P3_U7438 & P3_U7437 & P3_U7436 & P3_U7435; 
assign P3_U4165 = P3_U7442 & P3_U7441 & P3_U7440 & P3_U7439; 
assign P3_U4168 = P3_U7454 & P3_U7453 & P3_U7452 & P3_U7451; 
assign P3_U4169 = P3_U7458 & P3_U7457 & P3_U7456 & P3_U7455; 
assign P3_U4172 = P3_U7470 & P3_U7469 & P3_U7468 & P3_U7467; 
assign P3_U4173 = P3_U7474 & P3_U7473 & P3_U7472 & P3_U7471; 
assign P3_U4176 = P3_U7486 & P3_U7485 & P3_U7484 & P3_U7483; 
assign P3_U4177 = P3_U7490 & P3_U7489 & P3_U7488 & P3_U7487; 
assign P3_U4180 = P3_U7502 & P3_U7501 & P3_U7500 & P3_U7499; 
assign P3_U4181 = P3_U7506 & P3_U7505 & P3_U7504 & P3_U7503; 
assign P3_U4186 = P3_U7528 & P3_U7527 & P3_U7526 & P3_U7525; 
assign P3_U4187 = P3_U7532 & P3_U7531 & P3_U7530 & P3_U7529; 
assign P3_U4190 = P3_U7544 & P3_U7543 & P3_U7542 & P3_U7541; 
assign P3_U4191 = P3_U7548 & P3_U7547 & P3_U7546 & P3_U7545; 
assign P3_U4194 = P3_U7560 & P3_U7559 & P3_U7558 & P3_U7557; 
assign P3_U4195 = P3_U7564 & P3_U7563 & P3_U7562 & P3_U7561; 
assign P3_U4198 = P3_U7576 & P3_U7575 & P3_U7574 & P3_U7573; 
assign P3_U4199 = P3_U7580 & P3_U7579 & P3_U7578 & P3_U7577; 
assign P3_U4202 = P3_U7592 & P3_U7591 & P3_U7590 & P3_U7589; 
assign P3_U4203 = P3_U7596 & P3_U7595 & P3_U7594 & P3_U7593; 
assign P3_U4206 = P3_U7608 & P3_U7607 & P3_U7606 & P3_U7605; 
assign P3_U4207 = P3_U7612 & P3_U7611 & P3_U7610 & P3_U7609; 
assign P3_U4210 = P3_U7624 & P3_U7623 & P3_U7622 & P3_U7621; 
assign P3_U4211 = P3_U7628 & P3_U7627 & P3_U7626 & P3_U7625; 
assign P3_U4214 = P3_U7640 & P3_U7639 & P3_U7638 & P3_U7637; 
assign P3_U4215 = P3_U7644 & P3_U7643 & P3_U7642 & P3_U7641; 
assign P3_U4216 = P3_U7649 & P3_U7648 & P3_U7647 & P3_U7646; 
assign P3_U4217 = P3_U7653 & P3_U7652 & P3_U7651 & P3_U7650; 
assign P3_U4220 = P3_U7665 & P3_U7664 & P3_U7663 & P3_U7662; 
assign P3_U4221 = P3_U7669 & P3_U7668 & P3_U7667 & P3_U7666; 
assign P3_U4224 = P3_U7681 & P3_U7680 & P3_U7679 & P3_U7678; 
assign P3_U4225 = P3_U7685 & P3_U7684 & P3_U7683 & P3_U7682; 
assign P3_U4228 = P3_U7697 & P3_U7696 & P3_U7695 & P3_U7694; 
assign P3_U4229 = P3_U7701 & P3_U7700 & P3_U7699 & P3_U7698; 
assign P3_U4232 = P3_U7713 & P3_U7712 & P3_U7711 & P3_U7710; 
assign P3_U4233 = P3_U7717 & P3_U7716 & P3_U7715 & P3_U7714; 
assign P3_U4236 = P3_U7729 & P3_U7728 & P3_U7727 & P3_U7726; 
assign P3_U4237 = P3_U7733 & P3_U7732 & P3_U7731 & P3_U7730; 
assign P3_U4240 = P3_U7745 & P3_U7744 & P3_U7743 & P3_U7742; 
assign P3_U4241 = P3_U7749 & P3_U7748 & P3_U7747 & P3_U7746; 
assign P3_U4244 = P3_U7761 & P3_U7760 & P3_U7759 & P3_U7758; 
assign P3_U4245 = P3_U7765 & P3_U7764 & P3_U7763 & P3_U7762; 
assign P3_U4331 = ~(P3_U2458 & P3_U4653); 
assign P3_U4488 = ~P3_U3108; 
assign P3_U4505 = ~P3_U3104; 
assign P3_U4522 = ~P3_U3102; 
assign P3_U4539 = ~P3_U3101; 
assign P3_U4556 = ~P3_U3107; 
assign P3_U4573 = ~P3_U3218; 
assign P3_U4590 = ~P3_U3110; 
assign P3_U4607 = ~P3_U3074; 
assign P3_U4645 = ~P3_U3155; 
assign P3_U4821 = ~P3_U3070; 
assign P3_U5028 = ~P3_U3071; 
assign P3_U5128 = ~(P3_U4342 & P3_U2458); 
assign P3_U5180 = ~(P3_U4343 & P3_U2458); 
assign P3_U5282 = ~(P3_U2460 & P3_U4653); 
assign P3_U5333 = ~(P3_U2460 & P3_U4342); 
assign P3_U5384 = ~(P3_U2460 & P3_U4343); 
assign P3_U7395 = ~(P3_U2532 & P3_INSTQUEUE_REG_7__7__SCAN_IN); 
assign P3_U7396 = ~(P3_U2531 & P3_INSTQUEUE_REG_6__7__SCAN_IN); 
assign P3_U7397 = ~(P3_U2530 & P3_INSTQUEUE_REG_5__7__SCAN_IN); 
assign P3_U7398 = ~(P3_U2529 & P3_INSTQUEUE_REG_4__7__SCAN_IN); 
assign P3_U7399 = ~(P3_U2527 & P3_INSTQUEUE_REG_3__7__SCAN_IN); 
assign P3_U7400 = ~(P3_U2525 & P3_INSTQUEUE_REG_2__7__SCAN_IN); 
assign P3_U7401 = ~(P3_U2523 & P3_INSTQUEUE_REG_1__7__SCAN_IN); 
assign P3_U7402 = ~(P3_U2521 & P3_INSTQUEUE_REG_0__7__SCAN_IN); 
assign P3_U7411 = ~(P3_U2532 & P3_INSTQUEUE_REG_7__6__SCAN_IN); 
assign P3_U7412 = ~(P3_U2531 & P3_INSTQUEUE_REG_6__6__SCAN_IN); 
assign P3_U7413 = ~(P3_U2530 & P3_INSTQUEUE_REG_5__6__SCAN_IN); 
assign P3_U7414 = ~(P3_U2529 & P3_INSTQUEUE_REG_4__6__SCAN_IN); 
assign P3_U7415 = ~(P3_U2527 & P3_INSTQUEUE_REG_3__6__SCAN_IN); 
assign P3_U7416 = ~(P3_U2525 & P3_INSTQUEUE_REG_2__6__SCAN_IN); 
assign P3_U7417 = ~(P3_U2523 & P3_INSTQUEUE_REG_1__6__SCAN_IN); 
assign P3_U7418 = ~(P3_U2521 & P3_INSTQUEUE_REG_0__6__SCAN_IN); 
assign P3_U7427 = ~(P3_U2532 & P3_INSTQUEUE_REG_7__5__SCAN_IN); 
assign P3_U7428 = ~(P3_U2531 & P3_INSTQUEUE_REG_6__5__SCAN_IN); 
assign P3_U7429 = ~(P3_U2530 & P3_INSTQUEUE_REG_5__5__SCAN_IN); 
assign P3_U7430 = ~(P3_U2529 & P3_INSTQUEUE_REG_4__5__SCAN_IN); 
assign P3_U7431 = ~(P3_U2527 & P3_INSTQUEUE_REG_3__5__SCAN_IN); 
assign P3_U7432 = ~(P3_U2525 & P3_INSTQUEUE_REG_2__5__SCAN_IN); 
assign P3_U7433 = ~(P3_U2523 & P3_INSTQUEUE_REG_1__5__SCAN_IN); 
assign P3_U7434 = ~(P3_U2521 & P3_INSTQUEUE_REG_0__5__SCAN_IN); 
assign P3_U7443 = ~(P3_U2532 & P3_INSTQUEUE_REG_7__4__SCAN_IN); 
assign P3_U7444 = ~(P3_U2531 & P3_INSTQUEUE_REG_6__4__SCAN_IN); 
assign P3_U7445 = ~(P3_U2530 & P3_INSTQUEUE_REG_5__4__SCAN_IN); 
assign P3_U7446 = ~(P3_U2529 & P3_INSTQUEUE_REG_4__4__SCAN_IN); 
assign P3_U7447 = ~(P3_U2527 & P3_INSTQUEUE_REG_3__4__SCAN_IN); 
assign P3_U7448 = ~(P3_U2525 & P3_INSTQUEUE_REG_2__4__SCAN_IN); 
assign P3_U7449 = ~(P3_U2523 & P3_INSTQUEUE_REG_1__4__SCAN_IN); 
assign P3_U7450 = ~(P3_U2521 & P3_INSTQUEUE_REG_0__4__SCAN_IN); 
assign P3_U7459 = ~(P3_U2532 & P3_INSTQUEUE_REG_7__3__SCAN_IN); 
assign P3_U7460 = ~(P3_U2531 & P3_INSTQUEUE_REG_6__3__SCAN_IN); 
assign P3_U7461 = ~(P3_U2530 & P3_INSTQUEUE_REG_5__3__SCAN_IN); 
assign P3_U7462 = ~(P3_U2529 & P3_INSTQUEUE_REG_4__3__SCAN_IN); 
assign P3_U7463 = ~(P3_U2527 & P3_INSTQUEUE_REG_3__3__SCAN_IN); 
assign P3_U7464 = ~(P3_U2525 & P3_INSTQUEUE_REG_2__3__SCAN_IN); 
assign P3_U7465 = ~(P3_U2523 & P3_INSTQUEUE_REG_1__3__SCAN_IN); 
assign P3_U7466 = ~(P3_U2521 & P3_INSTQUEUE_REG_0__3__SCAN_IN); 
assign P3_U7475 = ~(P3_U2532 & P3_INSTQUEUE_REG_7__2__SCAN_IN); 
assign P3_U7476 = ~(P3_U2531 & P3_INSTQUEUE_REG_6__2__SCAN_IN); 
assign P3_U7477 = ~(P3_U2530 & P3_INSTQUEUE_REG_5__2__SCAN_IN); 
assign P3_U7478 = ~(P3_U2529 & P3_INSTQUEUE_REG_4__2__SCAN_IN); 
assign P3_U7479 = ~(P3_U2527 & P3_INSTQUEUE_REG_3__2__SCAN_IN); 
assign P3_U7480 = ~(P3_U2525 & P3_INSTQUEUE_REG_2__2__SCAN_IN); 
assign P3_U7481 = ~(P3_U2523 & P3_INSTQUEUE_REG_1__2__SCAN_IN); 
assign P3_U7482 = ~(P3_U2521 & P3_INSTQUEUE_REG_0__2__SCAN_IN); 
assign P3_U7491 = ~(P3_U2532 & P3_INSTQUEUE_REG_7__1__SCAN_IN); 
assign P3_U7492 = ~(P3_U2531 & P3_INSTQUEUE_REG_6__1__SCAN_IN); 
assign P3_U7493 = ~(P3_U2530 & P3_INSTQUEUE_REG_5__1__SCAN_IN); 
assign P3_U7494 = ~(P3_U2529 & P3_INSTQUEUE_REG_4__1__SCAN_IN); 
assign P3_U7495 = ~(P3_U2527 & P3_INSTQUEUE_REG_3__1__SCAN_IN); 
assign P3_U7496 = ~(P3_U2525 & P3_INSTQUEUE_REG_2__1__SCAN_IN); 
assign P3_U7497 = ~(P3_U2523 & P3_INSTQUEUE_REG_1__1__SCAN_IN); 
assign P3_U7498 = ~(P3_U2521 & P3_INSTQUEUE_REG_0__1__SCAN_IN); 
assign P3_U7507 = ~(P3_U2532 & P3_INSTQUEUE_REG_7__0__SCAN_IN); 
assign P3_U7508 = ~(P3_U2531 & P3_INSTQUEUE_REG_6__0__SCAN_IN); 
assign P3_U7509 = ~(P3_U2530 & P3_INSTQUEUE_REG_5__0__SCAN_IN); 
assign P3_U7510 = ~(P3_U2529 & P3_INSTQUEUE_REG_4__0__SCAN_IN); 
assign P3_U7511 = ~(P3_U2527 & P3_INSTQUEUE_REG_3__0__SCAN_IN); 
assign P3_U7512 = ~(P3_U2525 & P3_INSTQUEUE_REG_2__0__SCAN_IN); 
assign P3_U7513 = ~(P3_U2523 & P3_INSTQUEUE_REG_1__0__SCAN_IN); 
assign P3_U7514 = ~(P3_U2521 & P3_INSTQUEUE_REG_0__0__SCAN_IN); 
assign P3_U7517 = ~(P3_U2562 & P3_INSTQUEUE_REG_0__7__SCAN_IN); 
assign P3_U7518 = ~(P3_U2561 & P3_INSTQUEUE_REG_1__7__SCAN_IN); 
assign P3_U7519 = ~(P3_U2560 & P3_INSTQUEUE_REG_2__7__SCAN_IN); 
assign P3_U7520 = ~(P3_U2559 & P3_INSTQUEUE_REG_3__7__SCAN_IN); 
assign P3_U7521 = ~(P3_U2557 & P3_INSTQUEUE_REG_4__7__SCAN_IN); 
assign P3_U7522 = ~(P3_U2556 & P3_INSTQUEUE_REG_5__7__SCAN_IN); 
assign P3_U7523 = ~(P3_U2555 & P3_INSTQUEUE_REG_6__7__SCAN_IN); 
assign P3_U7524 = ~(P3_U2554 & P3_INSTQUEUE_REG_7__7__SCAN_IN); 
assign P3_U7533 = ~(P3_U2562 & P3_INSTQUEUE_REG_0__6__SCAN_IN); 
assign P3_U7534 = ~(P3_U2561 & P3_INSTQUEUE_REG_1__6__SCAN_IN); 
assign P3_U7535 = ~(P3_U2560 & P3_INSTQUEUE_REG_2__6__SCAN_IN); 
assign P3_U7536 = ~(P3_U2559 & P3_INSTQUEUE_REG_3__6__SCAN_IN); 
assign P3_U7537 = ~(P3_U2557 & P3_INSTQUEUE_REG_4__6__SCAN_IN); 
assign P3_U7538 = ~(P3_U2556 & P3_INSTQUEUE_REG_5__6__SCAN_IN); 
assign P3_U7539 = ~(P3_U2555 & P3_INSTQUEUE_REG_6__6__SCAN_IN); 
assign P3_U7540 = ~(P3_U2554 & P3_INSTQUEUE_REG_7__6__SCAN_IN); 
assign P3_U7549 = ~(P3_U2562 & P3_INSTQUEUE_REG_0__5__SCAN_IN); 
assign P3_U7550 = ~(P3_U2561 & P3_INSTQUEUE_REG_1__5__SCAN_IN); 
assign P3_U7551 = ~(P3_U2560 & P3_INSTQUEUE_REG_2__5__SCAN_IN); 
assign P3_U7552 = ~(P3_U2559 & P3_INSTQUEUE_REG_3__5__SCAN_IN); 
assign P3_U7553 = ~(P3_U2557 & P3_INSTQUEUE_REG_4__5__SCAN_IN); 
assign P3_U7554 = ~(P3_U2556 & P3_INSTQUEUE_REG_5__5__SCAN_IN); 
assign P3_U7555 = ~(P3_U2555 & P3_INSTQUEUE_REG_6__5__SCAN_IN); 
assign P3_U7556 = ~(P3_U2554 & P3_INSTQUEUE_REG_7__5__SCAN_IN); 
assign P3_U7565 = ~(P3_U2562 & P3_INSTQUEUE_REG_0__4__SCAN_IN); 
assign P3_U7566 = ~(P3_U2561 & P3_INSTQUEUE_REG_1__4__SCAN_IN); 
assign P3_U7567 = ~(P3_U2560 & P3_INSTQUEUE_REG_2__4__SCAN_IN); 
assign P3_U7568 = ~(P3_U2559 & P3_INSTQUEUE_REG_3__4__SCAN_IN); 
assign P3_U7569 = ~(P3_U2557 & P3_INSTQUEUE_REG_4__4__SCAN_IN); 
assign P3_U7570 = ~(P3_U2556 & P3_INSTQUEUE_REG_5__4__SCAN_IN); 
assign P3_U7571 = ~(P3_U2555 & P3_INSTQUEUE_REG_6__4__SCAN_IN); 
assign P3_U7572 = ~(P3_U2554 & P3_INSTQUEUE_REG_7__4__SCAN_IN); 
assign P3_U7581 = ~(P3_U2562 & P3_INSTQUEUE_REG_0__3__SCAN_IN); 
assign P3_U7582 = ~(P3_U2561 & P3_INSTQUEUE_REG_1__3__SCAN_IN); 
assign P3_U7583 = ~(P3_U2560 & P3_INSTQUEUE_REG_2__3__SCAN_IN); 
assign P3_U7584 = ~(P3_U2559 & P3_INSTQUEUE_REG_3__3__SCAN_IN); 
assign P3_U7585 = ~(P3_U2557 & P3_INSTQUEUE_REG_4__3__SCAN_IN); 
assign P3_U7586 = ~(P3_U2556 & P3_INSTQUEUE_REG_5__3__SCAN_IN); 
assign P3_U7587 = ~(P3_U2555 & P3_INSTQUEUE_REG_6__3__SCAN_IN); 
assign P3_U7588 = ~(P3_U2554 & P3_INSTQUEUE_REG_7__3__SCAN_IN); 
assign P3_U7597 = ~(P3_U2562 & P3_INSTQUEUE_REG_0__2__SCAN_IN); 
assign P3_U7598 = ~(P3_U2561 & P3_INSTQUEUE_REG_1__2__SCAN_IN); 
assign P3_U7599 = ~(P3_U2560 & P3_INSTQUEUE_REG_2__2__SCAN_IN); 
assign P3_U7600 = ~(P3_U2559 & P3_INSTQUEUE_REG_3__2__SCAN_IN); 
assign P3_U7601 = ~(P3_U2557 & P3_INSTQUEUE_REG_4__2__SCAN_IN); 
assign P3_U7602 = ~(P3_U2556 & P3_INSTQUEUE_REG_5__2__SCAN_IN); 
assign P3_U7603 = ~(P3_U2555 & P3_INSTQUEUE_REG_6__2__SCAN_IN); 
assign P3_U7604 = ~(P3_U2554 & P3_INSTQUEUE_REG_7__2__SCAN_IN); 
assign P3_U7613 = ~(P3_U2562 & P3_INSTQUEUE_REG_0__1__SCAN_IN); 
assign P3_U7614 = ~(P3_U2561 & P3_INSTQUEUE_REG_1__1__SCAN_IN); 
assign P3_U7615 = ~(P3_U2560 & P3_INSTQUEUE_REG_2__1__SCAN_IN); 
assign P3_U7616 = ~(P3_U2559 & P3_INSTQUEUE_REG_3__1__SCAN_IN); 
assign P3_U7617 = ~(P3_U2557 & P3_INSTQUEUE_REG_4__1__SCAN_IN); 
assign P3_U7618 = ~(P3_U2556 & P3_INSTQUEUE_REG_5__1__SCAN_IN); 
assign P3_U7619 = ~(P3_U2555 & P3_INSTQUEUE_REG_6__1__SCAN_IN); 
assign P3_U7620 = ~(P3_U2554 & P3_INSTQUEUE_REG_7__1__SCAN_IN); 
assign P3_U7629 = ~(P3_U2562 & P3_INSTQUEUE_REG_0__0__SCAN_IN); 
assign P3_U7630 = ~(P3_U2561 & P3_INSTQUEUE_REG_1__0__SCAN_IN); 
assign P3_U7631 = ~(P3_U2560 & P3_INSTQUEUE_REG_2__0__SCAN_IN); 
assign P3_U7632 = ~(P3_U2559 & P3_INSTQUEUE_REG_3__0__SCAN_IN); 
assign P3_U7633 = ~(P3_U2557 & P3_INSTQUEUE_REG_4__0__SCAN_IN); 
assign P3_U7634 = ~(P3_U2556 & P3_INSTQUEUE_REG_5__0__SCAN_IN); 
assign P3_U7635 = ~(P3_U2555 & P3_INSTQUEUE_REG_6__0__SCAN_IN); 
assign P3_U7636 = ~(P3_U2554 & P3_INSTQUEUE_REG_7__0__SCAN_IN); 
assign P3_U7654 = ~(P3_U2572 & P3_INSTQUEUE_REG_0__7__SCAN_IN); 
assign P3_U7655 = ~(P3_U2571 & P3_INSTQUEUE_REG_1__7__SCAN_IN); 
assign P3_U7656 = ~(P3_U2570 & P3_INSTQUEUE_REG_2__7__SCAN_IN); 
assign P3_U7657 = ~(P3_U2569 & P3_INSTQUEUE_REG_3__7__SCAN_IN); 
assign P3_U7658 = ~(P3_U2567 & P3_INSTQUEUE_REG_4__7__SCAN_IN); 
assign P3_U7659 = ~(P3_U2566 & P3_INSTQUEUE_REG_5__7__SCAN_IN); 
assign P3_U7660 = ~(P3_U2565 & P3_INSTQUEUE_REG_6__7__SCAN_IN); 
assign P3_U7661 = ~(P3_U2564 & P3_INSTQUEUE_REG_7__7__SCAN_IN); 
assign P3_U7670 = ~(P3_U2572 & P3_INSTQUEUE_REG_0__6__SCAN_IN); 
assign P3_U7671 = ~(P3_U2571 & P3_INSTQUEUE_REG_1__6__SCAN_IN); 
assign P3_U7672 = ~(P3_U2570 & P3_INSTQUEUE_REG_2__6__SCAN_IN); 
assign P3_U7673 = ~(P3_U2569 & P3_INSTQUEUE_REG_3__6__SCAN_IN); 
assign P3_U7674 = ~(P3_U2567 & P3_INSTQUEUE_REG_4__6__SCAN_IN); 
assign P3_U7675 = ~(P3_U2566 & P3_INSTQUEUE_REG_5__6__SCAN_IN); 
assign P3_U7676 = ~(P3_U2565 & P3_INSTQUEUE_REG_6__6__SCAN_IN); 
assign P3_U7677 = ~(P3_U2564 & P3_INSTQUEUE_REG_7__6__SCAN_IN); 
assign P3_U7686 = ~(P3_U2572 & P3_INSTQUEUE_REG_0__5__SCAN_IN); 
assign P3_U7687 = ~(P3_U2571 & P3_INSTQUEUE_REG_1__5__SCAN_IN); 
assign P3_U7688 = ~(P3_U2570 & P3_INSTQUEUE_REG_2__5__SCAN_IN); 
assign P3_U7689 = ~(P3_U2569 & P3_INSTQUEUE_REG_3__5__SCAN_IN); 
assign P3_U7690 = ~(P3_U2567 & P3_INSTQUEUE_REG_4__5__SCAN_IN); 
assign P3_U7691 = ~(P3_U2566 & P3_INSTQUEUE_REG_5__5__SCAN_IN); 
assign P3_U7692 = ~(P3_U2565 & P3_INSTQUEUE_REG_6__5__SCAN_IN); 
assign P3_U7693 = ~(P3_U2564 & P3_INSTQUEUE_REG_7__5__SCAN_IN); 
assign P3_U7702 = ~(P3_U2572 & P3_INSTQUEUE_REG_0__4__SCAN_IN); 
assign P3_U7703 = ~(P3_U2571 & P3_INSTQUEUE_REG_1__4__SCAN_IN); 
assign P3_U7704 = ~(P3_U2570 & P3_INSTQUEUE_REG_2__4__SCAN_IN); 
assign P3_U7705 = ~(P3_U2569 & P3_INSTQUEUE_REG_3__4__SCAN_IN); 
assign P3_U7706 = ~(P3_U2567 & P3_INSTQUEUE_REG_4__4__SCAN_IN); 
assign P3_U7707 = ~(P3_U2566 & P3_INSTQUEUE_REG_5__4__SCAN_IN); 
assign P3_U7708 = ~(P3_U2565 & P3_INSTQUEUE_REG_6__4__SCAN_IN); 
assign P3_U7709 = ~(P3_U2564 & P3_INSTQUEUE_REG_7__4__SCAN_IN); 
assign P3_U7718 = ~(P3_U2572 & P3_INSTQUEUE_REG_0__3__SCAN_IN); 
assign P3_U7719 = ~(P3_U2571 & P3_INSTQUEUE_REG_1__3__SCAN_IN); 
assign P3_U7720 = ~(P3_U2570 & P3_INSTQUEUE_REG_2__3__SCAN_IN); 
assign P3_U7721 = ~(P3_U2569 & P3_INSTQUEUE_REG_3__3__SCAN_IN); 
assign P3_U7722 = ~(P3_U2567 & P3_INSTQUEUE_REG_4__3__SCAN_IN); 
assign P3_U7723 = ~(P3_U2566 & P3_INSTQUEUE_REG_5__3__SCAN_IN); 
assign P3_U7724 = ~(P3_U2565 & P3_INSTQUEUE_REG_6__3__SCAN_IN); 
assign P3_U7725 = ~(P3_U2564 & P3_INSTQUEUE_REG_7__3__SCAN_IN); 
assign P3_U7734 = ~(P3_U2572 & P3_INSTQUEUE_REG_0__2__SCAN_IN); 
assign P3_U7735 = ~(P3_U2571 & P3_INSTQUEUE_REG_1__2__SCAN_IN); 
assign P3_U7736 = ~(P3_U2570 & P3_INSTQUEUE_REG_2__2__SCAN_IN); 
assign P3_U7737 = ~(P3_U2569 & P3_INSTQUEUE_REG_3__2__SCAN_IN); 
assign P3_U7738 = ~(P3_U2567 & P3_INSTQUEUE_REG_4__2__SCAN_IN); 
assign P3_U7739 = ~(P3_U2566 & P3_INSTQUEUE_REG_5__2__SCAN_IN); 
assign P3_U7740 = ~(P3_U2565 & P3_INSTQUEUE_REG_6__2__SCAN_IN); 
assign P3_U7741 = ~(P3_U2564 & P3_INSTQUEUE_REG_7__2__SCAN_IN); 
assign P3_U7750 = ~(P3_U2572 & P3_INSTQUEUE_REG_0__1__SCAN_IN); 
assign P3_U7751 = ~(P3_U2571 & P3_INSTQUEUE_REG_1__1__SCAN_IN); 
assign P3_U7752 = ~(P3_U2570 & P3_INSTQUEUE_REG_2__1__SCAN_IN); 
assign P3_U7753 = ~(P3_U2569 & P3_INSTQUEUE_REG_3__1__SCAN_IN); 
assign P3_U7754 = ~(P3_U2567 & P3_INSTQUEUE_REG_4__1__SCAN_IN); 
assign P3_U7755 = ~(P3_U2566 & P3_INSTQUEUE_REG_5__1__SCAN_IN); 
assign P3_U7756 = ~(P3_U2565 & P3_INSTQUEUE_REG_6__1__SCAN_IN); 
assign P3_U7757 = ~(P3_U2564 & P3_INSTQUEUE_REG_7__1__SCAN_IN); 
assign P3_U7766 = ~(P3_U2572 & P3_INSTQUEUE_REG_0__0__SCAN_IN); 
assign P3_U7767 = ~(P3_U2571 & P3_INSTQUEUE_REG_1__0__SCAN_IN); 
assign P3_U7768 = ~(P3_U2570 & P3_INSTQUEUE_REG_2__0__SCAN_IN); 
assign P3_U7769 = ~(P3_U2569 & P3_INSTQUEUE_REG_3__0__SCAN_IN); 
assign P3_U7770 = ~(P3_U2567 & P3_INSTQUEUE_REG_4__0__SCAN_IN); 
assign P3_U7771 = ~(P3_U2566 & P3_INSTQUEUE_REG_5__0__SCAN_IN); 
assign P3_U7772 = ~(P3_U2565 & P3_INSTQUEUE_REG_6__0__SCAN_IN); 
assign P3_U7773 = ~(P3_U2564 & P3_INSTQUEUE_REG_7__0__SCAN_IN); 
assign P3_U7966 = ~(P3_U7965 & P3_U4657); 
assign P3_U7973 = ~(P3_U3218 & P3_U3107); 
assign P2_U2353 = P2_U4343 & P2_U2439; 
assign P2_U2357 = P2_U3712 & P2_U2458; 
assign P2_U2376 = P2_U3873 & P2_U2436; 
assign P2_U2450 = P2_U2354 & P2_U7871; 
assign P2_U2658 = P2_U2354 & P2_U2598; 
assign P2_U2659 = P2_U2354 & P2_U2597; 
assign P2_U2660 = P2_U2354 & P2_U2596; 
assign P2_U2661 = P2_U2354 & P2_U2595; 
assign P2_U2662 = P2_U2354 & P2_U2594; 
assign P2_U2663 = P2_U2354 & P2_U2593; 
assign P2_U2664 = P2_U2354 & P2_U2592; 
assign P2_U2665 = P2_U2354 & P2_U2591; 
assign P2_U2674 = P2_U2355 & P2_INSTQUEUE_REG_0__7__SCAN_IN; 
assign P2_U2675 = P2_U2355 & P2_INSTQUEUE_REG_0__6__SCAN_IN; 
assign P2_U2676 = P2_U2355 & P2_INSTQUEUE_REG_0__5__SCAN_IN; 
assign P2_U2677 = P2_U2355 & P2_INSTQUEUE_REG_0__4__SCAN_IN; 
assign P2_U2678 = P2_U2355 & P2_INSTQUEUE_REG_0__3__SCAN_IN; 
assign P2_U2679 = P2_U2355 & P2_INSTQUEUE_REG_0__2__SCAN_IN; 
assign P2_U2680 = P2_U2355 & P2_INSTQUEUE_REG_0__1__SCAN_IN; 
assign P2_U3288 = ~(P2_U2457 & P2_U7859 & P2_U2458); 
assign P2_U3527 = ~(P2_U3283 & P2_U3289); 
assign P2_U3574 = ~(P2_U5571 & P2_U3295 & P2_U3521); 
assign P2_U3868 = P2_U5573 & P2_U5571; 
assign P2_U4193 = P2_U6873 & P2_U6872 & P2_U6871 & P2_U6870; 
assign P2_U4194 = P2_U6877 & P2_U6876 & P2_U6875 & P2_U6874; 
assign P2_U4197 = P2_U6889 & P2_U6888 & P2_U6887 & P2_U6886; 
assign P2_U4198 = P2_U6893 & P2_U6892 & P2_U6891 & P2_U6890; 
assign P2_U4201 = P2_U6905 & P2_U6904 & P2_U6903 & P2_U6902; 
assign P2_U4202 = P2_U6909 & P2_U6908 & P2_U6907 & P2_U6906; 
assign P2_U4205 = P2_U6921 & P2_U6920 & P2_U6919 & P2_U6918; 
assign P2_U4206 = P2_U6925 & P2_U6924 & P2_U6923 & P2_U6922; 
assign P2_U4209 = P2_U6937 & P2_U6936 & P2_U6935 & P2_U6934; 
assign P2_U4210 = P2_U6941 & P2_U6940 & P2_U6939 & P2_U6938; 
assign P2_U4213 = P2_U6953 & P2_U6952 & P2_U6951 & P2_U6950; 
assign P2_U4214 = P2_U6957 & P2_U6956 & P2_U6955 & P2_U6954; 
assign P2_U4217 = P2_U6969 & P2_U6968 & P2_U6967 & P2_U6966; 
assign P2_U4218 = P2_U6973 & P2_U6972 & P2_U6971 & P2_U6970; 
assign P2_U4221 = P2_U6985 & P2_U6984 & P2_U6983 & P2_U6982; 
assign P2_U4222 = P2_U6989 & P2_U6988 & P2_U6987 & P2_U6986; 
assign P2_U4225 = P2_U7001 & P2_U7000 & P2_U6999 & P2_U6998; 
assign P2_U4226 = P2_U7005 & P2_U7004 & P2_U7003 & P2_U7002; 
assign P2_U4229 = P2_U7019 & P2_U7018 & P2_U7017 & P2_U7016; 
assign P2_U4230 = P2_U7023 & P2_U7022 & P2_U7021 & P2_U7020; 
assign P2_U4233 = P2_U7035 & P2_U7034 & P2_U7033 & P2_U7032; 
assign P2_U4234 = P2_U7039 & P2_U7038 & P2_U7037 & P2_U7036; 
assign P2_U4237 = P2_U7051 & P2_U7050 & P2_U7049 & P2_U7048; 
assign P2_U4238 = P2_U7055 & P2_U7054 & P2_U7053 & P2_U7052; 
assign P2_U4241 = P2_U7067 & P2_U7066 & P2_U7065 & P2_U7064; 
assign P2_U4242 = P2_U7071 & P2_U7070 & P2_U7069 & P2_U7068; 
assign P2_U4245 = P2_U7083 & P2_U7082 & P2_U7081 & P2_U7080; 
assign P2_U4246 = P2_U7087 & P2_U7086 & P2_U7085 & P2_U7084; 
assign P2_U4249 = P2_U7099 & P2_U7098 & P2_U7097 & P2_U7096; 
assign P2_U4250 = P2_U7103 & P2_U7102 & P2_U7101 & P2_U7100; 
assign P2_U4253 = P2_U7115 & P2_U7114 & P2_U7113 & P2_U7112; 
assign P2_U4254 = P2_U7119 & P2_U7118 & P2_U7117 & P2_U7116; 
assign P2_U4257 = P2_U7131 & P2_U7130 & P2_U7129 & P2_U7128; 
assign P2_U4258 = P2_U7135 & P2_U7134 & P2_U7133 & P2_U7132; 
assign P2_U4287 = P2_U7212 & P2_U7211 & P2_U7210 & P2_U7209; 
assign P2_U4288 = P2_U7216 & P2_U7215 & P2_U7214 & P2_U7213; 
assign P2_U4295 = P2_U7246 & P2_U7245 & P2_U7244 & P2_U7243; 
assign P2_U4296 = P2_U7250 & P2_U7249 & P2_U7248 & P2_U7247; 
assign P2_U4303 = P2_U7280 & P2_U7279 & P2_U7278 & P2_U7277; 
assign P2_U4304 = P2_U7284 & P2_U7283 & P2_U7282 & P2_U7281; 
assign P2_U4311 = P2_U7314 & P2_U7313 & P2_U7312 & P2_U7311; 
assign P2_U4312 = P2_U7318 & P2_U7317 & P2_U7316 & P2_U7315; 
assign P2_U4319 = P2_U7348 & P2_U7347 & P2_U7346 & P2_U7345; 
assign P2_U4320 = P2_U7352 & P2_U7351 & P2_U7350 & P2_U7349; 
assign P2_U4327 = P2_U7382 & P2_U7381 & P2_U7380 & P2_U7379; 
assign P2_U4328 = P2_U7386 & P2_U7385 & P2_U7384 & P2_U7383; 
assign P2_U4335 = P2_U7416 & P2_U7415 & P2_U7414 & P2_U7413; 
assign P2_U4336 = P2_U7420 & P2_U7419 & P2_U7418 & P2_U7417; 
assign P2_U4341 = P2_U7430 & P2_U3571; 
assign P2_U4390 = P2_U7731 & P2_U3536; 
assign P2_U4391 = P2_U7735 & P2_U3536; 
assign P2_U4412 = ~P2_U3571; 
assign P2_U4417 = ~P2_U3283; 
assign P2_U4419 = ~P2_U3536; 
assign P2_U4427 = ~P2_U3289; 
assign P2_U4429 = ~P2_U3294; 
assign P2_U4460 = ~(P2_U2438 & P2_U3295); 
assign P2_U4476 = ~P2_U3281; 
assign P2_U4597 = ~(P2_U3294 & P2_U3286); 
assign P2_U4601 = ~P2_U3295; 
assign P2_U4886 = ~P2_U3380; 
assign P2_U5001 = ~P2_U3403; 
assign P2_U5115 = ~P2_U3429; 
assign P2_U5229 = ~P2_U3452; 
assign P2_U5344 = ~P2_U3475; 
assign P2_U5459 = ~P2_U3498; 
assign P2_U5574 = ~(P2_U7895 & P2_U3521 & P2_U3255 & P2_U3289); 
assign P2_U5586 = ~(P2_U2617 & P2_U3295 & P2_U3878); 
assign P2_U5587 = ~(P2_U3295 & P2_U3255); 
assign P2_U5590 = ~P2_U3525; 
assign P2_U5591 = ~(P2_U7738 & P2_U3278); 
assign P2_U5596 = ~(P2_U3295 & P2_U7873); 
assign P2_U5600 = ~(P2_U5597 & P2_U3280); 
assign P2_U6845 = ~P2_U2715; 
assign P2_U6846 = ~(P2_U2715 & P2_U3536); 
assign P2_U6848 = ~(P2_U4184 & P2_U2356); 
assign P2_U6858 = ~(P2_U3286 & P2_U3294 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U7008 = ~(P2_U2586 & P2_INSTQUEUE_REG_0__7__SCAN_IN); 
assign P2_U7009 = ~(P2_U2585 & P2_INSTQUEUE_REG_1__7__SCAN_IN); 
assign P2_U7010 = ~(P2_U2584 & P2_INSTQUEUE_REG_2__7__SCAN_IN); 
assign P2_U7011 = ~(P2_U2583 & P2_INSTQUEUE_REG_3__7__SCAN_IN); 
assign P2_U7012 = ~(P2_U2581 & P2_INSTQUEUE_REG_4__7__SCAN_IN); 
assign P2_U7013 = ~(P2_U2580 & P2_INSTQUEUE_REG_5__7__SCAN_IN); 
assign P2_U7014 = ~(P2_U2579 & P2_INSTQUEUE_REG_6__7__SCAN_IN); 
assign P2_U7015 = ~(P2_U2578 & P2_INSTQUEUE_REG_7__7__SCAN_IN); 
assign P2_U7024 = ~(P2_U2586 & P2_INSTQUEUE_REG_0__6__SCAN_IN); 
assign P2_U7025 = ~(P2_U2585 & P2_INSTQUEUE_REG_1__6__SCAN_IN); 
assign P2_U7026 = ~(P2_U2584 & P2_INSTQUEUE_REG_2__6__SCAN_IN); 
assign P2_U7027 = ~(P2_U2583 & P2_INSTQUEUE_REG_3__6__SCAN_IN); 
assign P2_U7028 = ~(P2_U2581 & P2_INSTQUEUE_REG_4__6__SCAN_IN); 
assign P2_U7029 = ~(P2_U2580 & P2_INSTQUEUE_REG_5__6__SCAN_IN); 
assign P2_U7030 = ~(P2_U2579 & P2_INSTQUEUE_REG_6__6__SCAN_IN); 
assign P2_U7031 = ~(P2_U2578 & P2_INSTQUEUE_REG_7__6__SCAN_IN); 
assign P2_U7040 = ~(P2_U2586 & P2_INSTQUEUE_REG_0__5__SCAN_IN); 
assign P2_U7041 = ~(P2_U2585 & P2_INSTQUEUE_REG_1__5__SCAN_IN); 
assign P2_U7042 = ~(P2_U2584 & P2_INSTQUEUE_REG_2__5__SCAN_IN); 
assign P2_U7043 = ~(P2_U2583 & P2_INSTQUEUE_REG_3__5__SCAN_IN); 
assign P2_U7044 = ~(P2_U2581 & P2_INSTQUEUE_REG_4__5__SCAN_IN); 
assign P2_U7045 = ~(P2_U2580 & P2_INSTQUEUE_REG_5__5__SCAN_IN); 
assign P2_U7046 = ~(P2_U2579 & P2_INSTQUEUE_REG_6__5__SCAN_IN); 
assign P2_U7047 = ~(P2_U2578 & P2_INSTQUEUE_REG_7__5__SCAN_IN); 
assign P2_U7056 = ~(P2_U2586 & P2_INSTQUEUE_REG_0__4__SCAN_IN); 
assign P2_U7057 = ~(P2_U2585 & P2_INSTQUEUE_REG_1__4__SCAN_IN); 
assign P2_U7058 = ~(P2_U2584 & P2_INSTQUEUE_REG_2__4__SCAN_IN); 
assign P2_U7059 = ~(P2_U2583 & P2_INSTQUEUE_REG_3__4__SCAN_IN); 
assign P2_U7060 = ~(P2_U2581 & P2_INSTQUEUE_REG_4__4__SCAN_IN); 
assign P2_U7061 = ~(P2_U2580 & P2_INSTQUEUE_REG_5__4__SCAN_IN); 
assign P2_U7062 = ~(P2_U2579 & P2_INSTQUEUE_REG_6__4__SCAN_IN); 
assign P2_U7063 = ~(P2_U2578 & P2_INSTQUEUE_REG_7__4__SCAN_IN); 
assign P2_U7072 = ~(P2_U2586 & P2_INSTQUEUE_REG_0__3__SCAN_IN); 
assign P2_U7073 = ~(P2_U2585 & P2_INSTQUEUE_REG_1__3__SCAN_IN); 
assign P2_U7074 = ~(P2_U2584 & P2_INSTQUEUE_REG_2__3__SCAN_IN); 
assign P2_U7075 = ~(P2_U2583 & P2_INSTQUEUE_REG_3__3__SCAN_IN); 
assign P2_U7076 = ~(P2_U2581 & P2_INSTQUEUE_REG_4__3__SCAN_IN); 
assign P2_U7077 = ~(P2_U2580 & P2_INSTQUEUE_REG_5__3__SCAN_IN); 
assign P2_U7078 = ~(P2_U2579 & P2_INSTQUEUE_REG_6__3__SCAN_IN); 
assign P2_U7079 = ~(P2_U2578 & P2_INSTQUEUE_REG_7__3__SCAN_IN); 
assign P2_U7088 = ~(P2_U2586 & P2_INSTQUEUE_REG_0__2__SCAN_IN); 
assign P2_U7089 = ~(P2_U2585 & P2_INSTQUEUE_REG_1__2__SCAN_IN); 
assign P2_U7090 = ~(P2_U2584 & P2_INSTQUEUE_REG_2__2__SCAN_IN); 
assign P2_U7091 = ~(P2_U2583 & P2_INSTQUEUE_REG_3__2__SCAN_IN); 
assign P2_U7092 = ~(P2_U2581 & P2_INSTQUEUE_REG_4__2__SCAN_IN); 
assign P2_U7093 = ~(P2_U2580 & P2_INSTQUEUE_REG_5__2__SCAN_IN); 
assign P2_U7094 = ~(P2_U2579 & P2_INSTQUEUE_REG_6__2__SCAN_IN); 
assign P2_U7095 = ~(P2_U2578 & P2_INSTQUEUE_REG_7__2__SCAN_IN); 
assign P2_U7104 = ~(P2_U2586 & P2_INSTQUEUE_REG_0__1__SCAN_IN); 
assign P2_U7105 = ~(P2_U2585 & P2_INSTQUEUE_REG_1__1__SCAN_IN); 
assign P2_U7106 = ~(P2_U2584 & P2_INSTQUEUE_REG_2__1__SCAN_IN); 
assign P2_U7107 = ~(P2_U2583 & P2_INSTQUEUE_REG_3__1__SCAN_IN); 
assign P2_U7108 = ~(P2_U2581 & P2_INSTQUEUE_REG_4__1__SCAN_IN); 
assign P2_U7109 = ~(P2_U2580 & P2_INSTQUEUE_REG_5__1__SCAN_IN); 
assign P2_U7110 = ~(P2_U2579 & P2_INSTQUEUE_REG_6__1__SCAN_IN); 
assign P2_U7111 = ~(P2_U2578 & P2_INSTQUEUE_REG_7__1__SCAN_IN); 
assign P2_U7120 = ~(P2_U2586 & P2_INSTQUEUE_REG_0__0__SCAN_IN); 
assign P2_U7121 = ~(P2_U2585 & P2_INSTQUEUE_REG_1__0__SCAN_IN); 
assign P2_U7122 = ~(P2_U2584 & P2_INSTQUEUE_REG_2__0__SCAN_IN); 
assign P2_U7123 = ~(P2_U2583 & P2_INSTQUEUE_REG_3__0__SCAN_IN); 
assign P2_U7124 = ~(P2_U2581 & P2_INSTQUEUE_REG_4__0__SCAN_IN); 
assign P2_U7125 = ~(P2_U2580 & P2_INSTQUEUE_REG_5__0__SCAN_IN); 
assign P2_U7126 = ~(P2_U2579 & P2_INSTQUEUE_REG_6__0__SCAN_IN); 
assign P2_U7127 = ~(P2_U2578 & P2_INSTQUEUE_REG_7__0__SCAN_IN); 
assign P2_U7166 = ~(P2_U2355 & P2_INSTQUEUE_REG_0__0__SCAN_IN); 
assign P2_U7426 = ~(P2_U2439 & P2_U3295); 
assign P2_U7736 = ~(P2_U3295 & P2_U7873 & P2_U3525); 
assign P2_U7744 = ~(P2_U7745 & P2_U3278); 
assign P2_U8117 = ~(P2_U2438 & P2_U7873); 
assign P2_U8348 = ~(P2_U7867 & P2_U3525); 
assign P2_U8359 = ~(P2_R2238_U22 & P2_U3283); 
assign P2_U8367 = ~(P2_R2337_U64 & P2_U3284); 
assign P1_U2353 = P1_U4231 & P1_STATE2_REG_2__SCAN_IN; 
assign P1_U2447 = P1_U3577 & P1_U2452; 
assign P1_U2678 = ~(P1_U7456 & P1_U3284); 
assign P1_U2722 = ~(P1_U4159 & P1_U4192); 
assign P1_U3244 = ~(P1_U3391 & P1_U3394 & P1_U5463); 
assign P1_U3279 = ~(P1_U3559 & P1_U3558); 
assign P1_U3286 = ~(P1_U2389 & P1_U3283); 
assign P1_U3291 = ~(P1_U4190 & P1_U3284); 
assign P1_U3396 = ~(P1_U3741 & P1_U4247); 
assign P1_U3411 = ~(P1_U4190 & P1_U2452); 
assign P1_U3422 = ~(P1_U4210 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U3423 = ~(P1_U4503 & P1_U3391); 
assign P1_U3734 = P1_U4210 & P1_U3257; 
assign P1_U3754 = P1_U5558 & P1_U3257; 
assign P1_U3759 = P1_U4186 & P1_U3284; 
assign P1_U3866 = P1_U2449 & P1_STATE2_REG_0__SCAN_IN; 
assign P1_U3889 = P1_U4494 & P1_U4186; 
assign P1_U3968 = P1_U3287 & P1_STATE2_REG_2__SCAN_IN; 
assign P1_U3972 = P1_U6629 & P1_U6628 & P1_U6627 & P1_U6626; 
assign P1_U3973 = P1_U6633 & P1_U6632 & P1_U6631 & P1_U6630; 
assign P1_U3976 = P1_U6645 & P1_U6644 & P1_U6643 & P1_U6642; 
assign P1_U3977 = P1_U6649 & P1_U6648 & P1_U6647 & P1_U6646; 
assign P1_U3980 = P1_U6661 & P1_U6660 & P1_U6659 & P1_U6658; 
assign P1_U3981 = P1_U6665 & P1_U6664 & P1_U6663 & P1_U6662; 
assign P1_U3984 = P1_U6677 & P1_U6676 & P1_U6675 & P1_U6674; 
assign P1_U3985 = P1_U7613 & P1_U6680 & P1_U6679 & P1_U6678; 
assign P1_U3988 = P1_U6692 & P1_U6691 & P1_U6690 & P1_U6689; 
assign P1_U3989 = P1_U6696 & P1_U6695 & P1_U6694 & P1_U6693; 
assign P1_U3992 = P1_U6708 & P1_U6707 & P1_U6706 & P1_U6705; 
assign P1_U3993 = P1_U6712 & P1_U6711 & P1_U6710 & P1_U6709; 
assign P1_U3996 = P1_U6724 & P1_U6723 & P1_U6722 & P1_U6721; 
assign P1_U3997 = P1_U6728 & P1_U6727 & P1_U6726 & P1_U6725; 
assign P1_U4000 = P1_U6740 & P1_U6739 & P1_U6738 & P1_U6737; 
assign P1_U4001 = P1_U6744 & P1_U6743 & P1_U6742 & P1_U6741; 
assign P1_U4029 = P1_U6895 & P1_U6894 & P1_U6893 & P1_U6892; 
assign P1_U4030 = P1_U6899 & P1_U6898 & P1_U6897 & P1_U6896; 
assign P1_U4033 = P1_U6913 & P1_U6912 & P1_U6911 & P1_U6910; 
assign P1_U4034 = P1_U6917 & P1_U6916 & P1_U6915 & P1_U6914; 
assign P1_U4037 = P1_U6944 & P1_U6943 & P1_U6942 & P1_U6941; 
assign P1_U4038 = P1_U6948 & P1_U6947 & P1_U6946 & P1_U6945; 
assign P1_U4041 = P1_U6961 & P1_U6960 & P1_U6959 & P1_U6958; 
assign P1_U4042 = P1_U6965 & P1_U6964 & P1_U6963 & P1_U6962; 
assign P1_U4045 = P1_U6978 & P1_U6977 & P1_U6976 & P1_U6975; 
assign P1_U4046 = P1_U6982 & P1_U6981 & P1_U6980 & P1_U6979; 
assign P1_U4049 = P1_U6995 & P1_U6994 & P1_U6993 & P1_U6992; 
assign P1_U4050 = P1_U6999 & P1_U6998 & P1_U6997 & P1_U6996; 
assign P1_U4053 = P1_U7010 & P1_U7009 & P1_U7008 & P1_U7007; 
assign P1_U4054 = P1_U7014 & P1_U7013 & P1_U7012 & P1_U7011; 
assign P1_U4057 = P1_U7027 & P1_U7026 & P1_U7025 & P1_U7024; 
assign P1_U4058 = P1_U7031 & P1_U7030 & P1_U7029 & P1_U7028; 
assign P1_U4121 = P1_U7223 & P1_U7222 & P1_U7221 & P1_U7220; 
assign P1_U4122 = P1_U7227 & P1_U7226 & P1_U7225 & P1_U7224; 
assign P1_U4125 = P1_U7240 & P1_U7239 & P1_U7238 & P1_U7237; 
assign P1_U4126 = P1_U7244 & P1_U7243 & P1_U7242 & P1_U7241; 
assign P1_U4129 = P1_U7257 & P1_U7256 & P1_U7255 & P1_U7254; 
assign P1_U4130 = P1_U7261 & P1_U7260 & P1_U7259 & P1_U7258; 
assign P1_U4133 = P1_U7274 & P1_U7273 & P1_U7272 & P1_U7271; 
assign P1_U4134 = P1_U7278 & P1_U7277 & P1_U7276 & P1_U7275; 
assign P1_U4137 = P1_U7289 & P1_U7288 & P1_U7287 & P1_U7286; 
assign P1_U4138 = P1_U7293 & P1_U7292 & P1_U7291 & P1_U7290; 
assign P1_U4141 = P1_U7306 & P1_U7305 & P1_U7304 & P1_U7303; 
assign P1_U4142 = P1_U7310 & P1_U7309 & P1_U7308 & P1_U7307; 
assign P1_U4145 = P1_U7323 & P1_U7322 & P1_U7321 & P1_U7320; 
assign P1_U4146 = P1_U7327 & P1_U7326 & P1_U7325 & P1_U7324; 
assign P1_U4149 = P1_U7340 & P1_U7339 & P1_U7338 & P1_U7337; 
assign P1_U4150 = P1_U7344 & P1_U7343 & P1_U7342 & P1_U7341; 
assign P1_U4153 = P1_U3284 & P1_U3419; 
assign P1_U4188 = ~P1_U3439; 
assign P1_U4189 = ~P1_U3393; 
assign P1_U4191 = ~P1_U3449; 
assign P1_U4199 = ~P1_U3289; 
assign P1_U4206 = ~P1_U3418; 
assign P1_U4208 = ~P1_U3282; 
assign P1_U4234 = ~P1_U3395; 
assign P1_U4236 = ~P1_U3398; 
assign P1_U4249 = ~P1_U3287; 
assign P1_U4250 = ~P1_U3397; 
assign P1_U4253 = ~P1_U3409; 
assign P1_U4254 = ~P1_U3419; 
assign P1_U4500 = ~(P1_U3272 & P1_U3390 & P1_U3287); 
assign P1_U4553 = ~(P1_U4545 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U4670 = ~(P1_U4664 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U4779 = ~P1_U3345; 
assign P1_U4790 = ~(P1_U3345 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U4847 = ~(P1_U4836 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U4894 = ~P1_U3352; 
assign P1_U4905 = ~(P1_U3352 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U4962 = ~(P1_U4951 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U5008 = ~P1_U3362; 
assign P1_U5018 = ~(P1_U3362 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U5075 = ~(P1_U5064 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U5122 = ~P1_U3369; 
assign P1_U5133 = ~(P1_U3369 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U5190 = ~(P1_U5179 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U5237 = ~P1_U3376; 
assign P1_U5248 = ~(P1_U3376 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U5305 = ~(P1_U5294 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U5352 = ~P1_U3383; 
assign P1_U5363 = ~(P1_U3383 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U5420 = ~(P1_U5409 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U5462 = ~(P1_U3391 & P1_U3394 & P1_U4503); 
assign P1_U5465 = ~(P1_U4494 & P1_U3289); 
assign P1_U5467 = ~(P1_U3732 & P1_U2452); 
assign P1_U5471 = ~(P1_U2449 & P1_U7494); 
assign P1_U5472 = ~(P1_U4257 & P1_U4503); 
assign P1_U5489 = ~(P1_U7704 & P1_U7703 & P1_U7494); 
assign P1_U5491 = ~(P1_U4400 & P1_U3394 & P1_U3409); 
assign P1_U5495 = ~(P1_U3395 & P1_U5494); 
assign P1_U5497 = ~(P1_U4257 & P1_U4503); 
assign P1_U5561 = ~(P1_U4235 & P1_U4503 & P1_U4192); 
assign P1_U5959 = ~(U210 & P1_U3282); 
assign P1_U6746 = ~(P1_U3412 & P1_U6745); 
assign P1_U6762 = ~(P1_R2337_U66 & P1_U2352); 
assign P1_U6900 = ~(P1_U2554 & P1_INSTQUEUE_REG_7__1__SCAN_IN); 
assign P1_U6901 = ~(P1_U2553 & P1_INSTQUEUE_REG_6__1__SCAN_IN); 
assign P1_U6902 = ~(P1_U2552 & P1_INSTQUEUE_REG_5__1__SCAN_IN); 
assign P1_U6903 = ~(P1_U2551 & P1_INSTQUEUE_REG_4__1__SCAN_IN); 
assign P1_U6904 = ~(P1_U2549 & P1_INSTQUEUE_REG_3__1__SCAN_IN); 
assign P1_U6905 = ~(P1_U2548 & P1_INSTQUEUE_REG_2__1__SCAN_IN); 
assign P1_U6906 = ~(P1_U2547 & P1_INSTQUEUE_REG_1__1__SCAN_IN); 
assign P1_U6907 = ~(P1_U2546 & P1_INSTQUEUE_REG_0__1__SCAN_IN); 
assign P1_U6909 = ~(P1_U3405 & P1_U3418); 
assign P1_U6918 = ~(P1_U2554 & P1_INSTQUEUE_REG_7__0__SCAN_IN); 
assign P1_U6919 = ~(P1_U2553 & P1_INSTQUEUE_REG_6__0__SCAN_IN); 
assign P1_U6920 = ~(P1_U2552 & P1_INSTQUEUE_REG_5__0__SCAN_IN); 
assign P1_U6921 = ~(P1_U2551 & P1_INSTQUEUE_REG_4__0__SCAN_IN); 
assign P1_U6922 = ~(P1_U2549 & P1_INSTQUEUE_REG_3__0__SCAN_IN); 
assign P1_U6923 = ~(P1_U2548 & P1_INSTQUEUE_REG_2__0__SCAN_IN); 
assign P1_U6924 = ~(P1_U2547 & P1_INSTQUEUE_REG_1__0__SCAN_IN); 
assign P1_U6925 = ~(P1_U2546 & P1_INSTQUEUE_REG_0__0__SCAN_IN); 
assign P1_U6949 = ~(P1_U2554 & P1_INSTQUEUE_REG_7__7__SCAN_IN); 
assign P1_U6950 = ~(P1_U2553 & P1_INSTQUEUE_REG_6__7__SCAN_IN); 
assign P1_U6951 = ~(P1_U2552 & P1_INSTQUEUE_REG_5__7__SCAN_IN); 
assign P1_U6952 = ~(P1_U2551 & P1_INSTQUEUE_REG_4__7__SCAN_IN); 
assign P1_U6953 = ~(P1_U2549 & P1_INSTQUEUE_REG_3__7__SCAN_IN); 
assign P1_U6954 = ~(P1_U2548 & P1_INSTQUEUE_REG_2__7__SCAN_IN); 
assign P1_U6955 = ~(P1_U2547 & P1_INSTQUEUE_REG_1__7__SCAN_IN); 
assign P1_U6956 = ~(P1_U2546 & P1_INSTQUEUE_REG_0__7__SCAN_IN); 
assign P1_U6966 = ~(P1_U2554 & P1_INSTQUEUE_REG_7__6__SCAN_IN); 
assign P1_U6967 = ~(P1_U2553 & P1_INSTQUEUE_REG_6__6__SCAN_IN); 
assign P1_U6968 = ~(P1_U2552 & P1_INSTQUEUE_REG_5__6__SCAN_IN); 
assign P1_U6969 = ~(P1_U2551 & P1_INSTQUEUE_REG_4__6__SCAN_IN); 
assign P1_U6970 = ~(P1_U2549 & P1_INSTQUEUE_REG_3__6__SCAN_IN); 
assign P1_U6971 = ~(P1_U2548 & P1_INSTQUEUE_REG_2__6__SCAN_IN); 
assign P1_U6972 = ~(P1_U2547 & P1_INSTQUEUE_REG_1__6__SCAN_IN); 
assign P1_U6973 = ~(P1_U2546 & P1_INSTQUEUE_REG_0__6__SCAN_IN); 
assign P1_U6983 = ~(P1_U2554 & P1_INSTQUEUE_REG_7__5__SCAN_IN); 
assign P1_U6984 = ~(P1_U2553 & P1_INSTQUEUE_REG_6__5__SCAN_IN); 
assign P1_U6985 = ~(P1_U2552 & P1_INSTQUEUE_REG_5__5__SCAN_IN); 
assign P1_U6986 = ~(P1_U2551 & P1_INSTQUEUE_REG_4__5__SCAN_IN); 
assign P1_U6987 = ~(P1_U2549 & P1_INSTQUEUE_REG_3__5__SCAN_IN); 
assign P1_U6988 = ~(P1_U2548 & P1_INSTQUEUE_REG_2__5__SCAN_IN); 
assign P1_U6989 = ~(P1_U2547 & P1_INSTQUEUE_REG_1__5__SCAN_IN); 
assign P1_U6990 = ~(P1_U2546 & P1_INSTQUEUE_REG_0__5__SCAN_IN); 
assign P1_U7000 = ~(P1_U2554 & P1_INSTQUEUE_REG_7__4__SCAN_IN); 
assign P1_U7001 = ~(P1_U2553 & P1_INSTQUEUE_REG_6__4__SCAN_IN); 
assign P1_U7002 = ~(P1_U2552 & P1_INSTQUEUE_REG_5__4__SCAN_IN); 
assign P1_U7003 = ~(P1_U2551 & P1_INSTQUEUE_REG_4__4__SCAN_IN); 
assign P1_U7004 = ~(P1_U2549 & P1_INSTQUEUE_REG_3__4__SCAN_IN); 
assign P1_U7005 = ~(P1_U2548 & P1_INSTQUEUE_REG_2__4__SCAN_IN); 
assign P1_U7006 = ~(P1_U2547 & P1_INSTQUEUE_REG_1__4__SCAN_IN); 
assign P1_U7015 = ~(P1_U2554 & P1_INSTQUEUE_REG_7__3__SCAN_IN); 
assign P1_U7016 = ~(P1_U2553 & P1_INSTQUEUE_REG_6__3__SCAN_IN); 
assign P1_U7017 = ~(P1_U2552 & P1_INSTQUEUE_REG_5__3__SCAN_IN); 
assign P1_U7018 = ~(P1_U2551 & P1_INSTQUEUE_REG_4__3__SCAN_IN); 
assign P1_U7019 = ~(P1_U2549 & P1_INSTQUEUE_REG_3__3__SCAN_IN); 
assign P1_U7020 = ~(P1_U2548 & P1_INSTQUEUE_REG_2__3__SCAN_IN); 
assign P1_U7021 = ~(P1_U2547 & P1_INSTQUEUE_REG_1__3__SCAN_IN); 
assign P1_U7022 = ~(P1_U2546 & P1_INSTQUEUE_REG_0__3__SCAN_IN); 
assign P1_U7032 = ~(P1_U2554 & P1_INSTQUEUE_REG_7__2__SCAN_IN); 
assign P1_U7033 = ~(P1_U2553 & P1_INSTQUEUE_REG_6__2__SCAN_IN); 
assign P1_U7034 = ~(P1_U2552 & P1_INSTQUEUE_REG_5__2__SCAN_IN); 
assign P1_U7035 = ~(P1_U2551 & P1_INSTQUEUE_REG_4__2__SCAN_IN); 
assign P1_U7036 = ~(P1_U2549 & P1_INSTQUEUE_REG_3__2__SCAN_IN); 
assign P1_U7037 = ~(P1_U2548 & P1_INSTQUEUE_REG_2__2__SCAN_IN); 
assign P1_U7038 = ~(P1_U2547 & P1_INSTQUEUE_REG_1__2__SCAN_IN); 
assign P1_U7039 = ~(P1_U2546 & P1_INSTQUEUE_REG_0__2__SCAN_IN); 
assign P1_U7048 = ~(P1_U4192 & P1_INSTQUEUE_REG_0__7__SCAN_IN); 
assign P1_U7050 = ~(P1_U4192 & P1_INSTQUEUE_REG_0__6__SCAN_IN); 
assign P1_U7052 = ~(P1_U4192 & P1_INSTQUEUE_REG_0__5__SCAN_IN); 
assign P1_U7055 = ~(P1_U4192 & P1_INSTQUEUE_REG_0__3__SCAN_IN); 
assign P1_U7057 = ~(P1_U4192 & P1_INSTQUEUE_REG_0__2__SCAN_IN); 
assign P1_U7059 = ~(P1_U4192 & P1_INSTQUEUE_REG_0__1__SCAN_IN); 
assign P1_U7062 = ~(P1_U4192 & P1_INSTQUEUE_REG_0__0__SCAN_IN); 
assign P1_U7082 = ~(P1_U4066 & P1_U4065 & P1_U4064 & P1_U4063); 
assign P1_U7086 = ~(P1_U4503 & P1_U3278); 
assign P1_U7088 = ~(P1_U4400 & P1_U4503 & P1_U4154 & P1_U3394); 
assign P1_U7114 = ~(P1_U4082 & P1_U4081 & P1_U4080 & P1_U4079); 
assign P1_U7131 = ~(P1_U4086 & P1_U4085 & P1_U4084 & P1_U4083); 
assign P1_U7163 = ~(P1_U4095 & P1_U4094 & P1_U4093 & P1_U4092); 
assign P1_U7180 = ~(P1_U4099 & P1_U4098 & P1_U4097 & P1_U4096); 
assign P1_U7197 = ~(P1_U4103 & P1_U4102 & P1_U4101 & P1_U4100); 
assign P1_U7214 = ~(P1_U4107 & P1_U4106 & P1_U4105 & P1_U4104); 
assign P1_U7228 = ~(P1_U2592 & P1_INSTQUEUE_REG_0__7__SCAN_IN); 
assign P1_U7229 = ~(P1_U2591 & P1_INSTQUEUE_REG_1__7__SCAN_IN); 
assign P1_U7230 = ~(P1_U2590 & P1_INSTQUEUE_REG_2__7__SCAN_IN); 
assign P1_U7231 = ~(P1_U2589 & P1_INSTQUEUE_REG_3__7__SCAN_IN); 
assign P1_U7232 = ~(P1_U2587 & P1_INSTQUEUE_REG_4__7__SCAN_IN); 
assign P1_U7233 = ~(P1_U2586 & P1_INSTQUEUE_REG_5__7__SCAN_IN); 
assign P1_U7234 = ~(P1_U2585 & P1_INSTQUEUE_REG_6__7__SCAN_IN); 
assign P1_U7235 = ~(P1_U2584 & P1_INSTQUEUE_REG_7__7__SCAN_IN); 
assign P1_U7245 = ~(P1_U2592 & P1_INSTQUEUE_REG_0__6__SCAN_IN); 
assign P1_U7246 = ~(P1_U2591 & P1_INSTQUEUE_REG_1__6__SCAN_IN); 
assign P1_U7247 = ~(P1_U2590 & P1_INSTQUEUE_REG_2__6__SCAN_IN); 
assign P1_U7248 = ~(P1_U2589 & P1_INSTQUEUE_REG_3__6__SCAN_IN); 
assign P1_U7249 = ~(P1_U2587 & P1_INSTQUEUE_REG_4__6__SCAN_IN); 
assign P1_U7250 = ~(P1_U2586 & P1_INSTQUEUE_REG_5__6__SCAN_IN); 
assign P1_U7251 = ~(P1_U2585 & P1_INSTQUEUE_REG_6__6__SCAN_IN); 
assign P1_U7252 = ~(P1_U2584 & P1_INSTQUEUE_REG_7__6__SCAN_IN); 
assign P1_U7262 = ~(P1_U2592 & P1_INSTQUEUE_REG_0__5__SCAN_IN); 
assign P1_U7263 = ~(P1_U2591 & P1_INSTQUEUE_REG_1__5__SCAN_IN); 
assign P1_U7264 = ~(P1_U2590 & P1_INSTQUEUE_REG_2__5__SCAN_IN); 
assign P1_U7265 = ~(P1_U2589 & P1_INSTQUEUE_REG_3__5__SCAN_IN); 
assign P1_U7266 = ~(P1_U2587 & P1_INSTQUEUE_REG_4__5__SCAN_IN); 
assign P1_U7267 = ~(P1_U2586 & P1_INSTQUEUE_REG_5__5__SCAN_IN); 
assign P1_U7268 = ~(P1_U2585 & P1_INSTQUEUE_REG_6__5__SCAN_IN); 
assign P1_U7269 = ~(P1_U2584 & P1_INSTQUEUE_REG_7__5__SCAN_IN); 
assign P1_U7279 = ~(P1_U2591 & P1_INSTQUEUE_REG_1__4__SCAN_IN); 
assign P1_U7280 = ~(P1_U2590 & P1_INSTQUEUE_REG_2__4__SCAN_IN); 
assign P1_U7281 = ~(P1_U2589 & P1_INSTQUEUE_REG_3__4__SCAN_IN); 
assign P1_U7282 = ~(P1_U2587 & P1_INSTQUEUE_REG_4__4__SCAN_IN); 
assign P1_U7283 = ~(P1_U2586 & P1_INSTQUEUE_REG_5__4__SCAN_IN); 
assign P1_U7284 = ~(P1_U2585 & P1_INSTQUEUE_REG_6__4__SCAN_IN); 
assign P1_U7285 = ~(P1_U2584 & P1_INSTQUEUE_REG_7__4__SCAN_IN); 
assign P1_U7294 = ~(P1_U2592 & P1_INSTQUEUE_REG_0__3__SCAN_IN); 
assign P1_U7295 = ~(P1_U2591 & P1_INSTQUEUE_REG_1__3__SCAN_IN); 
assign P1_U7296 = ~(P1_U2590 & P1_INSTQUEUE_REG_2__3__SCAN_IN); 
assign P1_U7297 = ~(P1_U2589 & P1_INSTQUEUE_REG_3__3__SCAN_IN); 
assign P1_U7298 = ~(P1_U2587 & P1_INSTQUEUE_REG_4__3__SCAN_IN); 
assign P1_U7299 = ~(P1_U2586 & P1_INSTQUEUE_REG_5__3__SCAN_IN); 
assign P1_U7300 = ~(P1_U2585 & P1_INSTQUEUE_REG_6__3__SCAN_IN); 
assign P1_U7301 = ~(P1_U2584 & P1_INSTQUEUE_REG_7__3__SCAN_IN); 
assign P1_U7311 = ~(P1_U2592 & P1_INSTQUEUE_REG_0__2__SCAN_IN); 
assign P1_U7312 = ~(P1_U2591 & P1_INSTQUEUE_REG_1__2__SCAN_IN); 
assign P1_U7313 = ~(P1_U2590 & P1_INSTQUEUE_REG_2__2__SCAN_IN); 
assign P1_U7314 = ~(P1_U2589 & P1_INSTQUEUE_REG_3__2__SCAN_IN); 
assign P1_U7315 = ~(P1_U2587 & P1_INSTQUEUE_REG_4__2__SCAN_IN); 
assign P1_U7316 = ~(P1_U2586 & P1_INSTQUEUE_REG_5__2__SCAN_IN); 
assign P1_U7317 = ~(P1_U2585 & P1_INSTQUEUE_REG_6__2__SCAN_IN); 
assign P1_U7318 = ~(P1_U2584 & P1_INSTQUEUE_REG_7__2__SCAN_IN); 
assign P1_U7328 = ~(P1_U2592 & P1_INSTQUEUE_REG_0__1__SCAN_IN); 
assign P1_U7329 = ~(P1_U2591 & P1_INSTQUEUE_REG_1__1__SCAN_IN); 
assign P1_U7330 = ~(P1_U2590 & P1_INSTQUEUE_REG_2__1__SCAN_IN); 
assign P1_U7331 = ~(P1_U2589 & P1_INSTQUEUE_REG_3__1__SCAN_IN); 
assign P1_U7332 = ~(P1_U2587 & P1_INSTQUEUE_REG_4__1__SCAN_IN); 
assign P1_U7333 = ~(P1_U2586 & P1_INSTQUEUE_REG_5__1__SCAN_IN); 
assign P1_U7334 = ~(P1_U2585 & P1_INSTQUEUE_REG_6__1__SCAN_IN); 
assign P1_U7335 = ~(P1_U2584 & P1_INSTQUEUE_REG_7__1__SCAN_IN); 
assign P1_U7345 = ~(P1_U2592 & P1_INSTQUEUE_REG_0__0__SCAN_IN); 
assign P1_U7346 = ~(P1_U2591 & P1_INSTQUEUE_REG_1__0__SCAN_IN); 
assign P1_U7347 = ~(P1_U2590 & P1_INSTQUEUE_REG_2__0__SCAN_IN); 
assign P1_U7348 = ~(P1_U2589 & P1_INSTQUEUE_REG_3__0__SCAN_IN); 
assign P1_U7349 = ~(P1_U2587 & P1_INSTQUEUE_REG_4__0__SCAN_IN); 
assign P1_U7350 = ~(P1_U2586 & P1_INSTQUEUE_REG_5__0__SCAN_IN); 
assign P1_U7351 = ~(P1_U2585 & P1_INSTQUEUE_REG_6__0__SCAN_IN); 
assign P1_U7352 = ~(P1_U2584 & P1_INSTQUEUE_REG_7__0__SCAN_IN); 
assign P1_U7358 = ~(P1_U4190 & P1_U2452); 
assign P1_U7362 = ~(P1_U2451 & P1_U4210); 
assign P1_U7373 = ~(P1_SUB_450_U22 & P1_U2354); 
assign P1_U7375 = ~(P1_SUB_450_U7 & P1_U2354); 
assign P1_U7385 = ~(P1_R2238_U22 & P1_U4192); 
assign P1_U7387 = ~(P1_U2451 & P1_U3284); 
assign P1_U7388 = ~(P1_R2238_U7 & P1_U4192); 
assign P1_U7390 = ~(P1_U3393 & P1_U3290); 
assign P1_U7391 = ~(P1_U3284 & P1_U3449); 
assign P1_U7490 = ~(P1_U7785 & P1_U7784 & P1_U4072); 
assign P1_U7614 = ~(P1_U2546 & P1_INSTQUEUE_REG_0__4__SCAN_IN); 
assign P1_U7616 = ~(P1_U4192 & P1_INSTQUEUE_REG_0__4__SCAN_IN); 
assign P1_U7618 = ~(P1_U4091 & P1_U4089 & P1_U4088 & P1_U4087); 
assign P1_U7619 = ~(P1_U2592 & P1_INSTQUEUE_REG_0__4__SCAN_IN); 
assign P1_U7627 = ~(P1_U5487 & P1_U4171); 
assign P1_U7628 = ~(P1_U3283 & P1_U3289); 
assign P1_U7631 = ~(P1_U5487 & P1_U4171); 
assign P3_ADD_526_U22 = ~(P3_ADD_526_U85 & P3_ADD_526_U120); 
assign P3_ADD_526_U110 = ~(P3_ADD_526_U120 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_526_U141 = ~(P3_ADD_526_U120 & P3_ADD_526_U18); 
assign P3_ADD_526_U144 = ~(P3_ADD_526_U125 & P3_ADD_526_U14); 
assign P3_ADD_552_U22 = ~(P3_ADD_552_U85 & P3_ADD_552_U120); 
assign P3_ADD_552_U110 = ~(P3_ADD_552_U120 & P3_EBX_REG_9__SCAN_IN); 
assign P3_ADD_552_U141 = ~(P3_ADD_552_U120 & P3_ADD_552_U18); 
assign P3_ADD_552_U144 = ~(P3_ADD_552_U125 & P3_ADD_552_U14); 
assign P3_ADD_546_U22 = ~(P3_ADD_546_U85 & P3_ADD_546_U120); 
assign P3_ADD_546_U110 = ~(P3_ADD_546_U120 & P3_EAX_REG_9__SCAN_IN); 
assign P3_ADD_546_U141 = ~(P3_ADD_546_U120 & P3_ADD_546_U18); 
assign P3_ADD_546_U144 = ~(P3_ADD_546_U125 & P3_ADD_546_U14); 
assign P3_ADD_476_U14 = ~(P3_ADD_476_U97 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_476_U130 = ~(P3_ADD_476_U97 & P3_ADD_476_U13); 
assign P3_ADD_531_U15 = ~(P3_ADD_531_U101 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_531_U137 = ~(P3_ADD_531_U101 & P3_ADD_531_U14); 
assign P3_SUB_320_U18 = P3_SUB_320_U92 & P3_SUB_320_U22; 
assign P3_SUB_320_U56 = ~P3_ADD_318_U66; 
assign P3_SUB_320_U84 = ~P3_SUB_320_U22; 
assign P3_SUB_320_U132 = ~(P3_ADD_318_U66 & P3_SUB_320_U22); 
assign P3_ADD_318_U14 = ~(P3_ADD_318_U97 & P3_PHYADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_318_U130 = ~(P3_ADD_318_U97 & P3_ADD_318_U13); 
assign P3_SUB_370_U21 = ~(P3_SUB_370_U61 & P3_SUB_370_U60); 
assign P3_SUB_370_U38 = ~P3_SUB_370_U27; 
assign P3_SUB_370_U40 = ~(P3_SUB_370_U39 & P3_SUB_370_U27); 
assign P3_SUB_370_U56 = ~(P3_SUB_370_U24 & P3_SUB_370_U27); 
assign P3_ADD_315_U14 = ~(P3_ADD_315_U94 & P3_PHYADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_315_U124 = ~(P3_ADD_315_U94 & P3_ADD_315_U13); 
assign P3_SUB_589_U6 = ~P3_U3301; 
assign P3_ADD_467_U14 = ~(P3_ADD_467_U97 & P3_REIP_REG_6__SCAN_IN); 
assign P3_ADD_467_U130 = ~(P3_ADD_467_U97 & P3_ADD_467_U13); 
assign P3_ADD_430_U14 = ~(P3_ADD_430_U97 & P3_REIP_REG_6__SCAN_IN); 
assign P3_ADD_430_U130 = ~(P3_ADD_430_U97 & P3_ADD_430_U13); 
assign P3_ADD_380_U15 = ~(P3_ADD_380_U101 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_380_U137 = ~(P3_ADD_380_U101 & P3_ADD_380_U14); 
assign P3_ADD_344_U15 = ~(P3_ADD_344_U101 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_344_U137 = ~(P3_ADD_344_U101 & P3_ADD_344_U14); 
assign P3_ADD_339_U14 = ~(P3_ADD_339_U97 & P3_PHYADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_339_U130 = ~(P3_ADD_339_U97 & P3_ADD_339_U13); 
assign P3_ADD_541_U14 = ~(P3_ADD_541_U97 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_541_U130 = ~(P3_ADD_541_U97 & P3_ADD_541_U13); 
assign P3_SUB_355_U21 = ~(P3_SUB_355_U61 & P3_SUB_355_U60); 
assign P3_SUB_355_U38 = ~P3_SUB_355_U27; 
assign P3_SUB_355_U40 = ~(P3_SUB_355_U39 & P3_SUB_355_U27); 
assign P3_SUB_355_U56 = ~(P3_SUB_355_U24 & P3_SUB_355_U27); 
assign P3_SUB_450_U18 = ~(P3_SUB_450_U58 & P3_SUB_450_U57); 
assign P3_SUB_450_U36 = ~P3_SUB_450_U24; 
assign P3_SUB_450_U38 = ~(P3_SUB_450_U37 & P3_SUB_450_U24); 
assign P3_SUB_450_U53 = ~(P3_SUB_450_U21 & P3_SUB_450_U24); 
assign P3_SUB_485_U18 = ~(P3_SUB_485_U58 & P3_SUB_485_U57); 
assign P3_SUB_485_U36 = ~P3_SUB_485_U24; 
assign P3_SUB_485_U38 = ~(P3_SUB_485_U37 & P3_SUB_485_U24); 
assign P3_SUB_485_U53 = ~(P3_SUB_485_U21 & P3_SUB_485_U24); 
assign P3_ADD_515_U14 = ~(P3_ADD_515_U97 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_515_U130 = ~(P3_ADD_515_U97 & P3_ADD_515_U13); 
assign P3_ADD_394_U14 = ~(P3_ADD_394_U100 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_394_U134 = ~(P3_ADD_394_U100 & P3_ADD_394_U13); 
assign P3_SUB_414_U20 = P3_SUB_414_U88 & P3_SUB_414_U24; 
assign P3_SUB_414_U28 = ~(P3_SUB_414_U52 & P3_SUB_414_U49 & P3_SUB_414_U86); 
assign P3_SUB_414_U125 = ~(P3_SUB_414_U86 & P3_SUB_414_U52); 
assign P3_SUB_414_U129 = ~(P3_SUB_414_U86 & P3_SUB_414_U52); 
assign P3_ADD_441_U14 = ~(P3_ADD_441_U97 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_441_U130 = ~(P3_ADD_441_U97 & P3_ADD_441_U13); 
assign P3_ADD_349_U15 = ~(P3_ADD_349_U101 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_349_U137 = ~(P3_ADD_349_U101 & P3_ADD_349_U14); 
assign P3_ADD_405_U14 = ~(P3_ADD_405_U100 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_405_U134 = ~(P3_ADD_405_U100 & P3_ADD_405_U13); 
assign P3_ADD_553_U15 = ~(P3_ADD_553_U101 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_553_U137 = ~(P3_ADD_553_U101 & P3_ADD_553_U14); 
assign P3_ADD_558_U15 = ~(P3_ADD_558_U101 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_558_U137 = ~(P3_ADD_558_U101 & P3_ADD_558_U14); 
assign P3_ADD_385_U15 = ~(P3_ADD_385_U101 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_385_U137 = ~(P3_ADD_385_U101 & P3_ADD_385_U14); 
assign P3_ADD_547_U15 = ~(P3_ADD_547_U101 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_547_U137 = ~(P3_ADD_547_U101 & P3_ADD_547_U14); 
assign P3_SUB_412_U18 = ~(P3_SUB_412_U58 & P3_SUB_412_U57); 
assign P3_SUB_412_U36 = ~P3_SUB_412_U24; 
assign P3_SUB_412_U38 = ~(P3_SUB_412_U37 & P3_SUB_412_U24); 
assign P3_SUB_412_U53 = ~(P3_SUB_412_U21 & P3_SUB_412_U24); 
assign P3_SUB_504_U18 = ~(P3_SUB_504_U58 & P3_SUB_504_U57); 
assign P3_SUB_504_U36 = ~P3_SUB_504_U24; 
assign P3_SUB_504_U38 = ~(P3_SUB_504_U37 & P3_SUB_504_U24); 
assign P3_SUB_504_U53 = ~(P3_SUB_504_U21 & P3_SUB_504_U24); 
assign P3_SUB_401_U21 = ~(P3_SUB_401_U61 & P3_SUB_401_U60); 
assign P3_SUB_401_U38 = ~P3_SUB_401_U27; 
assign P3_SUB_401_U40 = ~(P3_SUB_401_U39 & P3_SUB_401_U27); 
assign P3_SUB_401_U56 = ~(P3_SUB_401_U24 & P3_SUB_401_U27); 
assign P3_SUB_390_U21 = ~(P3_SUB_390_U61 & P3_SUB_390_U60); 
assign P3_SUB_390_U38 = ~P3_SUB_390_U27; 
assign P3_SUB_390_U40 = ~(P3_SUB_390_U39 & P3_SUB_390_U27); 
assign P3_SUB_390_U56 = ~(P3_SUB_390_U24 & P3_SUB_390_U27); 
assign P3_ADD_494_U14 = ~(P3_ADD_494_U97 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_494_U130 = ~(P3_ADD_494_U97 & P3_ADD_494_U13); 
assign P3_ADD_536_U14 = ~(P3_ADD_536_U97 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_536_U130 = ~(P3_ADD_536_U97 & P3_ADD_536_U13); 
assign P2_ADD_402_1132_U5 = ~P2_U2591; 
assign P2_ADD_402_1132_U7 = ~P2_U2592; 
assign P2_ADD_402_1132_U9 = ~P2_U2593; 
assign P2_ADD_402_1132_U11 = ~P2_U2594; 
assign P2_ADD_402_1132_U13 = ~P2_U2595; 
assign P2_ADD_402_1132_U15 = ~P2_U2596; 
assign P2_ADD_402_1132_U17 = ~P2_U2597; 
assign P2_ADD_402_1132_U26 = ~P2_U2598; 
assign P2_R2027_U15 = ~(P2_R2027_U101 & P2_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P2_R2027_U137 = ~(P2_R2027_U101 & P2_R2027_U14); 
assign P2_R2337_U15 = ~(P2_R2337_U98 & P2_PHYADDRPOINTER_REG_7__SCAN_IN); 
assign P2_R2337_U128 = ~(P2_R2337_U98 & P2_R2337_U14); 
assign P2_R2147_U10 = ~P2_U2752; 
assign P2_R2147_U15 = ~(P2_U2752 & P2_R2147_U11); 
assign P2_R2219_U9 = ~P2_U4428; 
assign P2_R2238_U21 = ~(P2_R2238_U61 & P2_R2238_U60); 
assign P2_R2238_U38 = ~P2_R2238_U27; 
assign P2_R2238_U40 = ~(P2_R2238_U39 & P2_R2238_U27); 
assign P2_R2238_U56 = ~(P2_R2238_U24 & P2_R2238_U27); 
assign P2_R1957_U56 = ~P2_U3657; 
assign P2_R1957_U59 = P2_R1957_U135 & P2_R1957_U134; 
assign P2_R1957_U84 = ~P2_R1957_U22; 
assign P2_R1957_U92 = ~(P2_U3658 & P2_R1957_U91); 
assign P2_R1957_U132 = ~(P2_U3657 & P2_R1957_U22); 
assign P2_SUB_450_U19 = ~(P2_SUB_450_U58 & P2_SUB_450_U57); 
assign P2_SUB_450_U36 = ~P2_SUB_450_U25; 
assign P2_SUB_450_U38 = ~(P2_SUB_450_U37 & P2_SUB_450_U25); 
assign P2_SUB_450_U53 = ~(P2_SUB_450_U22 & P2_SUB_450_U25); 
assign P2_ADD_394_U14 = ~(P2_ADD_394_U100 & P2_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P2_ADD_394_U128 = ~(P2_ADD_394_U100 & P2_ADD_394_U12); 
assign P1_R2027_U22 = ~(P1_R2027_U85 & P1_R2027_U120); 
assign P1_R2027_U110 = ~(P1_R2027_U120 & P1_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P1_R2027_U141 = ~(P1_R2027_U120 & P1_R2027_U18); 
assign P1_R2027_U144 = ~(P1_R2027_U125 & P1_R2027_U14); 
assign P1_R2099_U4 = ~P1_U4190; 
assign P1_R2337_U14 = ~(P1_R2337_U97 & P1_PHYADDRPOINTER_REG_6__SCAN_IN); 
assign P1_R2337_U130 = ~(P1_R2337_U97 & P1_R2337_U13); 
assign P1_R2096_U14 = ~(P1_R2096_U97 & P1_REIP_REG_6__SCAN_IN); 
assign P1_R2096_U130 = ~(P1_R2096_U97 & P1_R2096_U13); 
assign P1_R2238_U21 = ~(P1_R2238_U61 & P1_R2238_U60); 
assign P1_R2238_U38 = ~P1_R2238_U27; 
assign P1_R2238_U40 = ~(P1_R2238_U39 & P1_R2238_U27); 
assign P1_R2238_U56 = ~(P1_R2238_U24 & P1_R2238_U27); 
assign P1_SUB_450_U21 = ~(P1_SUB_450_U61 & P1_SUB_450_U60); 
assign P1_SUB_450_U38 = ~P1_SUB_450_U27; 
assign P1_SUB_450_U40 = ~(P1_SUB_450_U39 & P1_SUB_450_U27); 
assign P1_SUB_450_U56 = ~(P1_SUB_450_U24 & P1_SUB_450_U27); 
assign P1_ADD_405_U14 = ~(P1_ADD_405_U100 & P1_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P1_ADD_405_U128 = ~(P1_ADD_405_U100 & P1_ADD_405_U12); 
assign P1_ADD_515_U14 = ~(P1_ADD_515_U97 & P1_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P1_ADD_515_U124 = ~(P1_ADD_515_U97 & P1_ADD_515_U12); 
assign P3_U2412 = P3_U3218 & P3_U3107 & P3_U4539; 
assign P3_U2456 = P3_U4556 & P3_U4607; 
assign P3_U2461 = P3_U4573 & P3_U4522; 
assign P3_U2463 = P3_U4590 & P3_U4607; 
assign P3_U2490 = P3_U3156 & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN; 
assign P3_U3112 = ~(P3_U4505 & P3_U3108); 
assign P3_U3113 = ~(P3_U4607 & P3_U3110); 
assign P3_U3114 = ~(P3_U4488 & P3_U4505); 
assign P3_U3118 = ~(P3_U4488 & P3_U3104); 
assign P3_U3142 = ~(P3_U4331 & P3_U4655); 
assign P3_U3143 = ~(P3_U3156 & P3_U3128); 
assign P3_U3185 = ~(P3_U3180 & P3_U4331); 
assign P3_U3189 = ~(P3_U3186 & P3_U5128); 
assign P3_U3193 = ~(P3_U3190 & P3_U5180); 
assign P3_U3198 = ~(P3_U3196 & P3_U5282); 
assign P3_U3201 = ~(P3_U3199 & P3_U5333); 
assign P3_U3204 = ~(P3_U3202 & P3_U5384); 
assign P3_U3208 = ~(P3_U4539 & P3_U3102); 
assign P3_U3216 = ~(P3_U4590 & P3_U3074); 
assign P3_U3236 = ~(P3_U3101 & P3_U2630 & P3_U4505); 
assign P3_U3271 = ~(P3_U7967 & P3_U7966); 
assign P3_U3354 = P3_U4556 & P3_U3218; 
assign P3_U3359 = P3_U4539 & P3_U2630; 
assign P3_U3654 = P3_U4522 & P3_U3104; 
assign P3_U3660 = P3_U4556 & P3_U4539; 
assign P3_U3662 = P3_U4590 & P3_U3101; 
assign P3_U3663 = P3_U4556 & P3_U3101; 
assign P3_U3953 = P3_U4505 & P3_STATE2_REG_0__SCAN_IN; 
assign P3_U4154 = P3_U7398 & P3_U7397 & P3_U7396 & P3_U7395; 
assign P3_U4155 = P3_U7402 & P3_U7401 & P3_U7400 & P3_U7399; 
assign P3_U4158 = P3_U7414 & P3_U7413 & P3_U7412 & P3_U7411; 
assign P3_U4159 = P3_U7418 & P3_U7417 & P3_U7416 & P3_U7415; 
assign P3_U4162 = P3_U7430 & P3_U7429 & P3_U7428 & P3_U7427; 
assign P3_U4163 = P3_U7434 & P3_U7433 & P3_U7432 & P3_U7431; 
assign P3_U4166 = P3_U7446 & P3_U7445 & P3_U7444 & P3_U7443; 
assign P3_U4167 = P3_U7450 & P3_U7449 & P3_U7448 & P3_U7447; 
assign P3_U4170 = P3_U7462 & P3_U7461 & P3_U7460 & P3_U7459; 
assign P3_U4171 = P3_U7466 & P3_U7465 & P3_U7464 & P3_U7463; 
assign P3_U4174 = P3_U7478 & P3_U7477 & P3_U7476 & P3_U7475; 
assign P3_U4175 = P3_U7482 & P3_U7481 & P3_U7480 & P3_U7479; 
assign P3_U4178 = P3_U7494 & P3_U7493 & P3_U7492 & P3_U7491; 
assign P3_U4179 = P3_U7498 & P3_U7497 & P3_U7496 & P3_U7495; 
assign P3_U4182 = P3_U7510 & P3_U7509 & P3_U7508 & P3_U7507; 
assign P3_U4183 = P3_U7514 & P3_U7513 & P3_U7512 & P3_U7511; 
assign P3_U4184 = P3_U7520 & P3_U7519 & P3_U7518 & P3_U7517; 
assign P3_U4185 = P3_U7524 & P3_U7523 & P3_U7522 & P3_U7521; 
assign P3_U4188 = P3_U7536 & P3_U7535 & P3_U7534 & P3_U7533; 
assign P3_U4189 = P3_U7540 & P3_U7539 & P3_U7538 & P3_U7537; 
assign P3_U4192 = P3_U7552 & P3_U7551 & P3_U7550 & P3_U7549; 
assign P3_U4193 = P3_U7556 & P3_U7555 & P3_U7554 & P3_U7553; 
assign P3_U4196 = P3_U7568 & P3_U7567 & P3_U7566 & P3_U7565; 
assign P3_U4197 = P3_U7572 & P3_U7571 & P3_U7570 & P3_U7569; 
assign P3_U4200 = P3_U7584 & P3_U7583 & P3_U7582 & P3_U7581; 
assign P3_U4201 = P3_U7588 & P3_U7587 & P3_U7586 & P3_U7585; 
assign P3_U4204 = P3_U7600 & P3_U7599 & P3_U7598 & P3_U7597; 
assign P3_U4205 = P3_U7604 & P3_U7603 & P3_U7602 & P3_U7601; 
assign P3_U4208 = P3_U7616 & P3_U7615 & P3_U7614 & P3_U7613; 
assign P3_U4209 = P3_U7620 & P3_U7619 & P3_U7618 & P3_U7617; 
assign P3_U4212 = P3_U7632 & P3_U7631 & P3_U7630 & P3_U7629; 
assign P3_U4213 = P3_U7636 & P3_U7635 & P3_U7634 & P3_U7633; 
assign P3_U4218 = P3_U7657 & P3_U7656 & P3_U7655 & P3_U7654; 
assign P3_U4219 = P3_U7661 & P3_U7660 & P3_U7659 & P3_U7658; 
assign P3_U4222 = P3_U7673 & P3_U7672 & P3_U7671 & P3_U7670; 
assign P3_U4223 = P3_U7677 & P3_U7676 & P3_U7675 & P3_U7674; 
assign P3_U4226 = P3_U7689 & P3_U7688 & P3_U7687 & P3_U7686; 
assign P3_U4227 = P3_U7693 & P3_U7692 & P3_U7691 & P3_U7690; 
assign P3_U4230 = P3_U7705 & P3_U7704 & P3_U7703 & P3_U7702; 
assign P3_U4231 = P3_U7709 & P3_U7708 & P3_U7707 & P3_U7706; 
assign P3_U4234 = P3_U7721 & P3_U7720 & P3_U7719 & P3_U7718; 
assign P3_U4235 = P3_U7725 & P3_U7724 & P3_U7723 & P3_U7722; 
assign P3_U4238 = P3_U7737 & P3_U7736 & P3_U7735 & P3_U7734; 
assign P3_U4239 = P3_U7741 & P3_U7740 & P3_U7739 & P3_U7738; 
assign P3_U4242 = P3_U7753 & P3_U7752 & P3_U7751 & P3_U7750; 
assign P3_U4243 = P3_U7757 & P3_U7756 & P3_U7755 & P3_U7754; 
assign P3_U4246 = P3_U7769 & P3_U7768 & P3_U7767 & P3_U7766; 
assign P3_U4247 = P3_U7773 & P3_U7772 & P3_U7771 & P3_U7770; 
assign P3_U4297 = ~P3_U3111; 
assign P3_U4344 = ~P3_U3103; 
assign P3_U4349 = ~P3_U3235; 
assign P3_U4646 = ~P3_U3156; 
assign P3_U4664 = ~P3_U3146; 
assign P3_U4675 = ~(P3_U2445 & P3_U4662); 
assign P3_U4680 = ~(P3_U2443 & P3_U4662); 
assign P3_U4685 = ~(P3_U2442 & P3_U4662); 
assign P3_U4690 = ~(P3_U2441 & P3_U4662); 
assign P3_U4695 = ~(P3_U2440 & P3_U4662); 
assign P3_U4700 = ~(P3_U2439 & P3_U4662); 
assign P3_U4705 = ~(P3_U2438 & P3_U4662); 
assign P3_U4710 = ~(P3_U2437 & P3_U4662); 
assign P3_U4718 = ~P3_U3152; 
assign P3_U4727 = ~(P3_U4716 & P3_U2445); 
assign P3_U4732 = ~(P3_U4716 & P3_U2443); 
assign P3_U4737 = ~(P3_U4716 & P3_U2442); 
assign P3_U4742 = ~(P3_U4716 & P3_U2441); 
assign P3_U4747 = ~(P3_U4716 & P3_U2440); 
assign P3_U4752 = ~(P3_U4716 & P3_U2439); 
assign P3_U4757 = ~(P3_U4716 & P3_U2438); 
assign P3_U4762 = ~(P3_U4716 & P3_U2437); 
assign P3_U4770 = ~P3_U3160; 
assign P3_U4779 = ~(P3_U4768 & P3_U2445); 
assign P3_U4784 = ~(P3_U4768 & P3_U2443); 
assign P3_U4789 = ~(P3_U4768 & P3_U2442); 
assign P3_U4794 = ~(P3_U4768 & P3_U2441); 
assign P3_U4799 = ~(P3_U4768 & P3_U2440); 
assign P3_U4804 = ~(P3_U4768 & P3_U2439); 
assign P3_U4809 = ~(P3_U4768 & P3_U2438); 
assign P3_U4814 = ~(P3_U4768 & P3_U2437); 
assign P3_U4830 = ~(P3_U4820 & P3_U2445); 
assign P3_U4835 = ~(P3_U4820 & P3_U2443); 
assign P3_U4840 = ~(P3_U4820 & P3_U2442); 
assign P3_U4845 = ~(P3_U4820 & P3_U2441); 
assign P3_U4850 = ~(P3_U4820 & P3_U2440); 
assign P3_U4855 = ~(P3_U4820 & P3_U2439); 
assign P3_U4860 = ~(P3_U4820 & P3_U2438); 
assign P3_U4865 = ~(P3_U4820 & P3_U2437); 
assign P3_U4873 = ~P3_U3168; 
assign P3_U4882 = ~(P3_U4871 & P3_U2445); 
assign P3_U4887 = ~(P3_U4871 & P3_U2443); 
assign P3_U4892 = ~(P3_U4871 & P3_U2442); 
assign P3_U4897 = ~(P3_U4871 & P3_U2441); 
assign P3_U4902 = ~(P3_U4871 & P3_U2440); 
assign P3_U4907 = ~(P3_U4871 & P3_U2439); 
assign P3_U4912 = ~(P3_U4871 & P3_U2438); 
assign P3_U4917 = ~(P3_U4871 & P3_U2437); 
assign P3_U4925 = ~P3_U3172; 
assign P3_U4934 = ~(P3_U4923 & P3_U2445); 
assign P3_U4939 = ~(P3_U4923 & P3_U2443); 
assign P3_U4944 = ~(P3_U4923 & P3_U2442); 
assign P3_U4949 = ~(P3_U4923 & P3_U2441); 
assign P3_U4954 = ~(P3_U4923 & P3_U2440); 
assign P3_U4959 = ~(P3_U4923 & P3_U2439); 
assign P3_U4964 = ~(P3_U4923 & P3_U2438); 
assign P3_U4969 = ~(P3_U4923 & P3_U2437); 
assign P3_U4977 = ~P3_U3176; 
assign P3_U4986 = ~(P3_U4975 & P3_U2445); 
assign P3_U4991 = ~(P3_U4975 & P3_U2443); 
assign P3_U4996 = ~(P3_U4975 & P3_U2442); 
assign P3_U5001 = ~(P3_U4975 & P3_U2441); 
assign P3_U5006 = ~(P3_U4975 & P3_U2440); 
assign P3_U5011 = ~(P3_U4975 & P3_U2439); 
assign P3_U5016 = ~(P3_U4975 & P3_U2438); 
assign P3_U5021 = ~(P3_U4975 & P3_U2437); 
assign P3_U5037 = ~(P3_U5027 & P3_U2445); 
assign P3_U5042 = ~(P3_U5027 & P3_U2443); 
assign P3_U5047 = ~(P3_U5027 & P3_U2442); 
assign P3_U5052 = ~(P3_U5027 & P3_U2441); 
assign P3_U5057 = ~(P3_U5027 & P3_U2440); 
assign P3_U5062 = ~(P3_U5027 & P3_U2439); 
assign P3_U5067 = ~(P3_U5027 & P3_U2438); 
assign P3_U5072 = ~(P3_U5027 & P3_U2437); 
assign P3_U5086 = ~(P3_U4650 & P3_U2445); 
assign P3_U5091 = ~(P3_U4650 & P3_U2443); 
assign P3_U5096 = ~(P3_U4650 & P3_U2442); 
assign P3_U5101 = ~(P3_U4650 & P3_U2441); 
assign P3_U5106 = ~(P3_U4650 & P3_U2440); 
assign P3_U5111 = ~(P3_U4650 & P3_U2439); 
assign P3_U5116 = ~(P3_U4650 & P3_U2438); 
assign P3_U5121 = ~(P3_U4650 & P3_U2437); 
assign P3_U5138 = ~(P3_U5127 & P3_U2445); 
assign P3_U5143 = ~(P3_U5127 & P3_U2443); 
assign P3_U5148 = ~(P3_U5127 & P3_U2442); 
assign P3_U5153 = ~(P3_U5127 & P3_U2441); 
assign P3_U5158 = ~(P3_U5127 & P3_U2440); 
assign P3_U5163 = ~(P3_U5127 & P3_U2439); 
assign P3_U5168 = ~(P3_U5127 & P3_U2438); 
assign P3_U5173 = ~(P3_U5127 & P3_U2437); 
assign P3_U5190 = ~(P3_U5179 & P3_U2445); 
assign P3_U5195 = ~(P3_U5179 & P3_U2443); 
assign P3_U5200 = ~(P3_U5179 & P3_U2442); 
assign P3_U5205 = ~(P3_U5179 & P3_U2441); 
assign P3_U5210 = ~(P3_U5179 & P3_U2440); 
assign P3_U5215 = ~(P3_U5179 & P3_U2439); 
assign P3_U5220 = ~(P3_U5179 & P3_U2438); 
assign P3_U5225 = ~(P3_U5179 & P3_U2437); 
assign P3_U5232 = ~P3_U3072; 
assign P3_U5240 = ~(P3_U5231 & P3_U2445); 
assign P3_U5245 = ~(P3_U5231 & P3_U2443); 
assign P3_U5250 = ~(P3_U5231 & P3_U2442); 
assign P3_U5255 = ~(P3_U5231 & P3_U2441); 
assign P3_U5260 = ~(P3_U5231 & P3_U2440); 
assign P3_U5265 = ~(P3_U5231 & P3_U2439); 
assign P3_U5270 = ~(P3_U5231 & P3_U2438); 
assign P3_U5275 = ~(P3_U5231 & P3_U2437); 
assign P3_U5291 = ~(P3_U5281 & P3_U2445); 
assign P3_U5296 = ~(P3_U5281 & P3_U2443); 
assign P3_U5301 = ~(P3_U5281 & P3_U2442); 
assign P3_U5306 = ~(P3_U5281 & P3_U2441); 
assign P3_U5311 = ~(P3_U5281 & P3_U2440); 
assign P3_U5316 = ~(P3_U5281 & P3_U2439); 
assign P3_U5321 = ~(P3_U5281 & P3_U2438); 
assign P3_U5326 = ~(P3_U5281 & P3_U2437); 
assign P3_U5342 = ~(P3_U5332 & P3_U2445); 
assign P3_U5347 = ~(P3_U5332 & P3_U2443); 
assign P3_U5352 = ~(P3_U5332 & P3_U2442); 
assign P3_U5357 = ~(P3_U5332 & P3_U2441); 
assign P3_U5362 = ~(P3_U5332 & P3_U2440); 
assign P3_U5367 = ~(P3_U5332 & P3_U2439); 
assign P3_U5372 = ~(P3_U5332 & P3_U2438); 
assign P3_U5377 = ~(P3_U5332 & P3_U2437); 
assign P3_U5393 = ~(P3_U5383 & P3_U2445); 
assign P3_U5398 = ~(P3_U5383 & P3_U2443); 
assign P3_U5403 = ~(P3_U5383 & P3_U2442); 
assign P3_U5408 = ~(P3_U5383 & P3_U2441); 
assign P3_U5413 = ~(P3_U5383 & P3_U2440); 
assign P3_U5418 = ~(P3_U5383 & P3_U2439); 
assign P3_U5423 = ~(P3_U5383 & P3_U2438); 
assign P3_U5428 = ~(P3_U5383 & P3_U2437); 
assign P3_U5435 = ~P3_U3073; 
assign P3_U5443 = ~(P3_U5434 & P3_U2445); 
assign P3_U5448 = ~(P3_U5434 & P3_U2443); 
assign P3_U5453 = ~(P3_U5434 & P3_U2442); 
assign P3_U5458 = ~(P3_U5434 & P3_U2441); 
assign P3_U5463 = ~(P3_U5434 & P3_U2440); 
assign P3_U5468 = ~(P3_U5434 & P3_U2439); 
assign P3_U5473 = ~(P3_U5434 & P3_U2438); 
assign P3_U5478 = ~(P3_U5434 & P3_U2437); 
assign P3_U5508 = ~(P3_U4522 & P3_U4607 & P3_U4488); 
assign P3_U5513 = ~(P3_U4522 & P3_U4607); 
assign P3_U5514 = ~(P3_U4607 & P3_U3218); 
assign P3_U5516 = ~(P3_U4573 & P3_U4505); 
assign P3_U5519 = ~(P3_U4607 & P3_U3104 & P3_U4573); 
assign P3_U5600 = ~(P3_U4322 & P3_U3156); 
assign P3_U7386 = ~(P3_U4488 & P3_STATE2_REG_2__SCAN_IN); 
assign P3_U7916 = ~(P3_U4505 & P3_U3106); 
assign P3_U7917 = ~(P3_U4488 & P3_U4522); 
assign P3_U7974 = ~(P3_U4573 & P3_U4590); 
assign P2_U2451 = P2_U4601 & P2_U2457 & P2_U2438; 
assign P2_U2590 = P2_U5590 & P2_U2436; 
assign P2_U2607 = ~(P2_U4226 & P2_U4225 & P2_U4224 & P2_U4223); 
assign P2_U2608 = ~(P2_U4222 & P2_U4221 & P2_U4220 & P2_U4219); 
assign P2_U2609 = ~(P2_U4218 & P2_U4217 & P2_U4216 & P2_U4215); 
assign P2_U2610 = ~(P2_U4214 & P2_U4213 & P2_U4212 & P2_U4211); 
assign P2_U2611 = ~(P2_U4210 & P2_U4209 & P2_U4208 & P2_U4207); 
assign P2_U2612 = ~(P2_U4206 & P2_U4205 & P2_U4204 & P2_U4203); 
assign P2_U2613 = ~(P2_U4202 & P2_U4201 & P2_U4200 & P2_U4199); 
assign P2_U2614 = ~(P2_U4198 & P2_U4197 & P2_U4196 & P2_U4195); 
assign P2_U2681 = ~(P2_U7166 & P2_U4275); 
assign P2_U2707 = ~(P2_U4391 & P2_U7734); 
assign P2_U3242 = ~(P2_U4194 & P2_U4193 & P2_U4192 & P2_U4191); 
assign P2_U3282 = ~(P2_U2457 & P2_U7869 & P2_U4476); 
assign P2_U3293 = ~(P2_U2357 & P2_U3280); 
assign P2_U3539 = ~(P2_U4056 & P2_U2357); 
assign P2_U3550 = ~(P2_U4427 & P2_STATE2_REG_0__SCAN_IN); 
assign P2_U3575 = ~(P2_U4419 & P2_U7871); 
assign P2_U3576 = ~(P2_U4419 & P2_U3279); 
assign P2_U3656 = ~(P2_U8368 & P2_U8367); 
assign P2_U3709 = P2_U3710 & P2_U4417; 
assign P2_U3875 = P2_U3874 & P2_U4429; 
assign P2_U3876 = P2_U4429 & P2_U3279; 
assign P2_U3879 = P2_U5587 & P2_U5588 & P2_U3281; 
assign P2_U3886 = P2_U4601 & P2_U2449; 
assign P2_U4058 = P2_U2374 & P2_U4417; 
assign P2_U4185 = P2_U6848 & P2_U3301; 
assign P2_U4227 = P2_U7011 & P2_U7010 & P2_U7009 & P2_U7008; 
assign P2_U4228 = P2_U7015 & P2_U7014 & P2_U7013 & P2_U7012; 
assign P2_U4231 = P2_U7027 & P2_U7026 & P2_U7025 & P2_U7024; 
assign P2_U4232 = P2_U7031 & P2_U7030 & P2_U7029 & P2_U7028; 
assign P2_U4235 = P2_U7043 & P2_U7042 & P2_U7041 & P2_U7040; 
assign P2_U4236 = P2_U7047 & P2_U7046 & P2_U7045 & P2_U7044; 
assign P2_U4239 = P2_U7059 & P2_U7058 & P2_U7057 & P2_U7056; 
assign P2_U4240 = P2_U7063 & P2_U7062 & P2_U7061 & P2_U7060; 
assign P2_U4243 = P2_U7075 & P2_U7074 & P2_U7073 & P2_U7072; 
assign P2_U4244 = P2_U7079 & P2_U7078 & P2_U7077 & P2_U7076; 
assign P2_U4247 = P2_U7091 & P2_U7090 & P2_U7089 & P2_U7088; 
assign P2_U4248 = P2_U7095 & P2_U7094 & P2_U7093 & P2_U7092; 
assign P2_U4251 = P2_U7107 & P2_U7106 & P2_U7105 & P2_U7104; 
assign P2_U4252 = P2_U7111 & P2_U7110 & P2_U7109 & P2_U7108; 
assign P2_U4255 = P2_U7123 & P2_U7122 & P2_U7121 & P2_U7120; 
assign P2_U4256 = P2_U7127 & P2_U7126 & P2_U7125 & P2_U7124; 
assign P2_U4340 = P2_U7426 & P2_U4414 & P2_U7428; 
assign P2_U4376 = P2_U3255 & P2_U6845; 
assign P2_U4387 = P2_U7736 & P2_STATE2_REG_0__SCAN_IN; 
assign P2_U4413 = ~(P2_U4337 & P2_U4601); 
assign P2_U4420 = ~P2_U3288; 
assign P2_U4422 = ~(P2_U2376 & P2_U3278 & P2_U2450); 
assign P2_U4596 = ~P2_U3527; 
assign P2_U4598 = ~(P2_U4597 & P2_U3265); 
assign P2_U4599 = ~(P2_U2359 & P2_U3527); 
assign P2_U5572 = ~P2_U3574; 
assign P2_U5575 = ~(P2_U2357 & P2_U7871); 
assign P2_U5576 = ~(P2_U4417 & P2_U3574); 
assign P2_U5592 = ~(P2_U3521 & P2_U5591 & P2_U5573 & P2_U5571); 
assign P2_U5593 = ~(P2_U4417 & P2_U3574); 
assign P2_U5599 = ~(P2_U4427 & P2_U5598); 
assign P2_U5602 = ~(P2_U3527 & P2_U3278); 
assign P2_U5624 = ~(P2_U2449 & P2_U7861 & P2_U4429); 
assign P2_U6850 = ~(U211 & P2_U6846); 
assign P2_U7217 = ~(P2_U4288 & P2_U4287 & P2_U4286 & P2_U4285); 
assign P2_U7251 = ~(P2_U4296 & P2_U4295 & P2_U4294 & P2_U4293); 
assign P2_U7285 = ~(P2_U4304 & P2_U4303 & P2_U4302 & P2_U4301); 
assign P2_U7319 = ~(P2_U4312 & P2_U4311 & P2_U4310 & P2_U4309); 
assign P2_U7353 = ~(P2_U4320 & P2_U4319 & P2_U4318 & P2_U4317); 
assign P2_U7387 = ~(P2_U4328 & P2_U4327 & P2_U4326 & P2_U4325); 
assign P2_U7421 = ~(P2_U4336 & P2_U4335 & P2_U4334 & P2_U4333); 
assign P2_U7434 = ~(P2_U2353 & P2_REIP_REG_9__SCAN_IN); 
assign P2_U7435 = ~(P2_U4412 & P2_EAX_REG_9__SCAN_IN); 
assign P2_U7438 = ~(P2_U2353 & P2_REIP_REG_8__SCAN_IN); 
assign P2_U7439 = ~(P2_U4412 & P2_EAX_REG_8__SCAN_IN); 
assign P2_U7442 = ~(P2_U2353 & P2_REIP_REG_7__SCAN_IN); 
assign P2_U7443 = ~(P2_U4412 & P2_EAX_REG_7__SCAN_IN); 
assign P2_U7445 = ~(P2_U2353 & P2_REIP_REG_6__SCAN_IN); 
assign P2_U7446 = ~(P2_U4412 & P2_EAX_REG_6__SCAN_IN); 
assign P2_U7448 = ~(P2_U2353 & P2_REIP_REG_5__SCAN_IN); 
assign P2_U7449 = ~(P2_U4412 & P2_EAX_REG_5__SCAN_IN); 
assign P2_U7451 = ~(P2_U2353 & P2_REIP_REG_4__SCAN_IN); 
assign P2_U7452 = ~(P2_U4412 & P2_EAX_REG_4__SCAN_IN); 
assign P2_U7454 = ~(P2_U2353 & P2_REIP_REG_31__SCAN_IN); 
assign P2_U7455 = ~(P2_U4412 & P2_EAX_REG_31__SCAN_IN); 
assign P2_U7457 = ~(P2_U2353 & P2_REIP_REG_30__SCAN_IN); 
assign P2_U7458 = ~(P2_U4412 & P2_EAX_REG_30__SCAN_IN); 
assign P2_U7460 = ~(P2_U2353 & P2_REIP_REG_3__SCAN_IN); 
assign P2_U7461 = ~(P2_U4412 & P2_EAX_REG_3__SCAN_IN); 
assign P2_U7463 = ~(P2_U2353 & P2_REIP_REG_29__SCAN_IN); 
assign P2_U7464 = ~(P2_U4412 & P2_EAX_REG_29__SCAN_IN); 
assign P2_U7466 = ~(P2_U2353 & P2_REIP_REG_28__SCAN_IN); 
assign P2_U7467 = ~(P2_U4412 & P2_EAX_REG_28__SCAN_IN); 
assign P2_U7469 = ~(P2_U2353 & P2_REIP_REG_27__SCAN_IN); 
assign P2_U7470 = ~(P2_U4412 & P2_EAX_REG_27__SCAN_IN); 
assign P2_U7472 = ~(P2_U2353 & P2_REIP_REG_26__SCAN_IN); 
assign P2_U7473 = ~(P2_U4412 & P2_EAX_REG_26__SCAN_IN); 
assign P2_U7475 = ~(P2_U2353 & P2_REIP_REG_25__SCAN_IN); 
assign P2_U7476 = ~(P2_U4412 & P2_EAX_REG_25__SCAN_IN); 
assign P2_U7478 = ~(P2_U2353 & P2_REIP_REG_24__SCAN_IN); 
assign P2_U7479 = ~(P2_U4412 & P2_EAX_REG_24__SCAN_IN); 
assign P2_U7481 = ~(P2_U2353 & P2_REIP_REG_23__SCAN_IN); 
assign P2_U7482 = ~(P2_U4412 & P2_EAX_REG_23__SCAN_IN); 
assign P2_U7484 = ~(P2_U2353 & P2_REIP_REG_22__SCAN_IN); 
assign P2_U7485 = ~(P2_U4412 & P2_EAX_REG_22__SCAN_IN); 
assign P2_U7487 = ~(P2_U2353 & P2_REIP_REG_21__SCAN_IN); 
assign P2_U7488 = ~(P2_U4412 & P2_EAX_REG_21__SCAN_IN); 
assign P2_U7490 = ~(P2_U2353 & P2_REIP_REG_20__SCAN_IN); 
assign P2_U7491 = ~(P2_U4412 & P2_EAX_REG_20__SCAN_IN); 
assign P2_U7493 = ~(P2_U2353 & P2_REIP_REG_2__SCAN_IN); 
assign P2_U7494 = ~(P2_U4412 & P2_EAX_REG_2__SCAN_IN); 
assign P2_U7496 = ~(P2_U2353 & P2_REIP_REG_19__SCAN_IN); 
assign P2_U7497 = ~(P2_U4412 & P2_EAX_REG_19__SCAN_IN); 
assign P2_U7499 = ~(P2_U2353 & P2_REIP_REG_18__SCAN_IN); 
assign P2_U7500 = ~(P2_U4412 & P2_EAX_REG_18__SCAN_IN); 
assign P2_U7502 = ~(P2_U2353 & P2_REIP_REG_17__SCAN_IN); 
assign P2_U7503 = ~(P2_U4412 & P2_EAX_REG_17__SCAN_IN); 
assign P2_U7505 = ~(P2_U2353 & P2_REIP_REG_16__SCAN_IN); 
assign P2_U7506 = ~(P2_U4412 & P2_EAX_REG_16__SCAN_IN); 
assign P2_U7508 = ~(P2_U2353 & P2_REIP_REG_15__SCAN_IN); 
assign P2_U7509 = ~(P2_U4412 & P2_EAX_REG_15__SCAN_IN); 
assign P2_U7512 = ~(P2_U2353 & P2_REIP_REG_14__SCAN_IN); 
assign P2_U7513 = ~(P2_U4412 & P2_EAX_REG_14__SCAN_IN); 
assign P2_U7516 = ~(P2_U2353 & P2_REIP_REG_13__SCAN_IN); 
assign P2_U7517 = ~(P2_U4412 & P2_EAX_REG_13__SCAN_IN); 
assign P2_U7520 = ~(P2_U2353 & P2_REIP_REG_12__SCAN_IN); 
assign P2_U7521 = ~(P2_U4412 & P2_EAX_REG_12__SCAN_IN); 
assign P2_U7524 = ~(P2_U2353 & P2_REIP_REG_11__SCAN_IN); 
assign P2_U7525 = ~(P2_U4412 & P2_EAX_REG_11__SCAN_IN); 
assign P2_U7528 = ~(P2_U2353 & P2_REIP_REG_10__SCAN_IN); 
assign P2_U7529 = ~(P2_U4412 & P2_EAX_REG_10__SCAN_IN); 
assign P2_U7532 = ~(P2_U2353 & P2_REIP_REG_1__SCAN_IN); 
assign P2_U7533 = ~(P2_U4412 & P2_EAX_REG_1__SCAN_IN); 
assign P2_U7535 = ~(P2_U2353 & P2_REIP_REG_0__SCAN_IN); 
assign P2_U7536 = ~(P2_U4412 & P2_EAX_REG_0__SCAN_IN); 
assign P2_U7579 = ~(P2_U2617 & P2_U2450); 
assign P2_U7581 = ~(P2_U3525 & P2_U6845 & P2_U7867); 
assign P2_U7730 = ~(P2_R2238_U21 & P2_U2356); 
assign P2_U7740 = ~(P2_U3521 & P2_U7744 & P2_U5573 & P2_U5571); 
assign P2_U7882 = ~(P2_U5590 & P2_U4428); 
assign P2_U7883 = ~(P2_U5596 & P2_U3525); 
assign P2_U8068 = ~(P2_U7859 & P2_U5574); 
assign P2_U8074 = ~(P2_U3280 & P2_U5586); 
assign P2_U8118 = ~(P2_U8117 & P2_U8116); 
assign P2_U8357 = ~(P2_R2238_U21 & P2_U3283); 
assign P2_U8358 = ~(P2_SUB_450_U19 & P2_U4417); 
assign P2_U8360 = ~(P2_SUB_450_U20 & P2_U4417); 
assign P2_U8429 = ~(P2_R2238_U21 & P2_U3269); 
assign P1_U2431 = P1_U4199 & P1_U7494; 
assign P1_U3227 = ~(P1_U4001 & P1_U4000 & P1_U3999 & P1_U3998); 
assign P1_U3228 = ~(P1_U3997 & P1_U3996 & P1_U3995 & P1_U3994); 
assign P1_U3229 = ~(P1_U3993 & P1_U3992 & P1_U3991 & P1_U3990); 
assign P1_U3230 = ~(P1_U3989 & P1_U3988 & P1_U3987 & P1_U3986); 
assign P1_U3231 = ~(P1_U3985 & P1_U3984 & P1_U3983 & P1_U3982); 
assign P1_U3232 = ~(P1_U3981 & P1_U3980 & P1_U3979 & P1_U3978); 
assign P1_U3233 = ~(P1_U3977 & P1_U3976 & P1_U3975 & P1_U3974); 
assign P1_U3234 = ~(P1_U3973 & P1_U3972 & P1_U3971 & P1_U3970); 
assign P1_U3288 = ~(P1_U4249 & P1_U2447); 
assign P1_U3392 = ~(P1_U5490 & P1_U5489 & P1_U7628); 
assign P1_U3399 = ~(P1_U4199 & P1_U4477 & P1_U4234); 
assign P1_U3400 = ~(P1_U2449 & P1_U2447); 
assign P1_U3410 = ~(P1_U4253 & P1_U3278); 
assign P1_U3420 = ~(P1_U4206 & P1_U4477); 
assign P1_U3427 = ~(P1_U4249 & P1_U3886 & P1_U2452 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U3428 = ~(P1_U3866 & P1_U2447); 
assign P1_U3434 = ~(P1_U4206 & P1_U3271); 
assign P1_U3447 = ~(P1_U4231 & P1_U4400 & P1_U4250); 
assign P1_U3448 = ~(P1_U4231 & P1_U3278 & P1_U4250); 
assign P1_U3568 = P1_U4377 & P1_U4208; 
assign P1_U3578 = P1_U4249 & P1_U3283; 
assign P1_U3736 = P1_U5471 & P1_U5472; 
assign P1_U3756 = P1_U5563 & P1_U5561; 
assign P1_U3867 = P1_U4208 & P1_U2368; 
assign P1_U3969 = P1_U4235 & P1_U4206; 
assign P1_U4007 = P1_U6762 & P1_U6761; 
assign P1_U4031 = P1_U6903 & P1_U6902 & P1_U6901 & P1_U6900; 
assign P1_U4032 = P1_U6907 & P1_U6906 & P1_U6905 & P1_U6904; 
assign P1_U4035 = P1_U6921 & P1_U6920 & P1_U6919 & P1_U6918; 
assign P1_U4036 = P1_U6925 & P1_U6924 & P1_U6923 & P1_U6922; 
assign P1_U4039 = P1_U6952 & P1_U6951 & P1_U6950 & P1_U6949; 
assign P1_U4040 = P1_U6956 & P1_U6955 & P1_U6954 & P1_U6953; 
assign P1_U4043 = P1_U6969 & P1_U6968 & P1_U6967 & P1_U6966; 
assign P1_U4044 = P1_U6973 & P1_U6972 & P1_U6971 & P1_U6970; 
assign P1_U4047 = P1_U6986 & P1_U6985 & P1_U6984 & P1_U6983; 
assign P1_U4048 = P1_U6990 & P1_U6989 & P1_U6988 & P1_U6987; 
assign P1_U4051 = P1_U7003 & P1_U7002 & P1_U7001 & P1_U7000; 
assign P1_U4052 = P1_U7614 & P1_U7006 & P1_U7005 & P1_U7004; 
assign P1_U4055 = P1_U7018 & P1_U7017 & P1_U7016 & P1_U7015; 
assign P1_U4056 = P1_U7022 & P1_U7021 & P1_U7020 & P1_U7019; 
assign P1_U4059 = P1_U7035 & P1_U7034 & P1_U7033 & P1_U7032; 
assign P1_U4060 = P1_U7039 & P1_U7038 & P1_U7037 & P1_U7036; 
assign P1_U4062 = P1_U7062 & P1_STATE2_REG_0__SCAN_IN; 
assign P1_U4123 = P1_U7231 & P1_U7230 & P1_U7229 & P1_U7228; 
assign P1_U4124 = P1_U7235 & P1_U7234 & P1_U7233 & P1_U7232; 
assign P1_U4127 = P1_U7248 & P1_U7247 & P1_U7246 & P1_U7245; 
assign P1_U4128 = P1_U7252 & P1_U7251 & P1_U7250 & P1_U7249; 
assign P1_U4131 = P1_U7265 & P1_U7264 & P1_U7263 & P1_U7262; 
assign P1_U4132 = P1_U7269 & P1_U7268 & P1_U7267 & P1_U7266; 
assign P1_U4135 = P1_U7282 & P1_U7281 & P1_U7280 & P1_U7279; 
assign P1_U4136 = P1_U7619 & P1_U7285 & P1_U7284 & P1_U7283; 
assign P1_U4139 = P1_U7297 & P1_U7296 & P1_U7295 & P1_U7294; 
assign P1_U4140 = P1_U7301 & P1_U7300 & P1_U7299 & P1_U7298; 
assign P1_U4143 = P1_U7314 & P1_U7313 & P1_U7312 & P1_U7311; 
assign P1_U4144 = P1_U7318 & P1_U7317 & P1_U7316 & P1_U7315; 
assign P1_U4147 = P1_U7331 & P1_U7330 & P1_U7329 & P1_U7328; 
assign P1_U4148 = P1_U7335 & P1_U7334 & P1_U7333 & P1_U7332; 
assign P1_U4151 = P1_U7348 & P1_U7347 & P1_U7346 & P1_U7345; 
assign P1_U4152 = P1_U7352 & P1_U7351 & P1_U7350 & P1_U7349; 
assign P1_U4163 = P1_U7373 & P1_STATE2_REG_0__SCAN_IN; 
assign P1_U4164 = P1_U7375 & P1_U2603; 
assign P1_U4167 = P1_U7389 & P1_U7388 & P1_U7387; 
assign P1_U4197 = ~P1_U3396; 
assign P1_U4201 = ~P1_U3422; 
assign P1_U4256 = ~P1_U3291; 
assign P1_U4262 = ~P1_U3286; 
assign P1_U4263 = ~(P1_U4236 & P1_U4399); 
assign P1_U4264 = ~P1_U3411; 
assign P1_U4501 = ~(P1_U4500 & P1_U3257); 
assign P1_U4504 = ~(P1_U4196 & P1_U3286); 
assign P1_U4785 = ~(P1_U4779 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U4900 = ~(P1_U4894 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U5013 = ~(P1_U5008 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U5128 = ~(P1_U5122 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U5243 = ~(P1_U5237 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U5358 = ~(P1_U5352 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U5461 = ~P1_U3423; 
assign P1_U5464 = ~P1_U3244; 
assign P1_U5468 = ~(P1_U4208 & P1_U5462); 
assign P1_U5492 = ~(P1_U5491 & P1_U4171); 
assign P1_U5496 = ~(P1_U4208 & P1_U5462); 
assign P1_U5498 = ~(P1_U5495 & P1_U3271); 
assign P1_U5500 = ~(P1_U4190 & P1_U3244); 
assign P1_U6364 = ~(P1_U4249 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U6605 = ~(P1_U4208 & P1_U6604); 
assign P1_U6615 = ~(P1_U3968 & P1_U3291); 
assign P1_U6747 = ~(P1_U4188 & P1_EAX_REG_9__SCAN_IN); 
assign P1_U6750 = ~(P1_U4188 & P1_EAX_REG_8__SCAN_IN); 
assign P1_U6753 = ~(P1_U4188 & P1_EAX_REG_7__SCAN_IN); 
assign P1_U6756 = ~(P1_U4188 & P1_EAX_REG_6__SCAN_IN); 
assign P1_U6760 = ~(P1_U4188 & P1_EAX_REG_5__SCAN_IN); 
assign P1_U6764 = ~(P1_U4188 & P1_EAX_REG_4__SCAN_IN); 
assign P1_U6767 = ~(P1_U2353 & P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P1_U6768 = ~(P1_U4188 & P1_EAX_REG_31__SCAN_IN); 
assign P1_U6772 = ~(P1_U4188 & P1_EAX_REG_30__SCAN_IN); 
assign P1_U6776 = ~(P1_U4188 & P1_EAX_REG_3__SCAN_IN); 
assign P1_U6779 = ~(P1_U2353 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P1_U6781 = ~(P1_U4188 & P1_EAX_REG_29__SCAN_IN); 
assign P1_U6785 = ~(P1_U4188 & P1_EAX_REG_28__SCAN_IN); 
assign P1_U6789 = ~(P1_U4188 & P1_EAX_REG_27__SCAN_IN); 
assign P1_U6793 = ~(P1_U4188 & P1_EAX_REG_26__SCAN_IN); 
assign P1_U6797 = ~(P1_U4188 & P1_EAX_REG_25__SCAN_IN); 
assign P1_U6801 = ~(P1_U4188 & P1_EAX_REG_24__SCAN_IN); 
assign P1_U6805 = ~(P1_U4188 & P1_EAX_REG_23__SCAN_IN); 
assign P1_U6809 = ~(P1_U4188 & P1_EAX_REG_22__SCAN_IN); 
assign P1_U6813 = ~(P1_U4188 & P1_EAX_REG_21__SCAN_IN); 
assign P1_U6817 = ~(P1_U4188 & P1_EAX_REG_20__SCAN_IN); 
assign P1_U6821 = ~(P1_U4188 & P1_EAX_REG_2__SCAN_IN); 
assign P1_U6824 = ~(P1_U2353 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_U6826 = ~(P1_U4188 & P1_EAX_REG_19__SCAN_IN); 
assign P1_U6830 = ~(P1_U4188 & P1_EAX_REG_18__SCAN_IN); 
assign P1_U6834 = ~(P1_U4188 & P1_EAX_REG_17__SCAN_IN); 
assign P1_U6838 = ~(P1_U4188 & P1_EAX_REG_16__SCAN_IN); 
assign P1_U6841 = ~(P1_U4188 & P1_EAX_REG_15__SCAN_IN); 
assign P1_U6844 = ~(P1_U4188 & P1_EAX_REG_14__SCAN_IN); 
assign P1_U6847 = ~(P1_U4188 & P1_EAX_REG_13__SCAN_IN); 
assign P1_U6850 = ~(P1_U4188 & P1_EAX_REG_12__SCAN_IN); 
assign P1_U6853 = ~(P1_U4188 & P1_EAX_REG_11__SCAN_IN); 
assign P1_U6856 = ~(P1_U4188 & P1_EAX_REG_10__SCAN_IN); 
assign P1_U6860 = ~(P1_U4188 & P1_EAX_REG_1__SCAN_IN); 
assign P1_U6863 = ~(P1_U2353 & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U6865 = ~(P1_U4188 & P1_EAX_REG_0__SCAN_IN); 
assign P1_U6868 = ~(P1_U2353 & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U7084 = ~(P1_U4073 & P1_U4191); 
assign P1_U7089 = ~(P1_U4189 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U7354 = ~(P1_U4231 & P1_U2354 & P1_U4234); 
assign P1_U7360 = ~(P1_U4208 & P1_U7088); 
assign P1_U7361 = ~(P1_U4160 & P1_U4208); 
assign P1_U7371 = ~(P1_SUB_450_U21 & P1_U2354); 
assign P1_U7382 = ~(P1_R2238_U21 & P1_U4192); 
assign P1_U7392 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P1_U7393 = ~(P1_U7390 & P1_EBX_REG_9__SCAN_IN); 
assign P1_U7394 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P1_U7395 = ~(P1_U7390 & P1_EBX_REG_8__SCAN_IN); 
assign P1_U7396 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P1_U7397 = ~(P1_U7390 & P1_EBX_REG_7__SCAN_IN); 
assign P1_U7398 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P1_U7399 = ~(P1_U7390 & P1_EBX_REG_6__SCAN_IN); 
assign P1_U7400 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P1_U7401 = ~(P1_U7390 & P1_EBX_REG_5__SCAN_IN); 
assign P1_U7402 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P1_U7403 = ~(P1_U7390 & P1_EBX_REG_4__SCAN_IN); 
assign P1_U7404 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P1_U7405 = ~(P1_U7390 & P1_EBX_REG_31__SCAN_IN); 
assign P1_U7406 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P1_U7407 = ~(P1_U7390 & P1_EBX_REG_30__SCAN_IN); 
assign P1_U7408 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P1_U7409 = ~(P1_U7390 & P1_EBX_REG_3__SCAN_IN); 
assign P1_U7410 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P1_U7411 = ~(P1_U7390 & P1_EBX_REG_29__SCAN_IN); 
assign P1_U7412 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P1_U7413 = ~(P1_U7390 & P1_EBX_REG_28__SCAN_IN); 
assign P1_U7414 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P1_U7415 = ~(P1_U7390 & P1_EBX_REG_27__SCAN_IN); 
assign P1_U7416 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P1_U7417 = ~(P1_U7390 & P1_EBX_REG_26__SCAN_IN); 
assign P1_U7418 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P1_U7419 = ~(P1_U7390 & P1_EBX_REG_25__SCAN_IN); 
assign P1_U7420 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P1_U7421 = ~(P1_U7390 & P1_EBX_REG_24__SCAN_IN); 
assign P1_U7422 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P1_U7423 = ~(P1_U7390 & P1_EBX_REG_23__SCAN_IN); 
assign P1_U7424 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P1_U7425 = ~(P1_U7390 & P1_EBX_REG_22__SCAN_IN); 
assign P1_U7426 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P1_U7427 = ~(P1_U7390 & P1_EBX_REG_21__SCAN_IN); 
assign P1_U7428 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P1_U7429 = ~(P1_U7390 & P1_EBX_REG_20__SCAN_IN); 
assign P1_U7430 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P1_U7431 = ~(P1_U7390 & P1_EBX_REG_2__SCAN_IN); 
assign P1_U7432 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P1_U7433 = ~(P1_U7390 & P1_EBX_REG_19__SCAN_IN); 
assign P1_U7434 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P1_U7435 = ~(P1_U7390 & P1_EBX_REG_18__SCAN_IN); 
assign P1_U7436 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P1_U7437 = ~(P1_U7390 & P1_EBX_REG_17__SCAN_IN); 
assign P1_U7438 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P1_U7439 = ~(P1_U7390 & P1_EBX_REG_16__SCAN_IN); 
assign P1_U7440 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P1_U7441 = ~(P1_U7390 & P1_EBX_REG_15__SCAN_IN); 
assign P1_U7442 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P1_U7443 = ~(P1_U7390 & P1_EBX_REG_14__SCAN_IN); 
assign P1_U7444 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P1_U7445 = ~(P1_U7390 & P1_EBX_REG_13__SCAN_IN); 
assign P1_U7446 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P1_U7447 = ~(P1_U7390 & P1_EBX_REG_12__SCAN_IN); 
assign P1_U7448 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P1_U7449 = ~(P1_U7390 & P1_EBX_REG_11__SCAN_IN); 
assign P1_U7450 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P1_U7451 = ~(P1_U7390 & P1_EBX_REG_10__SCAN_IN); 
assign P1_U7452 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P1_U7453 = ~(P1_U7390 & P1_EBX_REG_1__SCAN_IN); 
assign P1_U7454 = ~(P1_U7391 & P1_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P1_U7455 = ~(P1_U7390 & P1_EBX_REG_0__SCAN_IN); 
assign P1_U7475 = ~(P1_U4236 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U7489 = ~(P1_U4236 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U7493 = ~P1_U3279; 
assign P1_U7630 = ~(P1_U4208 & P1_U7490); 
assign P1_U7700 = ~(P1_U5467 & P1_U4171); 
assign P3_ADD_526_U51 = ~(P3_ADD_526_U142 & P3_ADD_526_U141); 
assign P3_ADD_526_U52 = ~(P3_ADD_526_U144 & P3_ADD_526_U143); 
assign P3_ADD_526_U113 = ~P3_ADD_526_U22; 
assign P3_ADD_526_U140 = ~P3_ADD_526_U110; 
assign P3_ADD_526_U200 = ~(P3_ADD_526_U22 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_526_U201 = ~(P3_ADD_526_U110 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_552_U51 = ~(P3_ADD_552_U142 & P3_ADD_552_U141); 
assign P3_ADD_552_U52 = ~(P3_ADD_552_U144 & P3_ADD_552_U143); 
assign P3_ADD_552_U113 = ~P3_ADD_552_U22; 
assign P3_ADD_552_U140 = ~P3_ADD_552_U110; 
assign P3_ADD_552_U200 = ~(P3_ADD_552_U22 & P3_EBX_REG_11__SCAN_IN); 
assign P3_ADD_552_U201 = ~(P3_ADD_552_U110 & P3_EBX_REG_10__SCAN_IN); 
assign P3_ADD_546_U51 = ~(P3_ADD_546_U142 & P3_ADD_546_U141); 
assign P3_ADD_546_U52 = ~(P3_ADD_546_U144 & P3_ADD_546_U143); 
assign P3_ADD_546_U113 = ~P3_ADD_546_U22; 
assign P3_ADD_546_U140 = ~P3_ADD_546_U110; 
assign P3_ADD_546_U200 = ~(P3_ADD_546_U22 & P3_EAX_REG_11__SCAN_IN); 
assign P3_ADD_546_U201 = ~(P3_ADD_546_U110 & P3_EAX_REG_10__SCAN_IN); 
assign P3_GTE_401_U7 = P3_SUB_401_U21 & P3_GTE_401_U9; 
assign P3_ADD_391_1180_U4 = ~P3_U2613; 
assign P3_ADD_391_1180_U7 = ~P3_U2614; 
assign P3_ADD_391_1180_U9 = ~P3_U2615; 
assign P3_ADD_391_1180_U11 = ~P3_U2616; 
assign P3_ADD_391_1180_U13 = ~P3_U2617; 
assign P3_ADD_391_1180_U15 = ~P3_U2618; 
assign P3_ADD_391_1180_U17 = ~P3_U2619; 
assign P3_ADD_391_1180_U26 = ~P3_U2620; 
assign P3_ADD_476_U65 = ~(P3_ADD_476_U130 & P3_ADD_476_U129); 
assign P3_ADD_476_U98 = ~P3_ADD_476_U14; 
assign P3_ADD_476_U127 = ~(P3_ADD_476_U14 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_GTE_390_U7 = P3_SUB_390_U21 & P3_GTE_390_U9; 
assign P3_ADD_531_U69 = ~(P3_ADD_531_U137 & P3_ADD_531_U136); 
assign P3_ADD_531_U102 = ~P3_ADD_531_U15; 
assign P3_ADD_531_U134 = ~(P3_ADD_531_U15 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_SUB_320_U89 = ~(P3_SUB_320_U84 & P3_SUB_320_U56); 
assign P3_SUB_320_U133 = ~(P3_SUB_320_U84 & P3_SUB_320_U56); 
assign P3_ADD_318_U65 = ~(P3_ADD_318_U130 & P3_ADD_318_U129); 
assign P3_ADD_318_U98 = ~P3_ADD_318_U14; 
assign P3_ADD_318_U127 = ~(P3_ADD_318_U14 & P3_PHYADDRPOINTER_REG_7__SCAN_IN); 
assign P3_SUB_370_U16 = ~(P3_SUB_370_U41 & P3_SUB_370_U40); 
assign P3_SUB_370_U55 = ~(P3_SUB_370_U38 & P3_SUB_370_U54); 
assign P3_ADD_315_U62 = ~(P3_ADD_315_U124 & P3_ADD_315_U123); 
assign P3_ADD_315_U95 = ~P3_ADD_315_U14; 
assign P3_ADD_315_U121 = ~(P3_ADD_315_U14 & P3_PHYADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_467_U65 = ~(P3_ADD_467_U130 & P3_ADD_467_U129); 
assign P3_ADD_467_U98 = ~P3_ADD_467_U14; 
assign P3_ADD_467_U127 = ~(P3_ADD_467_U14 & P3_REIP_REG_7__SCAN_IN); 
assign P3_ADD_430_U65 = ~(P3_ADD_430_U130 & P3_ADD_430_U129); 
assign P3_ADD_430_U98 = ~P3_ADD_430_U14; 
assign P3_ADD_430_U127 = ~(P3_ADD_430_U14 & P3_REIP_REG_7__SCAN_IN); 
assign P3_ADD_380_U69 = ~(P3_ADD_380_U137 & P3_ADD_380_U136); 
assign P3_ADD_380_U102 = ~P3_ADD_380_U15; 
assign P3_ADD_380_U134 = ~(P3_ADD_380_U15 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_GTE_370_U7 = P3_SUB_370_U21 & P3_GTE_370_U9; 
assign P3_ADD_344_U69 = ~(P3_ADD_344_U137 & P3_ADD_344_U136); 
assign P3_ADD_344_U102 = ~P3_ADD_344_U15; 
assign P3_ADD_344_U134 = ~(P3_ADD_344_U15 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_339_U65 = ~(P3_ADD_339_U130 & P3_ADD_339_U129); 
assign P3_ADD_339_U98 = ~P3_ADD_339_U14; 
assign P3_ADD_339_U127 = ~(P3_ADD_339_U14 & P3_PHYADDRPOINTER_REG_7__SCAN_IN); 
assign P3_LT_589_U7 = P3_SUB_589_U7 & P3_SUB_589_U6; 
assign P3_ADD_541_U65 = ~(P3_ADD_541_U130 & P3_ADD_541_U129); 
assign P3_ADD_541_U98 = ~P3_ADD_541_U14; 
assign P3_ADD_541_U127 = ~(P3_ADD_541_U14 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_SUB_355_U16 = ~(P3_SUB_355_U41 & P3_SUB_355_U40); 
assign P3_SUB_355_U55 = ~(P3_SUB_355_U38 & P3_SUB_355_U54); 
assign P3_SUB_450_U14 = ~(P3_SUB_450_U39 & P3_SUB_450_U38); 
assign P3_SUB_450_U52 = ~(P3_SUB_450_U36 & P3_SUB_450_U51); 
assign P3_SUB_485_U14 = ~(P3_SUB_485_U39 & P3_SUB_485_U38); 
assign P3_SUB_485_U52 = ~(P3_SUB_485_U36 & P3_SUB_485_U51); 
assign P3_ADD_515_U65 = ~(P3_ADD_515_U130 & P3_ADD_515_U129); 
assign P3_ADD_515_U98 = ~P3_ADD_515_U14; 
assign P3_ADD_515_U127 = ~(P3_ADD_515_U14 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_394_U66 = ~(P3_ADD_394_U134 & P3_ADD_394_U133); 
assign P3_ADD_394_U101 = ~P3_ADD_394_U14; 
assign P3_ADD_394_U131 = ~(P3_ADD_394_U14 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_SUB_414_U53 = P3_SUB_414_U129 & P3_SUB_414_U128; 
assign P3_SUB_414_U93 = ~P3_SUB_414_U28; 
assign P3_SUB_414_U126 = ~(P3_SUB_414_U125 & P3_EBX_REG_10__SCAN_IN); 
assign P3_SUB_414_U158 = ~(P3_SUB_414_U28 & P3_EBX_REG_11__SCAN_IN); 
assign P3_ADD_441_U65 = ~(P3_ADD_441_U130 & P3_ADD_441_U129); 
assign P3_ADD_441_U98 = ~P3_ADD_441_U14; 
assign P3_ADD_441_U127 = ~(P3_ADD_441_U14 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_349_U69 = ~(P3_ADD_349_U137 & P3_ADD_349_U136); 
assign P3_ADD_349_U102 = ~P3_ADD_349_U15; 
assign P3_ADD_349_U134 = ~(P3_ADD_349_U15 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_405_U66 = ~(P3_ADD_405_U134 & P3_ADD_405_U133); 
assign P3_ADD_405_U101 = ~P3_ADD_405_U14; 
assign P3_ADD_405_U131 = ~(P3_ADD_405_U14 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_553_U69 = ~(P3_ADD_553_U137 & P3_ADD_553_U136); 
assign P3_ADD_553_U102 = ~P3_ADD_553_U15; 
assign P3_ADD_553_U134 = ~(P3_ADD_553_U15 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_558_U69 = ~(P3_ADD_558_U137 & P3_ADD_558_U136); 
assign P3_ADD_558_U102 = ~P3_ADD_558_U15; 
assign P3_ADD_558_U134 = ~(P3_ADD_558_U15 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_385_U69 = ~(P3_ADD_385_U137 & P3_ADD_385_U136); 
assign P3_ADD_385_U102 = ~P3_ADD_385_U15; 
assign P3_ADD_385_U134 = ~(P3_ADD_385_U15 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_547_U69 = ~(P3_ADD_547_U137 & P3_ADD_547_U136); 
assign P3_ADD_547_U102 = ~P3_ADD_547_U15; 
assign P3_ADD_547_U134 = ~(P3_ADD_547_U15 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_SUB_412_U14 = ~(P3_SUB_412_U39 & P3_SUB_412_U38); 
assign P3_SUB_412_U52 = ~(P3_SUB_412_U36 & P3_SUB_412_U51); 
assign P3_SUB_504_U14 = ~(P3_SUB_504_U39 & P3_SUB_504_U38); 
assign P3_SUB_504_U52 = ~(P3_SUB_504_U36 & P3_SUB_504_U51); 
assign P3_SUB_401_U16 = ~(P3_SUB_401_U41 & P3_SUB_401_U40); 
assign P3_SUB_401_U55 = ~(P3_SUB_401_U38 & P3_SUB_401_U54); 
assign P3_SUB_390_U16 = ~(P3_SUB_390_U41 & P3_SUB_390_U40); 
assign P3_SUB_390_U55 = ~(P3_SUB_390_U38 & P3_SUB_390_U54); 
assign P3_ADD_494_U65 = ~(P3_ADD_494_U130 & P3_ADD_494_U129); 
assign P3_ADD_494_U98 = ~P3_ADD_494_U14; 
assign P3_ADD_494_U127 = ~(P3_ADD_494_U14 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_536_U65 = ~(P3_ADD_536_U130 & P3_ADD_536_U129); 
assign P3_ADD_536_U98 = ~P3_ADD_536_U14; 
assign P3_ADD_536_U127 = ~(P3_ADD_536_U14 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_402_1132_U4 = ~P3_U2613; 
assign P3_ADD_402_1132_U7 = ~P3_U2614; 
assign P3_ADD_402_1132_U9 = ~P3_U2615; 
assign P3_ADD_402_1132_U11 = ~P3_U2616; 
assign P3_ADD_402_1132_U13 = ~P3_U2617; 
assign P3_ADD_402_1132_U15 = ~P3_U2618; 
assign P3_ADD_402_1132_U17 = ~P3_U2619; 
assign P3_ADD_402_1132_U26 = ~P3_U2620; 
assign P2_R2182_U22 = ~P2_U2675; 
assign P2_R2182_U24 = ~P2_U2676; 
assign P2_R2182_U35 = ~P2_U2674; 
assign P2_R2182_U43 = ~P2_U2679; 
assign P2_R2182_U47 = ~P2_U2680; 
assign P2_R2182_U49 = ~P2_U2678; 
assign P2_R2182_U51 = ~P2_U2677; 
assign P2_R2182_U53 = ~P2_U2665; 
assign P2_R2182_U55 = ~P2_U2664; 
assign P2_R2182_U57 = ~P2_U2663; 
assign P2_R2182_U59 = ~P2_U2662; 
assign P2_R2182_U61 = ~P2_U2661; 
assign P2_R2182_U63 = ~P2_U2660; 
assign P2_R2182_U65 = ~P2_U2659; 
assign P2_R2182_U107 = ~P2_U2658; 
assign P2_R2027_U69 = ~(P2_R2027_U137 & P2_R2027_U136); 
assign P2_R2027_U102 = ~P2_R2027_U15; 
assign P2_R2027_U134 = ~(P2_R2027_U15 & P2_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P2_R2337_U63 = ~(P2_R2337_U128 & P2_R2337_U127); 
assign P2_R2337_U99 = ~P2_R2337_U15; 
assign P2_R2337_U125 = ~(P2_R2337_U15 & P2_PHYADDRPOINTER_REG_8__SCAN_IN); 
assign P2_R2147_U16 = ~(P2_R2147_U13 & P2_R2147_U10); 
assign P2_R2238_U16 = ~(P2_R2238_U41 & P2_R2238_U40); 
assign P2_R2238_U55 = ~(P2_R2238_U38 & P2_R2238_U54); 
assign P2_R1957_U18 = P2_R1957_U92 & P2_R1957_U22; 
assign P2_R1957_U89 = ~(P2_R1957_U84 & P2_R1957_U56); 
assign P2_R1957_U133 = ~(P2_R1957_U84 & P2_R1957_U56); 
assign P2_SUB_450_U14 = ~(P2_SUB_450_U39 & P2_SUB_450_U38); 
assign P2_SUB_450_U52 = ~(P2_SUB_450_U36 & P2_SUB_450_U51); 
assign P2_ADD_394_U63 = ~(P2_ADD_394_U128 & P2_ADD_394_U127); 
assign P2_ADD_394_U101 = ~P2_ADD_394_U14; 
assign P2_ADD_394_U181 = ~(P2_ADD_394_U14 & P2_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P1_R2027_U51 = ~(P1_R2027_U142 & P1_R2027_U141); 
assign P1_R2027_U52 = ~(P1_R2027_U144 & P1_R2027_U143); 
assign P1_R2027_U113 = ~P1_R2027_U22; 
assign P1_R2027_U140 = ~P1_R2027_U110; 
assign P1_R2027_U200 = ~(P1_R2027_U22 & P1_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P1_R2027_U201 = ~(P1_R2027_U110 & P1_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P1_R2099_U5 = ~P1_U4189; 
assign P1_R2099_U6 = ~P1_U2678; 
assign P1_R2099_U146 = P1_U4190 | P1_U4189; 
assign P1_R2099_U148 = ~(P1_U4189 & P1_U4190); 
assign P1_R2099_U345 = ~(P1_U4189 & P1_R2099_U4); 
assign P1_R2167_U23 = ~P1_U2722; 
assign P1_R2337_U65 = ~(P1_R2337_U130 & P1_R2337_U129); 
assign P1_R2337_U98 = ~P1_R2337_U14; 
assign P1_R2337_U127 = ~(P1_R2337_U14 & P1_PHYADDRPOINTER_REG_7__SCAN_IN); 
assign P1_R2096_U65 = ~(P1_R2096_U130 & P1_R2096_U129); 
assign P1_R2096_U98 = ~P1_R2096_U14; 
assign P1_R2096_U127 = ~(P1_R2096_U14 & P1_REIP_REG_7__SCAN_IN); 
assign P1_R2238_U16 = ~(P1_R2238_U41 & P1_R2238_U40); 
assign P1_R2238_U55 = ~(P1_R2238_U38 & P1_R2238_U54); 
assign P1_SUB_450_U16 = ~(P1_SUB_450_U41 & P1_SUB_450_U40); 
assign P1_SUB_450_U55 = ~(P1_SUB_450_U38 & P1_SUB_450_U54); 
assign P1_ADD_405_U63 = ~(P1_ADD_405_U128 & P1_ADD_405_U127); 
assign P1_ADD_405_U101 = ~P1_ADD_405_U14; 
assign P1_ADD_405_U181 = ~(P1_ADD_405_U14 & P1_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P1_ADD_515_U62 = ~(P1_ADD_515_U124 & P1_ADD_515_U123); 
assign P1_ADD_515_U98 = ~P1_ADD_515_U14; 
assign P1_ADD_515_U177 = ~(P1_ADD_515_U14 & P1_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_U2363 = P3_U5442 & P3_U5435; 
assign P3_U2364 = P3_U5392 & P3_U3204; 
assign P3_U2365 = P3_U5341 & P3_U3201; 
assign P3_U2366 = P3_U5290 & P3_U3198; 
assign P3_U2367 = P3_U5239 & P3_U5232; 
assign P3_U2449 = P3_U4344 & P3_U4522; 
assign P3_U2452 = P3_U2463 & P3_U4522 & P3_U2412; 
assign P3_U2487 = P3_U3270 & P3_U3142; 
assign P3_U2493 = P3_U4646 & P3_U3128; 
assign P3_U2495 = P3_U4646 & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN; 
assign P3_U2514 = P3_U3218 & P3_U3216; 
assign P3_U2605 = ~(P3_U4215 & P3_U4214 & P3_U4213 & P3_U4212); 
assign P3_U2606 = ~(P3_U4211 & P3_U4210 & P3_U4209 & P3_U4208); 
assign P3_U2607 = ~(P3_U4207 & P3_U4206 & P3_U4205 & P3_U4204); 
assign P3_U2608 = ~(P3_U4203 & P3_U4202 & P3_U4201 & P3_U4200); 
assign P3_U2609 = ~(P3_U4199 & P3_U4198 & P3_U4197 & P3_U4196); 
assign P3_U2610 = ~(P3_U4195 & P3_U4194 & P3_U4193 & P3_U4192); 
assign P3_U2611 = ~(P3_U4191 & P3_U4190 & P3_U4189 & P3_U4188); 
assign P3_U2612 = ~(P3_U4187 & P3_U4186 & P3_U4185 & P3_U4184); 
assign P3_U2621 = ~(P3_U4183 & P3_U4182 & P3_U4181 & P3_U4180); 
assign P3_U2622 = ~(P3_U4179 & P3_U4178 & P3_U4177 & P3_U4176); 
assign P3_U2623 = ~(P3_U4175 & P3_U4174 & P3_U4173 & P3_U4172); 
assign P3_U2624 = ~(P3_U4171 & P3_U4170 & P3_U4169 & P3_U4168); 
assign P3_U2625 = ~(P3_U4167 & P3_U4166 & P3_U4165 & P3_U4164); 
assign P3_U2626 = ~(P3_U4163 & P3_U4162 & P3_U4161 & P3_U4160); 
assign P3_U2627 = ~(P3_U4159 & P3_U4158 & P3_U4157 & P3_U4156); 
assign P3_U2628 = ~(P3_U4155 & P3_U4154 & P3_U4153 & P3_U4152); 
assign P3_U3062 = ~(P3_U4247 & P3_U4246 & P3_U4245 & P3_U4244); 
assign P3_U3063 = ~(P3_U4243 & P3_U4242 & P3_U4241 & P3_U4240); 
assign P3_U3064 = ~(P3_U4239 & P3_U4238 & P3_U4237 & P3_U4236); 
assign P3_U3065 = ~(P3_U4235 & P3_U4234 & P3_U4233 & P3_U4232); 
assign P3_U3066 = ~(P3_U4231 & P3_U4230 & P3_U4229 & P3_U4228); 
assign P3_U3067 = ~(P3_U4227 & P3_U4226 & P3_U4225 & P3_U4224); 
assign P3_U3068 = ~(P3_U4223 & P3_U4222 & P3_U4221 & P3_U4220); 
assign P3_U3069 = ~(P3_U4219 & P3_U4218 & P3_U4217 & P3_U4216); 
assign P3_U3165 = ~(P3_U7965 & P3_U3142); 
assign P3_U3219 = ~(P3_U3662 & P3_U2461); 
assign P3_U3655 = P3_U3107 & P3_U3118; 
assign P3_U3661 = P3_U2461 & P3_U4297; 
assign P3_U3673 = P3_U4505 & P3_U2456; 
assign P3_U3691 = P3_U2456 & P3_U4590; 
assign P3_U4296 = ~P3_U3112; 
assign P3_U4323 = ~P3_U3114; 
assign P3_U4324 = ~P3_U3118; 
assign P3_U4348 = ~P3_U3236; 
assign P3_U4350 = ~P3_U3208; 
assign P3_U4351 = ~P3_U3216; 
assign P3_U4608 = ~P3_U3113; 
assign P3_U4621 = ~(P3_U3359 & P3_U7916); 
assign P3_U4647 = ~P3_U3143; 
assign P3_U4656 = ~P3_U3142; 
assign P3_U4659 = ~(P3_U3140 & P3_U3142); 
assign P3_U5078 = ~P3_U3185; 
assign P3_U5129 = ~P3_U3189; 
assign P3_U5181 = ~P3_U3193; 
assign P3_U5283 = ~P3_U3198; 
assign P3_U5334 = ~P3_U3201; 
assign P3_U5385 = ~P3_U3204; 
assign P3_U5510 = ~(P3_U7974 & P3_U7973 & P3_U3104); 
assign P3_U5515 = ~(P3_U5514 & P3_U3216 & P3_U4556); 
assign P3_U5517 = ~(P3_U4488 & P3_U5516); 
assign P3_U5518 = ~(P3_U3103 & P3_U3218 & P3_U3112); 
assign P3_U5523 = ~(P3_U3111 & P3_U3114); 
assign P3_U5587 = ~(P3_U5582 & P3_U3142); 
assign P3_U5602 = ~(P3_U5601 & P3_U5600); 
assign P3_U7376 = ~(P3_U3112 & P3_U3118); 
assign P3_U7385 = ~(P3_U3111 & P3_U3114 & P3_STATE2_REG_2__SCAN_IN); 
assign P3_U7968 = ~P3_U3271; 
assign P3_U7978 = ~(P3_U5513 & P3_U3107 & P3_U4590); 
assign P3_U7998 = ~(P3_U3271 & P3_U3143); 
assign P2_U2599 = ~(P2_U4258 & P2_U4257 & P2_U4256 & P2_U4255); 
assign P2_U2600 = ~(P2_U4254 & P2_U4253 & P2_U4252 & P2_U4251); 
assign P2_U2601 = ~(P2_U4250 & P2_U4249 & P2_U4248 & P2_U4247); 
assign P2_U2602 = ~(P2_U4246 & P2_U4245 & P2_U4244 & P2_U4243); 
assign P2_U2603 = ~(P2_U4242 & P2_U4241 & P2_U4240 & P2_U4239); 
assign P2_U2604 = ~(P2_U4238 & P2_U4237 & P2_U4236 & P2_U4235); 
assign P2_U2605 = ~(P2_U4234 & P2_U4233 & P2_U4232 & P2_U4231); 
assign P2_U2606 = ~(P2_U4230 & P2_U4229 & P2_U4228 & P2_U4227); 
assign P2_U2650 = P2_U2352 & P2_U3242; 
assign P2_U2651 = P2_U2352 & P2_U7217; 
assign P2_U2652 = P2_U2352 & P2_U7251; 
assign P2_U2653 = P2_U2352 & P2_U7285; 
assign P2_U2666 = P2_U2614 & P2_U2355; 
assign P2_U2667 = P2_U2613 & P2_U2355; 
assign P2_U2668 = P2_U2612 & P2_U2355; 
assign P2_U2669 = P2_U2611 & P2_U2355; 
assign P2_U2670 = P2_U2610 & P2_U2355; 
assign P2_U2671 = P2_U2609 & P2_U2355; 
assign P2_U2672 = P2_U2608 & P2_U2355; 
assign P2_U2673 = P2_U2607 & P2_U2355; 
assign P2_U2705 = ~(P2_U4390 & P2_U7730); 
assign P2_U2706 = ~(P2_U7732 & P2_U7733 & P2_U3550); 
assign P2_U2758 = P2_U4428 & P2_U3242; 
assign P2_U2759 = P2_U4428 & P2_U7217; 
assign P2_U2760 = P2_U4428 & P2_U7251; 
assign P2_U3254 = ~(P2_U2590 & P2_U4429); 
assign P2_U3296 = ~(P2_U2451 & P2_U4428); 
assign P2_U3522 = ~(P2_U2451 & P2_U4429); 
assign P2_U3549 = ~(P2_U2356 & P2_U4420); 
assign P2_U3554 = ~(P2_U4415 & P2_U3576); 
assign P2_U3572 = ~P2_U3242; 
assign P2_U3578 = ~(P2_U2590 & P2_U4428); 
assign P2_U3651 = ~(P2_U8358 & P2_U8357); 
assign P2_U3652 = ~(P2_U8360 & P2_U8359); 
assign P2_U3713 = P2_U4599 & P2_U4598; 
assign P2_U3869 = P2_U3868 & P2_U5576; 
assign P2_U3877 = P2_U7859 & P2_U5593; 
assign P2_U4338 = P2_U7425 & P2_U4413; 
assign P2_U4342 = P2_U4413 & P2_U4341; 
assign P2_U4346 = P2_U7442 & P2_U7443; 
assign P2_U4347 = P2_U7445 & P2_U7446; 
assign P2_U4348 = P2_U7448 & P2_U7449; 
assign P2_U4349 = P2_U7451 & P2_U7452; 
assign P2_U4350 = P2_U7454 & P2_U7455; 
assign P2_U4351 = P2_U7457 & P2_U7458; 
assign P2_U4352 = P2_U7460 & P2_U7461; 
assign P2_U4353 = P2_U7463 & P2_U7464; 
assign P2_U4354 = P2_U7466 & P2_U7467; 
assign P2_U4355 = P2_U7469 & P2_U7470; 
assign P2_U4356 = P2_U7472 & P2_U7473; 
assign P2_U4357 = P2_U7475 & P2_U7476; 
assign P2_U4358 = P2_U7478 & P2_U7479; 
assign P2_U4359 = P2_U7481 & P2_U7482; 
assign P2_U4360 = P2_U7484 & P2_U7485; 
assign P2_U4361 = P2_U7487 & P2_U7488; 
assign P2_U4362 = P2_U7490 & P2_U7491; 
assign P2_U4363 = P2_U7493 & P2_U7494; 
assign P2_U4364 = P2_U7496 & P2_U7497; 
assign P2_U4365 = P2_U7499 & P2_U7500; 
assign P2_U4366 = P2_U7502 & P2_U7503; 
assign P2_U4367 = P2_U7505 & P2_U7506; 
assign P2_U4374 = P2_U7532 & P2_U7533; 
assign P2_U4375 = P2_U7536 & P2_U7535; 
assign P2_U4383 = P2_U7579 & P2_U4422; 
assign P2_U4416 = ~P2_U3576; 
assign P2_U4418 = ~P2_U3550; 
assign P2_U4421 = ~P2_U3539; 
assign P2_U4424 = ~P2_U3282; 
assign P2_U4437 = ~(P2_U3875 & P2_U2376); 
assign P2_U4459 = ~P2_U3575; 
assign P2_U4470 = ~(P2_U3876 & P2_U2376); 
assign P2_U4475 = ~P2_U3293; 
assign P2_U5589 = ~(P2_U8075 & P2_U8074 & P2_U3879); 
assign P2_U5594 = ~(P2_U5592 & P2_U2616); 
assign P2_U5625 = ~(P2_U7882 & P2_U5624); 
assign P2_U5674 = ~(P2_U4427 & P2_U4420); 
assign P2_U7422 = ~(P2_U2352 & P2_U7319); 
assign P2_U7424 = ~(P2_U2352 & P2_U7353); 
assign P2_U7427 = ~(P2_U2352 & P2_U7387); 
assign P2_U7429 = ~(P2_U2352 & P2_U7421); 
assign P2_U7432 = ~(P2_U4414 & P2_U7431 & P2_U4413); 
assign P2_U7436 = ~(P2_U2352 & P2_U2608); 
assign P2_U7440 = ~(P2_U2352 & P2_U2607); 
assign P2_U7510 = ~(P2_U2352 & P2_U2614); 
assign P2_U7514 = ~(P2_U2352 & P2_U2613); 
assign P2_U7518 = ~(P2_U2352 & P2_U2612); 
assign P2_U7522 = ~(P2_U2352 & P2_U2611); 
assign P2_U7526 = ~(P2_U2352 & P2_U2610); 
assign P2_U7530 = ~(P2_U2352 & P2_U2609); 
assign P2_U7561 = ~(P2_U4596 & P2_U3294); 
assign P2_U7562 = ~(P2_U4428 & P2_U7285); 
assign P2_U7564 = ~(P2_U4428 & P2_U7319); 
assign P2_U7566 = ~(P2_U4428 & P2_U7353); 
assign P2_U7568 = ~(P2_U4428 & P2_U7387); 
assign P2_U7570 = ~(P2_U4428 & P2_U7421); 
assign P2_U7577 = ~(P2_U4377 & P2_U5572); 
assign P2_U7580 = ~(P2_U4376 & P2_U5592); 
assign P2_U7589 = ~(P2_U2590 & P2_U6845); 
assign P2_U7723 = ~(P2_U3550 & P2_U3536); 
assign P2_U7884 = ~(P2_U4596 & P2_U7883); 
assign P2_U8052 = ~(P2_U7871 & P2_U3293); 
assign P2_U8053 = ~(P2_U3253 & P2_U3282); 
assign P2_U8069 = ~(P2_U3280 & P2_U5575); 
assign P2_U8095 = ~(P2_U3886 & P2_U4597 & P2_U3255); 
assign P2_U8122 = ~(P2_U2616 & P2_U3282); 
assign P2_U8297 = ~(P2_U3242 & P2_U7873); 
assign P2_U8299 = ~(P2_U7217 & P2_U7873); 
assign P2_U8301 = ~(P2_U7251 & P2_U7873); 
assign P2_U8303 = ~(P2_U7285 & P2_U7873); 
assign P2_U8305 = ~(P2_U7319 & P2_U7873); 
assign P2_U8307 = ~(P2_U7353 & P2_U7873); 
assign P2_U8309 = ~(P2_U7387 & P2_U7873); 
assign P2_U8311 = ~(P2_U7421 & P2_U7873); 
assign P2_U8347 = ~(P2_U3255 & P2_U7740); 
assign P2_U8365 = ~(P2_R2337_U63 & P2_U3284); 
assign P1_U2355 = P1_U3234 & P1_U2450; 
assign P1_U2679 = ~(P1_U7405 & P1_U7404); 
assign P1_U2680 = ~(P1_U7407 & P1_U7406); 
assign P1_U2681 = ~(P1_U7411 & P1_U7410); 
assign P1_U2682 = ~(P1_U7413 & P1_U7412); 
assign P1_U2683 = ~(P1_U7415 & P1_U7414); 
assign P1_U2684 = ~(P1_U7417 & P1_U7416); 
assign P1_U2685 = ~(P1_U7419 & P1_U7418); 
assign P1_U2686 = ~(P1_U7421 & P1_U7420); 
assign P1_U2687 = ~(P1_U7423 & P1_U7422); 
assign P1_U2688 = ~(P1_U7425 & P1_U7424); 
assign P1_U2689 = ~(P1_U7427 & P1_U7426); 
assign P1_U2690 = ~(P1_U7429 & P1_U7428); 
assign P1_U2691 = ~(P1_U7433 & P1_U7432); 
assign P1_U2692 = ~(P1_U7435 & P1_U7434); 
assign P1_U2693 = ~(P1_U7437 & P1_U7436); 
assign P1_U2694 = ~(P1_U7439 & P1_U7438); 
assign P1_U2695 = ~(P1_U7441 & P1_U7440); 
assign P1_U2696 = ~(P1_U7443 & P1_U7442); 
assign P1_U2697 = ~(P1_U7445 & P1_U7444); 
assign P1_U2698 = ~(P1_U7447 & P1_U7446); 
assign P1_U2699 = ~(P1_U7449 & P1_U7448); 
assign P1_U2700 = ~(P1_U7451 & P1_U7450); 
assign P1_U2701 = ~(P1_U7393 & P1_U7392); 
assign P1_U2702 = ~(P1_U7395 & P1_U7394); 
assign P1_U2703 = ~(P1_U7397 & P1_U7396); 
assign P1_U2704 = ~(P1_U7399 & P1_U7398); 
assign P1_U2705 = ~(P1_U7401 & P1_U7400); 
assign P1_U2706 = ~(P1_U7403 & P1_U7402); 
assign P1_U2707 = ~(P1_U7409 & P1_U7408); 
assign P1_U2708 = ~(P1_U7431 & P1_U7430); 
assign P1_U2709 = ~(P1_U7453 & P1_U7452); 
assign P1_U2710 = ~(P1_U7455 & P1_U7454); 
assign P1_U2714 = ~(P1_U7386 & P1_U7385 & P1_U4166 & P1_U3434); 
assign P1_U3245 = ~(P1_U7086 & P1_U5464); 
assign P1_U3292 = ~(P1_U4256 & P1_U2431); 
assign P1_U3441 = ~P1_U3234; 
assign P1_U3446 = ~(P1_U4197 & P1_U4234); 
assign P1_U3742 = P1_U5496 & P1_U3393; 
assign P1_U3743 = P1_U5498 & P1_U5497; 
assign P1_U3745 = P1_U4263 & P1_U3397; 
assign P1_U4006 = P1_U6760 & P1_U4007; 
assign P1_U4008 = P1_U6764 & P1_U6765; 
assign P1_U4010 = P1_U6776 & P1_U6777; 
assign P1_U4021 = P1_U6821 & P1_U6822; 
assign P1_U4027 = P1_U6860 & P1_U6861; 
assign P1_U4067 = P1_U4256 & P1_STATE2_REG_0__SCAN_IN; 
assign P1_U4111 = P1_U7089 & P1_U3427; 
assign P1_U4158 = P1_U4157 & P1_U7360; 
assign P1_U4162 = P1_U7371 & P1_U2603; 
assign P1_U4165 = P1_U7382 & P1_U7383; 
assign P1_U4193 = ~P1_U3434; 
assign P1_U4194 = ~P1_U3420; 
assign P1_U4202 = ~P1_U3428; 
assign P1_U4204 = ~P1_U3427; 
assign P1_U4205 = ~(P1_U3885 & P1_U4189 & P1_U4197); 
assign P1_U4212 = ~P1_U3447; 
assign P1_U4213 = ~P1_U3448; 
assign P1_U4214 = ~P1_U3400; 
assign P1_U4215 = ~P1_U3288; 
assign P1_U4217 = ~(P1_U3578 & P1_U2431); 
assign P1_U4218 = ~P1_U3399; 
assign P1_U4266 = ~P1_U3410; 
assign P1_U4505 = ~(P1_U4504 & P1_U3579); 
assign P1_U5466 = ~(P1_U5465 & P1_U3283 & P1_U5464); 
assign P1_U5520 = ~(P1_U2431 & P1_U4249); 
assign P1_U5565 = ~(P1_U4262 & P1_U4208); 
assign P1_U5566 = ~(P1_U4256 & P1_U2389); 
assign P1_U5568 = ~(P1_U4264 & P1_U4494); 
assign P1_U6606 = ~(P1_U3964 & P1_U6605); 
assign P1_U6758 = ~(P1_R2337_U65 & P1_U2352); 
assign P1_U6908 = ~(P1_U4032 & P1_U4031 & P1_U4030 & P1_U4029); 
assign P1_U6926 = ~(P1_U4036 & P1_U4035 & P1_U4034 & P1_U4033); 
assign P1_U6957 = ~(P1_U4040 & P1_U4039 & P1_U4038 & P1_U4037); 
assign P1_U6974 = ~(P1_U4044 & P1_U4043 & P1_U4042 & P1_U4041); 
assign P1_U6991 = ~(P1_U4048 & P1_U4047 & P1_U4046 & P1_U4045); 
assign P1_U7023 = ~(P1_U4056 & P1_U4055 & P1_U4054 & P1_U4053); 
assign P1_U7040 = ~(P1_U4060 & P1_U4059 & P1_U4058 & P1_U4057); 
assign P1_U7047 = ~(P1_U4206 & P1_U3234); 
assign P1_U7049 = ~(P1_U4206 & P1_U3233); 
assign P1_U7051 = ~(P1_U4206 & P1_U3232); 
assign P1_U7053 = ~(P1_U4206 & P1_U3231); 
assign P1_U7054 = ~(P1_U4206 & P1_U3230); 
assign P1_U7056 = ~(P1_U4206 & P1_U3229); 
assign P1_U7058 = ~(P1_U4206 & P1_U3228); 
assign P1_U7060 = ~(P1_U4206 & P1_U3227); 
assign P1_U7061 = ~(P1_U3234 & P1_U4400); 
assign P1_U7063 = ~(P1_U3428 & P1_U3427); 
assign P1_U7085 = ~(P1_U7084 & P1_U3422); 
assign P1_U7236 = ~(P1_U4124 & P1_U4123 & P1_U4122 & P1_U4121); 
assign P1_U7253 = ~(P1_U4128 & P1_U4127 & P1_U4126 & P1_U4125); 
assign P1_U7270 = ~(P1_U4132 & P1_U4131 & P1_U4130 & P1_U4129); 
assign P1_U7302 = ~(P1_U4140 & P1_U4139 & P1_U4138 & P1_U4137); 
assign P1_U7319 = ~(P1_U4144 & P1_U4143 & P1_U4142 & P1_U4141); 
assign P1_U7336 = ~(P1_U4148 & P1_U4147 & P1_U4146 & P1_U4145); 
assign P1_U7353 = ~(P1_U4152 & P1_U4151 & P1_U4150 & P1_U4149); 
assign P1_U7356 = ~(P1_U3396 & P1_U3410); 
assign P1_U7363 = ~(P1_U3420 & P1_U3434 & P1_U4195 & P1_U7362 & P1_U7361); 
assign P1_U7381 = ~(P1_U3420 & P1_U7380); 
assign P1_U7471 = ~(P1_U7084 & P1_U3422); 
assign P1_U7476 = ~(P1_U4264 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U7496 = ~(P1_U3734 & P1_U7493); 
assign P1_U7507 = ~(P1_U3759 & P1_U7493); 
assign P1_U7605 = ~(P1_U3867 & P1_U7493); 
assign P1_U7607 = ~(P1_U4208 & P1_U7493); 
assign P1_U7609 = ~(P1_U3279 & P1_U3400); 
assign P1_U7610 = ~(P1_U3754 & P1_U7493); 
assign P1_U7615 = ~(P1_U4052 & P1_U4051 & P1_U4050 & P1_U4049); 
assign P1_U7620 = ~(P1_U4136 & P1_U4135 & P1_U4134 & P1_U4133); 
assign P1_U7629 = ~P1_U3392; 
assign P1_U7632 = ~(P1_U7631 & P1_U7630); 
assign P3_ADD_526_U25 = ~(P3_ADD_526_U86 & P3_ADD_526_U113); 
assign P3_ADD_526_U109 = ~(P3_ADD_526_U113 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_526_U199 = ~(P3_ADD_526_U113 & P3_ADD_526_U21); 
assign P3_ADD_526_U202 = ~(P3_ADD_526_U140 & P3_ADD_526_U19); 
assign P3_ADD_552_U25 = ~(P3_ADD_552_U86 & P3_ADD_552_U113); 
assign P3_ADD_552_U109 = ~(P3_ADD_552_U113 & P3_EBX_REG_11__SCAN_IN); 
assign P3_ADD_552_U199 = ~(P3_ADD_552_U113 & P3_ADD_552_U21); 
assign P3_ADD_552_U202 = ~(P3_ADD_552_U140 & P3_ADD_552_U19); 
assign P3_ADD_546_U25 = ~(P3_ADD_546_U86 & P3_ADD_546_U113); 
assign P3_ADD_546_U109 = ~(P3_ADD_546_U113 & P3_EAX_REG_11__SCAN_IN); 
assign P3_ADD_546_U199 = ~(P3_ADD_546_U113 & P3_ADD_546_U21); 
assign P3_ADD_546_U202 = ~(P3_ADD_546_U140 & P3_ADD_546_U19); 
assign P3_ADD_476_U16 = ~(P3_ADD_476_U98 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_476_U128 = ~(P3_ADD_476_U98 & P3_ADD_476_U15); 
assign P3_ADD_531_U17 = ~(P3_ADD_531_U102 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_531_U135 = ~(P3_ADD_531_U102 & P3_ADD_531_U16); 
assign P3_SUB_320_U26 = ~P3_ADD_318_U65; 
assign P3_SUB_320_U57 = P3_SUB_320_U133 & P3_SUB_320_U132; 
assign P3_SUB_320_U90 = ~(P3_ADD_318_U65 & P3_SUB_320_U89); 
assign P3_ADD_318_U16 = ~(P3_ADD_318_U98 & P3_PHYADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_318_U128 = ~(P3_ADD_318_U98 & P3_ADD_318_U15); 
assign P3_SUB_370_U20 = ~(P3_SUB_370_U56 & P3_SUB_370_U55); 
assign P3_SUB_370_U42 = ~P3_SUB_370_U16; 
assign P3_SUB_370_U51 = ~(P3_SUB_370_U23 & P3_SUB_370_U16); 
assign P3_ADD_315_U17 = ~(P3_ADD_315_U95 & P3_PHYADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_315_U122 = ~(P3_ADD_315_U95 & P3_ADD_315_U15); 
assign P3_ADD_467_U16 = ~(P3_ADD_467_U98 & P3_REIP_REG_7__SCAN_IN); 
assign P3_ADD_467_U128 = ~(P3_ADD_467_U98 & P3_ADD_467_U15); 
assign P3_ADD_430_U16 = ~(P3_ADD_430_U98 & P3_REIP_REG_7__SCAN_IN); 
assign P3_ADD_430_U128 = ~(P3_ADD_430_U98 & P3_ADD_430_U15); 
assign P3_ADD_380_U17 = ~(P3_ADD_380_U102 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_380_U135 = ~(P3_ADD_380_U102 & P3_ADD_380_U16); 
assign P3_ADD_344_U17 = ~(P3_ADD_344_U102 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_344_U135 = ~(P3_ADD_344_U102 & P3_ADD_344_U16); 
assign P3_ADD_339_U16 = ~(P3_ADD_339_U98 & P3_PHYADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_339_U128 = ~(P3_ADD_339_U98 & P3_ADD_339_U15); 
assign P3_LT_589_U8 = ~(P3_LT_589_U7 | P3_SUB_589_U8 | P3_SUB_589_U9); 
assign P3_ADD_541_U16 = ~(P3_ADD_541_U98 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_541_U128 = ~(P3_ADD_541_U98 & P3_ADD_541_U15); 
assign P3_SUB_355_U20 = ~(P3_SUB_355_U56 & P3_SUB_355_U55); 
assign P3_SUB_355_U42 = ~P3_SUB_355_U16; 
assign P3_SUB_355_U51 = ~(P3_SUB_355_U23 & P3_SUB_355_U16); 
assign P3_SUB_450_U17 = ~(P3_SUB_450_U53 & P3_SUB_450_U52); 
assign P3_SUB_450_U40 = ~P3_SUB_450_U14; 
assign P3_SUB_450_U48 = ~(P3_SUB_450_U20 & P3_SUB_450_U14); 
assign P3_SUB_485_U17 = ~(P3_SUB_485_U53 & P3_SUB_485_U52); 
assign P3_SUB_485_U40 = ~P3_SUB_485_U14; 
assign P3_SUB_485_U48 = ~(P3_SUB_485_U20 & P3_SUB_485_U14); 
assign P3_ADD_515_U16 = ~(P3_ADD_515_U98 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_515_U128 = ~(P3_ADD_515_U98 & P3_ADD_515_U15); 
assign P3_ADD_394_U16 = ~(P3_ADD_394_U101 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_394_U132 = ~(P3_ADD_394_U101 & P3_ADD_394_U15); 
assign P3_SUB_414_U6 = P3_SUB_414_U126 & P3_SUB_414_U28; 
assign P3_SUB_414_U29 = ~(P3_SUB_414_U48 & P3_SUB_414_U81 & P3_SUB_414_U93); 
assign P3_SUB_414_U123 = ~(P3_SUB_414_U93 & P3_SUB_414_U81); 
assign P3_SUB_414_U159 = ~(P3_SUB_414_U93 & P3_SUB_414_U81); 
assign P3_ADD_441_U16 = ~(P3_ADD_441_U98 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_441_U128 = ~(P3_ADD_441_U98 & P3_ADD_441_U15); 
assign P3_ADD_349_U17 = ~(P3_ADD_349_U102 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_349_U135 = ~(P3_ADD_349_U102 & P3_ADD_349_U16); 
assign P3_ADD_405_U16 = ~(P3_ADD_405_U101 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_405_U132 = ~(P3_ADD_405_U101 & P3_ADD_405_U15); 
assign P3_ADD_553_U17 = ~(P3_ADD_553_U102 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_553_U135 = ~(P3_ADD_553_U102 & P3_ADD_553_U16); 
assign P3_ADD_558_U17 = ~(P3_ADD_558_U102 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_558_U135 = ~(P3_ADD_558_U102 & P3_ADD_558_U16); 
assign P3_ADD_385_U17 = ~(P3_ADD_385_U102 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_385_U135 = ~(P3_ADD_385_U102 & P3_ADD_385_U16); 
assign P3_ADD_547_U17 = ~(P3_ADD_547_U102 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_547_U135 = ~(P3_ADD_547_U102 & P3_ADD_547_U16); 
assign P3_SUB_412_U17 = ~(P3_SUB_412_U53 & P3_SUB_412_U52); 
assign P3_SUB_412_U40 = ~P3_SUB_412_U14; 
assign P3_SUB_412_U48 = ~(P3_SUB_412_U20 & P3_SUB_412_U14); 
assign P3_SUB_504_U17 = ~(P3_SUB_504_U53 & P3_SUB_504_U52); 
assign P3_SUB_504_U40 = ~P3_SUB_504_U14; 
assign P3_SUB_504_U48 = ~(P3_SUB_504_U20 & P3_SUB_504_U14); 
assign P3_SUB_401_U20 = ~(P3_SUB_401_U56 & P3_SUB_401_U55); 
assign P3_SUB_401_U42 = ~P3_SUB_401_U16; 
assign P3_SUB_401_U51 = ~(P3_SUB_401_U23 & P3_SUB_401_U16); 
assign P3_SUB_390_U20 = ~(P3_SUB_390_U56 & P3_SUB_390_U55); 
assign P3_SUB_390_U42 = ~P3_SUB_390_U16; 
assign P3_SUB_390_U51 = ~(P3_SUB_390_U23 & P3_SUB_390_U16); 
assign P3_ADD_494_U16 = ~(P3_ADD_494_U98 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_494_U128 = ~(P3_ADD_494_U98 & P3_ADD_494_U15); 
assign P3_ADD_536_U16 = ~(P3_ADD_536_U98 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_536_U128 = ~(P3_ADD_536_U98 & P3_ADD_536_U15); 
assign P2_R2182_U45 = ~P2_U2681; 
assign P2_R2027_U17 = ~(P2_R2027_U102 & P2_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P2_R2027_U135 = ~(P2_R2027_U102 & P2_R2027_U16); 
assign P2_R2337_U18 = ~(P2_R2337_U99 & P2_PHYADDRPOINTER_REG_8__SCAN_IN); 
assign P2_R2337_U126 = ~(P2_R2337_U99 & P2_R2337_U16); 
assign P2_R2147_U7 = ~(P2_R2147_U16 & P2_R2147_U15); 
assign P2_R2238_U20 = ~(P2_R2238_U56 & P2_R2238_U55); 
assign P2_R2238_U42 = ~P2_R2238_U16; 
assign P2_R2238_U51 = ~(P2_R2238_U23 & P2_R2238_U16); 
assign P2_R1957_U26 = ~P2_U3656; 
assign P2_R1957_U57 = P2_R1957_U133 & P2_R1957_U132; 
assign P2_R1957_U90 = ~(P2_U3656 & P2_R1957_U89); 
assign P2_SUB_450_U18 = ~(P2_SUB_450_U53 & P2_SUB_450_U52); 
assign P2_SUB_450_U40 = ~P2_SUB_450_U14; 
assign P2_SUB_450_U48 = ~(P2_SUB_450_U21 & P2_SUB_450_U14); 
assign P2_ADD_394_U16 = ~(P2_ADD_394_U101 & P2_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P2_ADD_394_U182 = ~(P2_ADD_394_U101 & P2_ADD_394_U15); 
assign P1_R2027_U25 = ~(P1_R2027_U86 & P1_R2027_U113); 
assign P1_R2027_U109 = ~(P1_R2027_U113 & P1_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P1_R2027_U199 = ~(P1_R2027_U113 & P1_R2027_U21); 
assign P1_R2027_U202 = ~(P1_R2027_U140 & P1_R2027_U19); 
assign P1_R2099_U346 = ~(P1_U4190 & P1_R2099_U5); 
assign P1_R2337_U16 = ~(P1_R2337_U98 & P1_PHYADDRPOINTER_REG_7__SCAN_IN); 
assign P1_R2337_U128 = ~(P1_R2337_U98 & P1_R2337_U15); 
assign P1_SUB_357_U6 = ~P1_U3233; 
assign P1_SUB_357_U7 = ~P1_U3228; 
assign P1_SUB_357_U8 = ~P1_U3234; 
assign P1_SUB_357_U9 = ~P1_U3232; 
assign P1_SUB_357_U10 = ~P1_U3227; 
assign P1_SUB_357_U11 = ~P1_U3230; 
assign P1_SUB_357_U12 = ~P1_U3229; 
assign P1_SUB_357_U13 = ~P1_U3231; 
assign P1_R2096_U16 = ~(P1_R2096_U98 & P1_REIP_REG_7__SCAN_IN); 
assign P1_R2096_U128 = ~(P1_R2096_U98 & P1_R2096_U15); 
assign P1_R2238_U20 = ~(P1_R2238_U56 & P1_R2238_U55); 
assign P1_R2238_U42 = ~P1_R2238_U16; 
assign P1_R2238_U51 = ~(P1_R2238_U23 & P1_R2238_U16); 
assign P1_SUB_450_U20 = ~(P1_SUB_450_U56 & P1_SUB_450_U55); 
assign P1_SUB_450_U42 = ~P1_SUB_450_U16; 
assign P1_SUB_450_U51 = ~(P1_SUB_450_U23 & P1_SUB_450_U16); 
assign P1_ADD_371_U4 = ~P1_U3227; 
assign P1_ADD_371_U7 = ~P1_U3228; 
assign P1_ADD_371_U8 = ~P1_U3230; 
assign P1_ADD_371_U10 = ~P1_U3231; 
assign P1_ADD_371_U12 = ~P1_U3232; 
assign P1_ADD_371_U13 = ~P1_U3233; 
assign P1_ADD_371_U15 = ~P1_U3229; 
assign P1_ADD_371_U16 = ~P1_U3234; 
assign P1_ADD_371_U22 = P1_U3234 & P1_U3233; 
assign P1_ADD_371_U26 = ~(P1_U3228 & P1_U3227); 
assign P1_ADD_371_U31 = ~(P1_U3228 & P1_U3227 & P1_U3229); 
assign P1_ADD_405_U16 = ~(P1_ADD_405_U101 & P1_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P1_ADD_405_U182 = ~(P1_ADD_405_U101 & P1_ADD_405_U15); 
assign P1_ADD_515_U16 = ~(P1_ADD_515_U98 & P1_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P1_ADD_515_U178 = ~(P1_ADD_515_U98 & P1_ADD_515_U15); 
assign P3_U2353 = P3_U3354 & P3_U2449; 
assign P3_U2450 = P3_U3660 & P3_U4351; 
assign P3_U2451 = P3_U4608 & P3_U3102 & P3_U2412; 
assign P3_U2462 = P3_U2412 & P3_U2449; 
assign P3_U2485 = P3_U4656 & P3_U3270; 
assign P3_U2488 = P3_U4657 & P3_U2487; 
assign P3_U2491 = P3_U4644 & P3_U2487; 
assign P3_U2494 = P3_U4645 & P3_U2487; 
assign P3_U2497 = P3_U2496 & P3_U2487; 
assign P3_U2509 = P3_U7965 & P3_U4656; 
assign P3_U3116 = ~(P3_U2452 & P3_U4297); 
assign P3_U3117 = ~(P3_U2452 & P3_U4296); 
assign P3_U3209 = ~(P3_U2514 & P3_U3113); 
assign P3_U3229 = ~(P3_U4323 & P3_U3218 & P3_U4350); 
assign P3_U3241 = ~P3_U2628; 
assign P3_U3355 = P3_U4323 & P3_U3101; 
assign P3_U3356 = P3_U4324 & P3_U3101; 
assign P3_U3361 = P3_U3235 & P3_U3236 & P3_U4621; 
assign P3_U3368 = P3_U3165 & P3_U4659; 
assign P3_U3664 = P3_U4573 & P3_U4324; 
assign P3_U3685 = P3_U5587 & P3_U5588; 
assign P3_U3688 = P3_U2456 & P3_U4296; 
assign P3_U3689 = P3_U2456 & P3_U4323; 
assign P3_U3690 = P3_U4608 & P3_U4556; 
assign P3_U4325 = ~P3_U3219; 
assign P3_U4333 = ~(P3_U4350 & P3_U3113); 
assign P3_U4339 = ~(P3_U3654 & P3_U4608); 
assign P3_U4658 = ~P3_U3165; 
assign P3_U4667 = ~(P3_U4657 & P3_U2487); 
assign P3_U4719 = ~(P3_U4644 & P3_U2487); 
assign P3_U4771 = ~(P3_U4645 & P3_U2487); 
assign P3_U4822 = ~(P3_U2496 & P3_U2487); 
assign P3_U5243 = ~(P3_U2367 & P3_U2420); 
assign P3_U5248 = ~(P3_U2367 & P3_U2419); 
assign P3_U5253 = ~(P3_U2367 & P3_U2418); 
assign P3_U5258 = ~(P3_U2367 & P3_U2417); 
assign P3_U5263 = ~(P3_U2367 & P3_U2416); 
assign P3_U5268 = ~(P3_U2367 & P3_U2415); 
assign P3_U5273 = ~(P3_U2367 & P3_U2414); 
assign P3_U5278 = ~(P3_U2367 & P3_U2413); 
assign P3_U5294 = ~(P3_U2366 & P3_U2420); 
assign P3_U5299 = ~(P3_U2366 & P3_U2419); 
assign P3_U5304 = ~(P3_U2366 & P3_U2418); 
assign P3_U5309 = ~(P3_U2366 & P3_U2417); 
assign P3_U5314 = ~(P3_U2366 & P3_U2416); 
assign P3_U5319 = ~(P3_U2366 & P3_U2415); 
assign P3_U5324 = ~(P3_U2366 & P3_U2414); 
assign P3_U5329 = ~(P3_U2366 & P3_U2413); 
assign P3_U5345 = ~(P3_U2365 & P3_U2420); 
assign P3_U5350 = ~(P3_U2365 & P3_U2419); 
assign P3_U5355 = ~(P3_U2365 & P3_U2418); 
assign P3_U5360 = ~(P3_U2365 & P3_U2417); 
assign P3_U5365 = ~(P3_U2365 & P3_U2416); 
assign P3_U5370 = ~(P3_U2365 & P3_U2415); 
assign P3_U5375 = ~(P3_U2365 & P3_U2414); 
assign P3_U5380 = ~(P3_U2365 & P3_U2413); 
assign P3_U5396 = ~(P3_U2364 & P3_U2420); 
assign P3_U5401 = ~(P3_U2364 & P3_U2419); 
assign P3_U5406 = ~(P3_U2364 & P3_U2418); 
assign P3_U5411 = ~(P3_U2364 & P3_U2417); 
assign P3_U5416 = ~(P3_U2364 & P3_U2416); 
assign P3_U5421 = ~(P3_U2364 & P3_U2415); 
assign P3_U5426 = ~(P3_U2364 & P3_U2414); 
assign P3_U5431 = ~(P3_U2364 & P3_U2413); 
assign P3_U5446 = ~(P3_U2363 & P3_U2420); 
assign P3_U5451 = ~(P3_U2363 & P3_U2419); 
assign P3_U5456 = ~(P3_U2363 & P3_U2418); 
assign P3_U5461 = ~(P3_U2363 & P3_U2417); 
assign P3_U5466 = ~(P3_U2363 & P3_U2416); 
assign P3_U5471 = ~(P3_U2363 & P3_U2415); 
assign P3_U5476 = ~(P3_U2363 & P3_U2414); 
assign P3_U5481 = ~(P3_U2363 & P3_U2413); 
assign P3_U5511 = ~(P3_U4323 & P3_U4344); 
assign P3_U5520 = ~(P3_U4324 & P3_U3103); 
assign P3_U5521 = ~(P3_U5518 & P3_U3102); 
assign P3_U5524 = ~(P3_U2452 & P3_U3108); 
assign P3_U5583 = ~(P3_U4647 & P3_U3271); 
assign P3_U5603 = ~(P3_U5602 & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P3_U5604 = ~(P3_U2493 & P3_U4322); 
assign P3_U7375 = ~(P3_U4296 & P3_U2631); 
assign P3_U7918 = ~(P3_U3208 & P3_U3219); 
assign P3_U7919 = ~(P3_U7376 & P3_U3105); 
assign P3_U7976 = ~(P3_U5515 & P3_U3101); 
assign P3_U7977 = ~(P3_U4556 & P3_U5517 & P3_U3110); 
assign P3_U7997 = ~(P3_U7968 & P3_U4647); 
assign P2_U2512 = P2_U8069 & P2_U8068 & P2_U3869; 
assign P2_U2589 = P2_U7581 & P2_U3550 & P2_U4457 & P2_U3549; 
assign P2_U2654 = ~(P2_U7423 & P2_U7422); 
assign P2_U2655 = ~(P2_U4338 & P2_U7424); 
assign P2_U2656 = ~(P2_U4340 & P2_U7427); 
assign P2_U2657 = ~(P2_U4342 & P2_U7429); 
assign P2_U2698 = P2_U3554 & P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P2_U3285 = ~(P2_U4424 & P2_U3709); 
assign P2_U3523 = ~(P2_U4475 & P2_U4427); 
assign P2_U3524 = ~(P2_U4429 & P2_U4475); 
assign P2_U3577 = ~(P2_U4424 & P2_U6845); 
assign P2_U3655 = ~(P2_U8366 & P2_U8365); 
assign P2_U3866 = P2_R2147_U7 & P2_U4466; 
assign P2_U3880 = P2_U5599 & P2_U3254; 
assign P2_U3895 = P2_U5674 & P2_U3578; 
assign P2_U4344 = P2_U7436 & P2_U7435; 
assign P2_U4345 = P2_U7440 & P2_U7439; 
assign P2_U4368 = P2_U7510 & P2_U7509; 
assign P2_U4369 = P2_U7514 & P2_U7513; 
assign P2_U4370 = P2_U7518 & P2_U7517; 
assign P2_U4371 = P2_U7522 & P2_U7521; 
assign P2_U4372 = P2_U7526 & P2_U7525; 
assign P2_U4373 = P2_U7530 & P2_U7529; 
assign P2_U4386 = P2_U7590 & P2_U7589; 
assign P2_U4426 = ~P2_U3549; 
assign P2_U4431 = ~P2_U3578; 
assign P2_U4432 = ~P2_U3254; 
assign P2_U4435 = ~P2_U3296; 
assign P2_U4436 = ~P2_U3522; 
assign P2_U4458 = ~(P2_U4378 & P2_U7577); 
assign P2_U4472 = ~(P2_U2376 & P2_U7871 & P2_U4416); 
assign P2_U4602 = ~(P2_U4424 & P2_U3253); 
assign P2_U5577 = ~(P2_U4428 & P2_U4424); 
assign P2_U5595 = ~(P2_U3877 & P2_U5594); 
assign P2_U5601 = ~(P2_U2436 & P2_U7884); 
assign P2_U5605 = ~(P2_U3296 & P2_U3522); 
assign P2_U5606 = ~(P2_U3578 & P2_U4437); 
assign P2_U5676 = ~(P2_U4417 & P2_U4424); 
assign P2_U5678 = ~(P2_U4428 & P2_U4424); 
assign P2_U6849 = ~(P2_U4418 & P2_U6847); 
assign P2_U7136 = ~P2_U3554; 
assign P2_U7142 = ~(P2_U2354 & P2_U2606); 
assign P2_U7143 = ~(P2_U2605 & P2_U2355); 
assign P2_U7144 = ~(P2_U2354 & P2_U2605); 
assign P2_U7145 = ~(P2_U2604 & P2_U2355); 
assign P2_U7146 = ~(P2_U2354 & P2_U2604); 
assign P2_U7147 = ~(P2_U2603 & P2_U2355); 
assign P2_U7148 = ~(P2_U2354 & P2_U2603); 
assign P2_U7152 = ~(P2_U2602 & P2_U2355); 
assign P2_U7153 = ~(P2_U2354 & P2_U2602); 
assign P2_U7154 = ~(P2_U2601 & P2_U2355); 
assign P2_U7155 = ~(P2_U2354 & P2_U2601); 
assign P2_U7156 = ~(P2_U2600 & P2_U2355); 
assign P2_U7157 = ~(P2_U2354 & P2_U2600); 
assign P2_U7158 = ~(P2_U2599 & P2_U2355); 
assign P2_U7159 = ~(P2_U2354 & P2_U2599); 
assign P2_U7433 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P2_U7437 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P2_U7441 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P2_U7444 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P2_U7447 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P2_U7450 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P2_U7453 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P2_U7456 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P2_U7459 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P2_U7462 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P2_U7465 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P2_U7468 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P2_U7471 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P2_U7474 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P2_U7477 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P2_U7480 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P2_U7483 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P2_U7486 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P2_U7489 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P2_U7492 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P2_U7495 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P2_U7498 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P2_U7501 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P2_U7504 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P2_U7507 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P2_U7511 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P2_U7515 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P2_U7519 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P2_U7523 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P2_U7527 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P2_U7531 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P2_U7534 = ~(P2_U7432 & P2_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P2_U7563 = ~(P2_U7561 & P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P2_U7565 = ~(P2_U7561 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7567 = ~(P2_U7561 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P2_U7569 = ~(P2_U7561 & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P2_U7571 = ~(P2_U7561 & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P2_U7572 = ~(P2_U7561 & P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P2_U7573 = ~(P2_U7561 & P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P2_U7574 = ~(P2_U7561 & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P2_U7575 = ~(P2_U7561 & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P2_U7576 = ~(P2_U7561 & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P2_U7586 = ~(P2_U4381 & P2_U4424); 
assign P2_U7591 = ~(P2_U2376 & P2_U7871 & P2_U4416); 
assign P2_U7728 = ~(P2_R2238_U20 & P2_U2356); 
assign P2_U7737 = ~(P2_U7590 & P2_U7589 & P2_U4422 & P2_U3272); 
assign P2_U7885 = ~(P2_U8348 & P2_U8347 & P2_U3253); 
assign P2_U7887 = ~(P2_U4459 & P2_U5589); 
assign P2_U7889 = ~(P2_U4459 & P2_U5589); 
assign P2_U7897 = ~(P2_U4429 & P2_U5589); 
assign P2_U8076 = ~(P2_U4424 & P2_U3253); 
assign P2_U8077 = ~(P2_U4475 & P2_U7871); 
assign P2_U8096 = ~(P2_U7869 & P2_U5625 & P2_U7867); 
assign P2_U8355 = ~(P2_R2238_U20 & P2_U3283); 
assign P2_U8356 = ~(P2_SUB_450_U18 & P2_U4417); 
assign P2_U8427 = ~(P2_R2238_U20 & P2_U3269); 
assign P1_U2520 = P1_U4219 & P1_U3446; 
assign P1_U2740 = P1_U7063 & P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign P1_U2745 = ~(P1_U7048 & P1_U7047); 
assign P1_U2746 = ~(P1_U7050 & P1_U7049); 
assign P1_U2747 = ~(P1_U7052 & P1_U7051); 
assign P1_U2748 = ~(P1_U7616 & P1_U7053); 
assign P1_U2749 = ~(P1_U7055 & P1_U7054); 
assign P1_U2750 = ~(P1_U7057 & P1_U7056); 
assign P1_U2752 = ~(P1_U4062 & P1_U7060 & P1_U7061); 
assign P1_U2753 = P1_U6957 & P1_U6909; 
assign P1_U2754 = P1_U6974 & P1_U6909; 
assign P1_U2755 = P1_U6991 & P1_U6909; 
assign P1_U2756 = P1_U7615 & P1_U6909; 
assign P1_U2757 = P1_U7023 & P1_U6909; 
assign P1_U2758 = P1_U7040 & P1_U6909; 
assign P1_U2759 = P1_U6909 & P1_U6908; 
assign P1_U2760 = P1_U6926 & P1_U6909; 
assign P1_U3421 = ~(P1_U4194 & P1_U2431); 
assign P1_U3443 = ~(P1_U2450 & P1_U3441); 
assign P1_U3451 = ~(P1_U4254 & P1_U4266); 
assign P1_U3580 = P1_U4217 & P1_U3400; 
assign P1_U3735 = P1_U7496 & P1_U4217; 
assign P1_U3744 = P1_U5500 & P1_U7627 & P1_U3742 & P1_U3743; 
assign P1_U3760 = P1_U3288 & P1_U4217 & P1_U3448; 
assign P1_U3761 = P1_U5566 & P1_U7507; 
assign P1_U4005 = P1_U6758 & P1_U6757; 
assign P1_U4211 = ~P1_U3446; 
assign P1_U4216 = ~P1_U3292; 
assign P1_U4239 = ~(P1_U4477 & P1_U7381); 
assign P1_U5469 = ~(P1_U3733 & P1_U7609); 
assign P1_U5493 = ~(P1_U7629 & P1_U5492); 
assign P1_U5501 = ~(P1_U3292 & P1_U4217); 
assign P1_U5504 = ~(P1_U4218 & P1_U3438); 
assign P1_U5505 = ~(P1_U4214 & P1_U3442); 
assign P1_U5513 = ~(P1_U4214 & P1_U3456); 
assign P1_U5521 = ~(P1_U3292 & P1_U5520); 
assign P1_U5524 = ~(P1_U4214 & P1_U3265); 
assign P1_U5567 = ~(P1_U4266 & P1_U4250); 
assign P1_U6150 = ~(P1_U4254 & P1_U4197 & P1_U4194); 
assign P1_U6607 = ~(P1_U6606 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U6608 = ~(P1_U4193 & P1_U3272); 
assign P1_U6890 = ~(P1_ADD_371_U4 & P1_U4208); 
assign P1_U6928 = ~(P1_U2355 & P1_SUB_357_U8); 
assign P1_U6930 = ~(P1_SUB_357_U6 & P1_U2355); 
assign P1_U6932 = ~(P1_SUB_357_U9 & P1_U2355); 
assign P1_U6934 = ~(P1_SUB_357_U13 & P1_U2355); 
assign P1_U6936 = ~(P1_SUB_357_U11 & P1_U2355); 
assign P1_U6939 = ~(P1_SUB_357_U12 & P1_U2355); 
assign P1_U7042 = ~(P1_SUB_357_U7 & P1_U2355); 
assign P1_U7045 = ~(P1_SUB_357_U10 & P1_U2355); 
assign P1_U7087 = ~P1_U3245; 
assign P1_U7090 = ~(P1_U4067 & P1_U3245); 
assign P1_U7357 = ~(P1_U4234 & P1_U7356); 
assign P1_U7368 = ~(P1_R2238_U20 & P1_U7363); 
assign P1_U7369 = ~(P1_SUB_450_U20 & P1_U2354); 
assign P1_U7370 = ~(P1_R2238_U21 & P1_U7363); 
assign P1_U7372 = ~(P1_R2238_U22 & P1_U7363); 
assign P1_U7374 = ~(P1_R2238_U7 & P1_U7363); 
assign P1_U7378 = ~(P1_R2238_U20 & P1_U4192); 
assign P1_U7473 = ~(P1_U4212 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U7474 = ~(P1_U4213 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U7477 = ~(P1_U7632 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U7480 = ~(P1_U7632 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U7486 = ~(P1_U5491 & P1_U4171 & P1_U4194); 
assign P1_U7488 = ~(P1_U4194 & P1_U3392); 
assign P1_U7504 = ~(P1_U7493 & P1_U7085); 
assign P1_U7505 = ~(P1_U7493 & P1_U7471); 
assign P1_U7606 = ~(P1_U7605 & P1_U3428); 
assign P1_U7608 = ~(P1_U7607 & P1_U3447); 
assign P1_U7611 = ~(P1_U3755 & P1_U7610); 
assign P1_U7699 = ~(P1_U4432 & P1_U5466); 
assign P1_U7717 = ~(P1_U4218 & P1_U3401); 
assign P1_U7725 = ~(P1_U4214 & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P3_ADD_526_U80 = ~(P3_ADD_526_U200 & P3_ADD_526_U199); 
assign P3_ADD_526_U81 = ~(P3_ADD_526_U202 & P3_ADD_526_U201); 
assign P3_ADD_526_U119 = ~P3_ADD_526_U25; 
assign P3_ADD_526_U139 = ~P3_ADD_526_U109; 
assign P3_ADD_526_U196 = ~(P3_ADD_526_U25 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_526_U197 = ~(P3_ADD_526_U109 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_552_U80 = ~(P3_ADD_552_U200 & P3_ADD_552_U199); 
assign P3_ADD_552_U81 = ~(P3_ADD_552_U202 & P3_ADD_552_U201); 
assign P3_ADD_552_U119 = ~P3_ADD_552_U25; 
assign P3_ADD_552_U139 = ~P3_ADD_552_U109; 
assign P3_ADD_552_U196 = ~(P3_ADD_552_U25 & P3_EBX_REG_13__SCAN_IN); 
assign P3_ADD_552_U197 = ~(P3_ADD_552_U109 & P3_EBX_REG_12__SCAN_IN); 
assign P3_ADD_546_U80 = ~(P3_ADD_546_U200 & P3_ADD_546_U199); 
assign P3_ADD_546_U81 = ~(P3_ADD_546_U202 & P3_ADD_546_U201); 
assign P3_ADD_546_U119 = ~P3_ADD_546_U25; 
assign P3_ADD_546_U139 = ~P3_ADD_546_U109; 
assign P3_ADD_546_U196 = ~(P3_ADD_546_U25 & P3_EAX_REG_13__SCAN_IN); 
assign P3_ADD_546_U197 = ~(P3_ADD_546_U109 & P3_EAX_REG_12__SCAN_IN); 
assign P3_ADD_391_1180_U5 = ~P3_U3069; 
assign P3_ADD_391_1180_U6 = ~(P3_U3069 & P3_U2613); 
assign P3_ADD_391_1180_U49 = ~(P3_U3069 & P3_ADD_391_1180_U4); 
assign P3_ADD_476_U64 = ~(P3_ADD_476_U128 & P3_ADD_476_U127); 
assign P3_ADD_476_U99 = ~P3_ADD_476_U16; 
assign P3_ADD_476_U125 = ~(P3_ADD_476_U16 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_531_U68 = ~(P3_ADD_531_U135 & P3_ADD_531_U134); 
assign P3_ADD_531_U103 = ~P3_ADD_531_U17; 
assign P3_ADD_531_U132 = ~(P3_ADD_531_U17 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_SUB_320_U23 = ~(P3_SUB_320_U26 & P3_SUB_320_U56 & P3_SUB_320_U84); 
assign P3_ADD_318_U64 = ~(P3_ADD_318_U128 & P3_ADD_318_U127); 
assign P3_ADD_318_U99 = ~P3_ADD_318_U16; 
assign P3_ADD_318_U125 = ~(P3_ADD_318_U16 & P3_PHYADDRPOINTER_REG_8__SCAN_IN); 
assign P3_SUB_370_U44 = ~(P3_SUB_370_U42 & P3_SUB_370_U43); 
assign P3_SUB_370_U50 = ~(P3_SUB_370_U49 & P3_SUB_370_U42); 
assign P3_ADD_315_U61 = ~(P3_ADD_315_U122 & P3_ADD_315_U121); 
assign P3_ADD_315_U96 = ~P3_ADD_315_U17; 
assign P3_ADD_315_U119 = ~(P3_ADD_315_U17 & P3_PHYADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_360_1242_U24 = ~P3_U2621; 
assign P3_ADD_360_1242_U27 = ~(P3_U2621 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_ADD_360_1242_U258 = ~(P3_U2621 & P3_ADD_360_1242_U25); 
assign P3_ADD_467_U64 = ~(P3_ADD_467_U128 & P3_ADD_467_U127); 
assign P3_ADD_467_U99 = ~P3_ADD_467_U16; 
assign P3_ADD_467_U125 = ~(P3_ADD_467_U16 & P3_REIP_REG_8__SCAN_IN); 
assign P3_ADD_430_U64 = ~(P3_ADD_430_U128 & P3_ADD_430_U127); 
assign P3_ADD_430_U99 = ~P3_ADD_430_U16; 
assign P3_ADD_430_U125 = ~(P3_ADD_430_U16 & P3_REIP_REG_8__SCAN_IN); 
assign P3_ADD_380_U68 = ~(P3_ADD_380_U135 & P3_ADD_380_U134); 
assign P3_ADD_380_U103 = ~P3_ADD_380_U17; 
assign P3_ADD_380_U132 = ~(P3_ADD_380_U17 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_344_U68 = ~(P3_ADD_344_U135 & P3_ADD_344_U134); 
assign P3_ADD_344_U103 = ~P3_ADD_344_U17; 
assign P3_ADD_344_U132 = ~(P3_ADD_344_U17 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_339_U64 = ~(P3_ADD_339_U128 & P3_ADD_339_U127); 
assign P3_ADD_339_U99 = ~P3_ADD_339_U16; 
assign P3_ADD_339_U125 = ~(P3_ADD_339_U16 & P3_PHYADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_360_U4 = ~P3_U2622; 
assign P3_ADD_360_U6 = ~P3_U2623; 
assign P3_ADD_360_U7 = ~(P3_U2623 & P3_U2622); 
assign P3_ADD_360_U8 = ~P3_U2624; 
assign P3_ADD_360_U10 = ~P3_U2625; 
assign P3_ADD_360_U12 = ~P3_U2626; 
assign P3_ADD_360_U14 = ~P3_U2628; 
assign P3_ADD_360_U15 = ~P3_U2627; 
assign P3_ADD_360_U22 = P3_U2628 & P3_U2627; 
assign P3_LT_589_U6 = P3_LT_589_U8 | P3_U2629; 
assign P3_ADD_541_U64 = ~(P3_ADD_541_U128 & P3_ADD_541_U127); 
assign P3_ADD_541_U99 = ~P3_ADD_541_U16; 
assign P3_ADD_541_U125 = ~(P3_ADD_541_U16 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_SUB_355_U44 = ~(P3_SUB_355_U42 & P3_SUB_355_U43); 
assign P3_SUB_355_U50 = ~(P3_SUB_355_U49 & P3_SUB_355_U42); 
assign P3_SUB_450_U42 = ~(P3_SUB_450_U40 & P3_SUB_450_U41); 
assign P3_SUB_450_U47 = ~(P3_SUB_450_U46 & P3_SUB_450_U40); 
assign P3_SUB_485_U42 = ~(P3_SUB_485_U40 & P3_SUB_485_U41); 
assign P3_SUB_485_U47 = ~(P3_SUB_485_U46 & P3_SUB_485_U40); 
assign P3_ADD_515_U64 = ~(P3_ADD_515_U128 & P3_ADD_515_U127); 
assign P3_ADD_515_U99 = ~P3_ADD_515_U16; 
assign P3_ADD_515_U125 = ~(P3_ADD_515_U16 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_394_U65 = ~(P3_ADD_394_U132 & P3_ADD_394_U131); 
assign P3_ADD_394_U102 = ~P3_ADD_394_U16; 
assign P3_ADD_394_U129 = ~(P3_ADD_394_U16 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_SUB_414_U82 = P3_SUB_414_U159 & P3_SUB_414_U158; 
assign P3_SUB_414_U94 = ~P3_SUB_414_U29; 
assign P3_SUB_414_U124 = ~(P3_SUB_414_U123 & P3_EBX_REG_12__SCAN_IN); 
assign P3_SUB_414_U156 = ~(P3_SUB_414_U29 & P3_EBX_REG_13__SCAN_IN); 
assign P3_ADD_441_U64 = ~(P3_ADD_441_U128 & P3_ADD_441_U127); 
assign P3_ADD_441_U99 = ~P3_ADD_441_U16; 
assign P3_ADD_441_U125 = ~(P3_ADD_441_U16 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_349_U68 = ~(P3_ADD_349_U135 & P3_ADD_349_U134); 
assign P3_ADD_349_U103 = ~P3_ADD_349_U17; 
assign P3_ADD_349_U132 = ~(P3_ADD_349_U17 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_405_U65 = ~(P3_ADD_405_U132 & P3_ADD_405_U131); 
assign P3_ADD_405_U102 = ~P3_ADD_405_U16; 
assign P3_ADD_405_U129 = ~(P3_ADD_405_U16 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_553_U68 = ~(P3_ADD_553_U135 & P3_ADD_553_U134); 
assign P3_ADD_553_U103 = ~P3_ADD_553_U17; 
assign P3_ADD_553_U132 = ~(P3_ADD_553_U17 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_558_U68 = ~(P3_ADD_558_U135 & P3_ADD_558_U134); 
assign P3_ADD_558_U103 = ~P3_ADD_558_U17; 
assign P3_ADD_558_U132 = ~(P3_ADD_558_U17 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_385_U68 = ~(P3_ADD_385_U135 & P3_ADD_385_U134); 
assign P3_ADD_385_U103 = ~P3_ADD_385_U17; 
assign P3_ADD_385_U132 = ~(P3_ADD_385_U17 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_547_U68 = ~(P3_ADD_547_U135 & P3_ADD_547_U134); 
assign P3_ADD_547_U103 = ~P3_ADD_547_U17; 
assign P3_ADD_547_U132 = ~(P3_ADD_547_U17 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_SUB_412_U42 = ~(P3_SUB_412_U40 & P3_SUB_412_U41); 
assign P3_SUB_412_U47 = ~(P3_SUB_412_U46 & P3_SUB_412_U40); 
assign P3_SUB_504_U42 = ~(P3_SUB_504_U40 & P3_SUB_504_U41); 
assign P3_SUB_504_U47 = ~(P3_SUB_504_U46 & P3_SUB_504_U40); 
assign P3_SUB_401_U44 = ~(P3_SUB_401_U42 & P3_SUB_401_U43); 
assign P3_SUB_401_U50 = ~(P3_SUB_401_U49 & P3_SUB_401_U42); 
assign P3_ADD_371_U4 = ~P3_U2621; 
assign P3_ADD_371_U7 = ~P3_U2622; 
assign P3_ADD_371_U8 = ~P3_U2624; 
assign P3_ADD_371_U10 = ~P3_U2625; 
assign P3_ADD_371_U12 = ~P3_U2626; 
assign P3_ADD_371_U14 = ~P3_U2628; 
assign P3_ADD_371_U15 = ~P3_U2627; 
assign P3_ADD_371_U16 = ~P3_U2623; 
assign P3_ADD_371_U22 = P3_U2628 & P3_U2627; 
assign P3_ADD_371_U26 = ~(P3_U2622 & P3_U2621); 
assign P3_ADD_371_U32 = ~(P3_U2622 & P3_U2621 & P3_U2623); 
assign P3_SUB_390_U44 = ~(P3_SUB_390_U42 & P3_SUB_390_U43); 
assign P3_SUB_390_U50 = ~(P3_SUB_390_U49 & P3_SUB_390_U42); 
assign P3_SUB_357_U6 = ~P3_U2627; 
assign P3_SUB_357_U7 = ~P3_U2622; 
assign P3_SUB_357_U8 = ~P3_U2628; 
assign P3_SUB_357_U9 = ~P3_U2626; 
assign P3_SUB_357_U10 = ~P3_U2621; 
assign P3_SUB_357_U11 = ~P3_U2624; 
assign P3_SUB_357_U12 = ~P3_U2623; 
assign P3_SUB_357_U13 = ~P3_U2625; 
assign P3_ADD_494_U64 = ~(P3_ADD_494_U128 & P3_ADD_494_U127); 
assign P3_ADD_494_U99 = ~P3_ADD_494_U16; 
assign P3_ADD_494_U125 = ~(P3_ADD_494_U16 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_536_U64 = ~(P3_ADD_536_U128 & P3_ADD_536_U127); 
assign P3_ADD_536_U99 = ~P3_ADD_536_U16; 
assign P3_ADD_536_U125 = ~(P3_ADD_536_U16 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_402_1132_U5 = ~P3_U3069; 
assign P3_ADD_402_1132_U6 = ~(P3_U3069 & P3_U2613); 
assign P3_ADD_402_1132_U49 = ~(P3_U3069 & P3_ADD_402_1132_U4); 
assign P2_ADD_402_1132_U4 = ~P2_U2606; 
assign P2_ADD_402_1132_U6 = ~(P2_U2591 & P2_U2606); 
assign P2_ADD_402_1132_U46 = ~(P2_U2606 & P2_ADD_402_1132_U5); 
assign P2_R2182_U23 = ~P2_U2671; 
assign P2_R2182_U25 = ~P2_U2666; 
assign P2_R2182_U26 = ~P2_U2667; 
assign P2_R2182_U33 = ~P2_U2670; 
assign P2_R2182_U34 = ~P2_U2672; 
assign P2_R2182_U36 = ~P2_U2673; 
assign P2_R2182_U38 = ~P2_U2668; 
assign P2_R2182_U39 = ~P2_U2669; 
assign P2_R2167_U7 = ~P2_U2706; 
assign P2_R2167_U10 = ~P2_U2705; 
assign P2_R2027_U68 = ~(P2_R2027_U135 & P2_R2027_U134); 
assign P2_R2027_U103 = ~P2_R2027_U17; 
assign P2_R2027_U132 = ~(P2_R2027_U17 & P2_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P2_R2337_U62 = ~(P2_R2337_U126 & P2_R2337_U125); 
assign P2_R2337_U100 = ~P2_R2337_U18; 
assign P2_R2337_U123 = ~(P2_R2337_U18 & P2_PHYADDRPOINTER_REG_9__SCAN_IN); 
assign P2_R2219_U20 = ~P2_U2760; 
assign P2_R2219_U21 = ~P2_U2759; 
assign P2_R2219_U22 = ~P2_U2758; 
assign P2_R2219_U58 = ~(P2_U2760 & P2_R2219_U9); 
assign P2_R2219_U62 = ~(P2_U2759 & P2_R2219_U9); 
assign P2_R2219_U67 = ~(P2_U2758 & P2_R2219_U9); 
assign P2_R2219_U82 = ~(P2_U2758 & P2_R2219_U9); 
assign P2_R2219_U87 = ~(P2_U2759 & P2_R2219_U9); 
assign P2_R2219_U92 = ~(P2_U2760 & P2_R2219_U9); 
assign P2_R2096_U60 = ~P2_U2653; 
assign P2_R2096_U62 = ~P2_U2652; 
assign P2_R2096_U64 = ~P2_U2651; 
assign P2_R2096_U66 = ~P2_U2650; 
assign P2_R2238_U44 = ~(P2_R2238_U42 & P2_R2238_U43); 
assign P2_R2238_U50 = ~(P2_R2238_U49 & P2_R2238_U42); 
assign P2_R1957_U23 = ~(P2_R1957_U84 & P2_R1957_U56 & P2_R1957_U26); 
assign P2_SUB_450_U42 = ~(P2_SUB_450_U40 & P2_SUB_450_U41); 
assign P2_SUB_450_U47 = ~(P2_SUB_450_U46 & P2_SUB_450_U40); 
assign P2_ADD_394_U89 = ~(P2_ADD_394_U182 & P2_ADD_394_U181); 
assign P2_ADD_394_U102 = ~P2_ADD_394_U16; 
assign P2_ADD_394_U161 = ~(P2_ADD_394_U16 & P2_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P1_R2027_U80 = ~(P1_R2027_U200 & P1_R2027_U199); 
assign P1_R2027_U81 = ~(P1_R2027_U202 & P1_R2027_U201); 
assign P1_R2027_U119 = ~P1_R2027_U25; 
assign P1_R2027_U139 = ~P1_R2027_U109; 
assign P1_R2027_U196 = ~(P1_R2027_U25 & P1_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P1_R2027_U197 = ~(P1_R2027_U109 & P1_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P1_R2144_U12 = ~P1_U2355; 
assign P1_R2099_U98 = ~(P1_R2099_U346 & P1_R2099_U345); 
assign P1_R2099_U99 = ~P1_U2702; 
assign P1_R2099_U100 = ~P1_U2710; 
assign P1_R2099_U101 = ~P1_U2709; 
assign P1_R2099_U102 = ~P1_U2708; 
assign P1_R2099_U103 = ~P1_U2707; 
assign P1_R2099_U104 = ~P1_U2706; 
assign P1_R2099_U105 = ~P1_U2705; 
assign P1_R2099_U106 = ~P1_U2704; 
assign P1_R2099_U107 = ~P1_U2703; 
assign P1_R2099_U108 = ~P1_U2701; 
assign P1_R2099_U113 = ~P1_U2682; 
assign P1_R2099_U114 = ~P1_U2683; 
assign P1_R2099_U115 = ~P1_U2684; 
assign P1_R2099_U116 = ~P1_U2685; 
assign P1_R2099_U117 = ~P1_U2686; 
assign P1_R2099_U118 = ~P1_U2687; 
assign P1_R2099_U119 = ~P1_U2688; 
assign P1_R2099_U120 = ~P1_U2689; 
assign P1_R2099_U121 = ~P1_U2690; 
assign P1_R2099_U122 = ~P1_U2691; 
assign P1_R2099_U123 = ~P1_U2692; 
assign P1_R2099_U124 = ~P1_U2700; 
assign P1_R2099_U125 = ~P1_U2699; 
assign P1_R2099_U126 = ~P1_U2698; 
assign P1_R2099_U127 = ~P1_U2697; 
assign P1_R2099_U128 = ~P1_U2696; 
assign P1_R2099_U129 = ~P1_U2695; 
assign P1_R2099_U130 = ~P1_U2694; 
assign P1_R2099_U131 = ~P1_U2693; 
assign P1_R2099_U132 = ~P1_U2680; 
assign P1_R2099_U133 = ~P1_U2681; 
assign P1_R2099_U134 = ~P1_U2679; 
assign P1_R2099_U183 = ~(P1_U2702 & P1_R2099_U4); 
assign P1_R2099_U186 = ~(P1_U2710 & P1_R2099_U4); 
assign P1_R2099_U189 = ~(P1_U2709 & P1_R2099_U4); 
assign P1_R2099_U192 = ~(P1_U2708 & P1_R2099_U4); 
assign P1_R2099_U195 = ~(P1_U2707 & P1_R2099_U4); 
assign P1_R2099_U198 = ~(P1_U2706 & P1_R2099_U4); 
assign P1_R2099_U201 = ~(P1_U2705 & P1_R2099_U4); 
assign P1_R2099_U204 = ~(P1_U2704 & P1_R2099_U4); 
assign P1_R2099_U207 = ~(P1_U2703 & P1_R2099_U4); 
assign P1_R2099_U210 = ~(P1_U2701 & P1_R2099_U4); 
assign P1_R2099_U227 = ~(P1_U2682 & P1_R2099_U4); 
assign P1_R2099_U230 = ~(P1_U2683 & P1_R2099_U4); 
assign P1_R2099_U233 = ~(P1_U2684 & P1_R2099_U4); 
assign P1_R2099_U236 = ~(P1_U2685 & P1_R2099_U4); 
assign P1_R2099_U239 = ~(P1_U2686 & P1_R2099_U4); 
assign P1_R2099_U242 = ~(P1_U2687 & P1_R2099_U4); 
assign P1_R2099_U245 = ~(P1_U2688 & P1_R2099_U4); 
assign P1_R2099_U248 = ~(P1_U2689 & P1_R2099_U4); 
assign P1_R2099_U251 = ~(P1_U2690 & P1_R2099_U4); 
assign P1_R2099_U254 = ~(P1_U2691 & P1_R2099_U4); 
assign P1_R2099_U257 = ~(P1_U2692 & P1_R2099_U4); 
assign P1_R2099_U260 = ~(P1_U2700 & P1_R2099_U4); 
assign P1_R2099_U263 = ~(P1_U2699 & P1_R2099_U4); 
assign P1_R2099_U266 = ~(P1_U2698 & P1_R2099_U4); 
assign P1_R2099_U269 = ~(P1_U2697 & P1_R2099_U4); 
assign P1_R2099_U272 = ~(P1_U2696 & P1_R2099_U4); 
assign P1_R2099_U275 = ~(P1_U2695 & P1_R2099_U4); 
assign P1_R2099_U278 = ~(P1_U2694 & P1_R2099_U4); 
assign P1_R2099_U281 = ~(P1_U2693 & P1_R2099_U4); 
assign P1_R2099_U284 = ~(P1_U2680 & P1_R2099_U4); 
assign P1_R2099_U287 = ~(P1_U2681 & P1_R2099_U4); 
assign P1_R2099_U290 = ~(P1_U2679 & P1_R2099_U4); 
assign P1_R2167_U7 = ~P1_U2714; 
assign P1_R2337_U64 = ~(P1_R2337_U128 & P1_R2337_U127); 
assign P1_R2337_U99 = ~P1_R2337_U16; 
assign P1_R2337_U125 = ~(P1_R2337_U16 & P1_PHYADDRPOINTER_REG_8__SCAN_IN); 
assign P1_R2096_U64 = ~(P1_R2096_U128 & P1_R2096_U127); 
assign P1_R2096_U99 = ~P1_R2096_U16; 
assign P1_R2096_U125 = ~(P1_R2096_U16 & P1_REIP_REG_8__SCAN_IN); 
assign P1_R2238_U44 = ~(P1_R2238_U42 & P1_R2238_U43); 
assign P1_R2238_U50 = ~(P1_R2238_U49 & P1_R2238_U42); 
assign P1_SUB_450_U44 = ~(P1_SUB_450_U42 & P1_SUB_450_U43); 
assign P1_SUB_450_U50 = ~(P1_SUB_450_U49 & P1_SUB_450_U42); 
assign P1_ADD_371_U23 = ~(P1_ADD_371_U15 & P1_ADD_371_U26); 
assign P1_ADD_371_U41 = ~(P1_U3228 & P1_ADD_371_U4); 
assign P1_ADD_371_U42 = ~(P1_U3227 & P1_ADD_371_U7); 
assign P1_ADD_405_U89 = ~(P1_ADD_405_U182 & P1_ADD_405_U181); 
assign P1_ADD_405_U102 = ~P1_ADD_405_U16; 
assign P1_ADD_405_U161 = ~(P1_ADD_405_U16 & P1_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P1_ADD_515_U89 = ~(P1_ADD_515_U178 & P1_ADD_515_U177); 
assign P1_ADD_515_U99 = ~P1_ADD_515_U16; 
assign P1_ADD_515_U159 = ~(P1_ADD_515_U16 & P1_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_U2354 = P3_U3688 & P3_U4325; 
assign P3_U2355 = P3_U3689 & P3_U4325; 
assign P3_U2356 = P3_U3355 & P3_U2353; 
assign P3_U2357 = P3_U4323 & P3_U2451; 
assign P3_U2359 = P3_U4324 & P3_U2462; 
assign P3_U2360 = P3_U4296 & P3_U2462; 
assign P3_U2361 = P3_U4297 & P3_U2462; 
assign P3_U2499 = P3_U4658 & P3_U4657; 
assign P3_U2500 = P3_U4658 & P3_U4644; 
assign P3_U2502 = P3_U4658 & P3_U4645; 
assign P3_U2503 = P3_U4658 & P3_U2496; 
assign P3_U2505 = P3_U4644 & P3_U2485; 
assign P3_U2506 = P3_U4645 & P3_U2485; 
assign P3_U2507 = P3_U2496 & P3_U2485; 
assign P3_U2510 = P3_U2509 & P3_U4657; 
assign P3_U2511 = P3_U2509 & P3_U4644; 
assign P3_U2512 = P3_U2509 & P3_U4645; 
assign P3_U2513 = P3_U2509 & P3_U2496; 
assign P3_U3109 = ~(P3_U2353 & P3_U4488); 
assign P3_U3115 = ~(P3_U2451 & P3_U4297); 
assign P3_U3119 = ~(P3_U3356 & P3_U2353); 
assign P3_U3181 = ~(P3_U2485 & P3_U4657); 
assign P3_U3217 = ~(P3_U2450 & P3_U4323); 
assign P3_U3232 = ~P3_LT_589_U6; 
assign P3_U3242 = ~(P3_U3661 & P3_U2450); 
assign P3_U3246 = ~(P3_U3663 & P3_U2449 & P3_U3664); 
assign P3_U3665 = P3_U5511 & P3_U5510 & P3_U5508; 
assign P3_U3666 = P3_U5519 & P3_U4339 & P3_U5520; 
assign P3_U4150 = P3_U7375 & P3_U2630; 
assign P3_U4303 = ~P3_U3117; 
assign P3_U4304 = ~P3_U3116; 
assign P3_U4341 = ~P3_U3229; 
assign P3_U4676 = ~(P3_U2436 & P3_U2488); 
assign P3_U4681 = ~(P3_U2434 & P3_U2488); 
assign P3_U4686 = ~(P3_U2432 & P3_U2488); 
assign P3_U4691 = ~(P3_U2430 & P3_U2488); 
assign P3_U4696 = ~(P3_U2428 & P3_U2488); 
assign P3_U4701 = ~(P3_U2426 & P3_U2488); 
assign P3_U4706 = ~(P3_U2424 & P3_U2488); 
assign P3_U4711 = ~(P3_U2422 & P3_U2488); 
assign P3_U4728 = ~(P3_U2491 & P3_U2436); 
assign P3_U4733 = ~(P3_U2491 & P3_U2434); 
assign P3_U4738 = ~(P3_U2491 & P3_U2432); 
assign P3_U4743 = ~(P3_U2491 & P3_U2430); 
assign P3_U4748 = ~(P3_U2491 & P3_U2428); 
assign P3_U4753 = ~(P3_U2491 & P3_U2426); 
assign P3_U4758 = ~(P3_U2491 & P3_U2424); 
assign P3_U4763 = ~(P3_U2491 & P3_U2422); 
assign P3_U4780 = ~(P3_U2494 & P3_U2436); 
assign P3_U4785 = ~(P3_U2494 & P3_U2434); 
assign P3_U4790 = ~(P3_U2494 & P3_U2432); 
assign P3_U4795 = ~(P3_U2494 & P3_U2430); 
assign P3_U4800 = ~(P3_U2494 & P3_U2428); 
assign P3_U4805 = ~(P3_U2494 & P3_U2426); 
assign P3_U4810 = ~(P3_U2494 & P3_U2424); 
assign P3_U4815 = ~(P3_U2494 & P3_U2422); 
assign P3_U4831 = ~(P3_U2497 & P3_U2436); 
assign P3_U4836 = ~(P3_U2497 & P3_U2434); 
assign P3_U4841 = ~(P3_U2497 & P3_U2432); 
assign P3_U4846 = ~(P3_U2497 & P3_U2430); 
assign P3_U4851 = ~(P3_U2497 & P3_U2428); 
assign P3_U4856 = ~(P3_U2497 & P3_U2426); 
assign P3_U4861 = ~(P3_U2497 & P3_U2424); 
assign P3_U4866 = ~(P3_U2497 & P3_U2422); 
assign P3_U4874 = ~(P3_U4658 & P3_U4657); 
assign P3_U4926 = ~(P3_U4658 & P3_U4644); 
assign P3_U4978 = ~(P3_U4658 & P3_U4645); 
assign P3_U5029 = ~(P3_U4658 & P3_U2496); 
assign P3_U5130 = ~(P3_U4644 & P3_U2485); 
assign P3_U5182 = ~(P3_U4645 & P3_U2485); 
assign P3_U5233 = ~(P3_U2496 & P3_U2485); 
assign P3_U5284 = ~(P3_U2509 & P3_U4657); 
assign P3_U5335 = ~(P3_U2509 & P3_U4644); 
assign P3_U5386 = ~(P3_U2509 & P3_U4645); 
assign P3_U5436 = ~(P3_U2509 & P3_U2496); 
assign P3_U5483 = ~(P3_U7917 & P3_U2514 & P3_U3655 & P3_U4339); 
assign P3_U5484 = ~P3_U3209; 
assign P3_U5485 = ~(P3_U4296 & P3_U3209); 
assign P3_U5526 = ~(P3_U2462 & P3_U3104); 
assign P3_U5527 = ~(P3_U3229 & P3_U3219); 
assign P3_U5532 = ~(P3_U2461 & P3_U5523 & P3_U2450); 
assign P3_U5533 = ~(P3_U3673 & P3_U7918); 
assign P3_U5536 = ~(P3_U3659 & P3_U5523 & P3_U2451); 
assign P3_U5550 = ~(P3_U5548 & P3_U5523 & P3_U2451); 
assign P3_U5578 = ~(P3_U2453 & P3_LT_589_U6 & P3_STATE2_REG_0__SCAN_IN); 
assign P3_U5606 = ~(P3_U5605 & P3_U5603 & P3_U5604); 
assign P3_U7999 = ~(P3_U7998 & P3_U7997); 
assign P2_U2358 = P2_U4431 & P2_STATE2_REG_0__SCAN_IN; 
assign P2_U2618 = ~(P2_U4350 & P2_U7453); 
assign P2_U2619 = ~(P2_U4351 & P2_U7456); 
assign P2_U2620 = ~(P2_U4353 & P2_U7462); 
assign P2_U2621 = ~(P2_U4354 & P2_U7465); 
assign P2_U2622 = ~(P2_U4355 & P2_U7468); 
assign P2_U2623 = ~(P2_U4356 & P2_U7471); 
assign P2_U2624 = ~(P2_U4357 & P2_U7474); 
assign P2_U2625 = ~(P2_U4358 & P2_U7477); 
assign P2_U2626 = ~(P2_U4359 & P2_U7480); 
assign P2_U2627 = ~(P2_U4360 & P2_U7483); 
assign P2_U2628 = ~(P2_U4361 & P2_U7486); 
assign P2_U2629 = ~(P2_U4362 & P2_U7489); 
assign P2_U2630 = ~(P2_U4364 & P2_U7495); 
assign P2_U2631 = ~(P2_U4365 & P2_U7498); 
assign P2_U2632 = ~(P2_U4366 & P2_U7501); 
assign P2_U2633 = ~(P2_U4367 & P2_U7504); 
assign P2_U2634 = ~(P2_U7508 & P2_U7507 & P2_U4368); 
assign P2_U2635 = ~(P2_U7512 & P2_U7511 & P2_U4369); 
assign P2_U2636 = ~(P2_U7516 & P2_U7515 & P2_U4370); 
assign P2_U2637 = ~(P2_U7520 & P2_U7519 & P2_U4371); 
assign P2_U2638 = ~(P2_U7524 & P2_U7523 & P2_U4372); 
assign P2_U2639 = ~(P2_U7528 & P2_U7527 & P2_U4373); 
assign P2_U2640 = ~(P2_U7434 & P2_U7433 & P2_U4344); 
assign P2_U2641 = ~(P2_U7438 & P2_U7437 & P2_U4345); 
assign P2_U2642 = ~(P2_U4346 & P2_U7441); 
assign P2_U2643 = ~(P2_U4347 & P2_U7444); 
assign P2_U2644 = ~(P2_U4348 & P2_U7447); 
assign P2_U2645 = ~(P2_U4349 & P2_U7450); 
assign P2_U2646 = ~(P2_U4352 & P2_U7459); 
assign P2_U2647 = ~(P2_U4363 & P2_U7492); 
assign P2_U2648 = ~(P2_U4374 & P2_U7531); 
assign P2_U2649 = ~(P2_U7534 & P2_U3300 & P2_U4375); 
assign P2_U2690 = ~(P2_U7144 & P2_U7143); 
assign P2_U2691 = ~(P2_U7146 & P2_U7145); 
assign P2_U2692 = ~(P2_U7148 & P2_U7147); 
assign P2_U2693 = ~(P2_U7153 & P2_U7152); 
assign P2_U2694 = ~(P2_U7155 & P2_U7154); 
assign P2_U2695 = ~(P2_U7157 & P2_U7156); 
assign P2_U2696 = ~(P2_U7159 & P2_U7158); 
assign P2_U2704 = ~(P2_U7729 & P2_U7728); 
assign P2_U2753 = ~(P2_U3286 & P2_U7572); 
assign P2_U2754 = ~(P2_U3286 & P2_U7573); 
assign P2_U2755 = ~(P2_U3286 & P2_U7574); 
assign P2_U2756 = ~(P2_U3286 & P2_U7575); 
assign P2_U2757 = ~(P2_U3286 & P2_U7576); 
assign P2_U2761 = ~(P2_U7563 & P2_U7562); 
assign P2_U2762 = ~(P2_U7565 & P2_U7564); 
assign P2_U2763 = ~(P2_U7567 & P2_U7566); 
assign P2_U2764 = ~(P2_U7569 & P2_U7568); 
assign P2_U2765 = ~(P2_U7571 & P2_U7570); 
assign P2_U3650 = ~(P2_U8356 & P2_U8355); 
assign P2_U3686 = ~(P2_U8428 & P2_U8427); 
assign P2_U3881 = P2_U5601 & P2_U5600 & P2_U3880; 
assign P2_U3882 = P2_U7897 & P2_U5602; 
assign P2_U4186 = P2_U4185 & P2_U6849; 
assign P2_U4382 = P2_U3577 & P2_U3539 & P2_U4472 & P2_U7587 & P2_U7586; 
assign P2_U4385 = P2_U7580 & P2_U4458; 
assign P2_U4388 = P2_U3573 & P2_U4458 & P2_U4457 & P2_U3549; 
assign P2_U4423 = ~P2_U3577; 
assign P2_U4425 = ~P2_U3285; 
assign P2_U4433 = ~P2_U3523; 
assign P2_U4434 = ~P2_U3524; 
assign P2_U4603 = ~(P2_U3524 & P2_U4602); 
assign P2_U4604 = ~(P2_U3523 & P2_U3522); 
assign P2_U5578 = ~(P2_U3524 & P2_U5577); 
assign P2_U5604 = ~(P2_U8077 & P2_U8076 & P2_U4470); 
assign P2_U5607 = ~(P2_U4395 & P2_U5605); 
assign P2_U5608 = ~(P2_U3581 & P2_U5606); 
assign P2_U5677 = ~(P2_U5676 & P2_U4470 & P2_U4437 & P2_U3524); 
assign P2_U5679 = ~(P2_U3296 & P2_U5678 & P2_U3523); 
assign P2_U7137 = ~(P2_U7136 & P2_U3300); 
assign P2_U7578 = ~(P2_U4432 & P2_STATE2_REG_0__SCAN_IN); 
assign P2_U7592 = ~(P2_U7591 & P2_U3285 & P2_U4422 & P2_U3539); 
assign P2_U7717 = ~(P2_U4387 & P2_U7885); 
assign P2_U7739 = ~(P2_U7591 & P2_U3285 & P2_U4422 & P2_U3539); 
assign P2_U7896 = ~(P2_U3255 & P2_U5595); 
assign P2_U8091 = ~(P2_U5616 & P2_U5605); 
assign P2_U8092 = ~(P2_U3530 & P2_U5606); 
assign P2_U8097 = ~(P2_U8096 & P2_U8095); 
assign P2_U8363 = ~(P2_R2337_U62 & P2_U3284); 
assign P1_U2518 = P1_U7700 & P1_U7699 & P1_U5468; 
assign P1_U2606 = P1_U7504 & P1_U3427; 
assign P1_U2614 = ~(P1_U6756 & P1_U4005); 
assign P1_U2712 = ~(P1_U7379 & P1_U7378); 
assign P1_U2713 = ~(P1_U4165 & P1_U4239); 
assign P1_U2715 = ~(P1_U4239 & P1_U4167); 
assign P1_U2719 = ~(P1_U4162 & P1_U7370); 
assign P1_U2720 = ~(P1_U4163 & P1_U7372); 
assign P1_U2721 = ~(P1_U4164 & P1_U7374); 
assign P1_U3425 = ~(P1_U4216 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U3746 = P1_U3411 & P1_U3288 & P1_U3745 & P1_U2520 & P1_U3279; 
assign P1_U3748 = P1_U5505 & P1_U5504; 
assign P1_U3757 = P1_U3398 & P1_U3399 & P1_U5567; 
assign P1_U3965 = P1_U6608 & P1_U3298; 
assign P1_U4061 = P1_U7059 & P1_U3443; 
assign P1_U4074 = P1_U7090 & P1_U7089; 
assign P1_U4076 = P1_U7475 & P1_U7476 & P1_U7474; 
assign P1_U4115 = P1_U7486 & P1_U7480 & P1_U7476 & P1_U7474; 
assign P1_U4117 = P1_U7090 & P1_U7089; 
assign P1_U4119 = P1_U7475 & P1_U7476 & P1_U7474; 
assign P1_U4155 = P1_U7357 & P1_U7358 & P1_U4263; 
assign P1_U4161 = P1_U7369 & P1_STATE2_REG_0__SCAN_IN; 
assign P1_U4200 = ~P1_U3421; 
assign P1_U4207 = ~P1_U3443; 
assign P1_U4506 = ~(P1_U3580 & P1_U4505); 
assign P1_U5502 = ~(P1_U3740 & P1_U5501); 
assign P1_U5522 = ~(P1_U5519 & P1_U5521); 
assign P1_U6755 = ~(P1_R2337_U64 & P1_U2352); 
assign P1_U7091 = ~P1_U3451; 
assign P1_U7092 = ~(P1_U3451 & P1_U5492 & P1_U7629); 
assign P1_U7355 = ~(P1_U4153 & P1_U7087); 
assign P1_U7472 = ~(P1_U4211 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U7497 = ~(P1_U3735 & P1_U5469); 
assign P1_U7508 = ~(P1_U3761 & P1_U5565 & P1_U3760); 
assign P1_U7706 = ~(P1_U4477 & P1_U5493); 
assign P1_U7716 = ~(P1_U5511 & P1_U5501); 
assign P1_U7726 = ~(P1_U5521 & P1_U3266); 
assign P3_ADD_526_U27 = ~(P3_ADD_526_U87 & P3_ADD_526_U119); 
assign P3_ADD_526_U108 = ~(P3_ADD_526_U119 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_526_U195 = ~(P3_ADD_526_U119 & P3_ADD_526_U24); 
assign P3_ADD_526_U198 = ~(P3_ADD_526_U139 & P3_ADD_526_U20); 
assign P3_ADD_552_U27 = ~(P3_ADD_552_U87 & P3_ADD_552_U119); 
assign P3_ADD_552_U108 = ~(P3_ADD_552_U119 & P3_EBX_REG_13__SCAN_IN); 
assign P3_ADD_552_U195 = ~(P3_ADD_552_U119 & P3_ADD_552_U24); 
assign P3_ADD_552_U198 = ~(P3_ADD_552_U139 & P3_ADD_552_U20); 
assign P3_ADD_546_U27 = ~(P3_ADD_546_U87 & P3_ADD_546_U119); 
assign P3_ADD_546_U108 = ~(P3_ADD_546_U119 & P3_EAX_REG_13__SCAN_IN); 
assign P3_ADD_546_U195 = ~(P3_ADD_546_U119 & P3_ADD_546_U24); 
assign P3_ADD_546_U198 = ~(P3_ADD_546_U139 & P3_ADD_546_U20); 
assign P3_ADD_391_1180_U28 = ~P3_ADD_391_1180_U6; 
assign P3_ADD_391_1180_U47 = ~(P3_U2614 & P3_ADD_391_1180_U6); 
assign P3_ADD_391_1180_U50 = ~(P3_U2613 & P3_ADD_391_1180_U5); 
assign P3_ADD_476_U19 = ~(P3_ADD_476_U99 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_476_U126 = ~(P3_ADD_476_U99 & P3_ADD_476_U17); 
assign P3_ADD_531_U19 = ~(P3_ADD_531_U103 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_531_U133 = ~(P3_ADD_531_U103 & P3_ADD_531_U18); 
assign P3_SUB_320_U19 = P3_SUB_320_U90 & P3_SUB_320_U23; 
assign P3_SUB_320_U54 = ~P3_ADD_318_U64; 
assign P3_SUB_320_U85 = ~P3_SUB_320_U23; 
assign P3_SUB_320_U130 = ~(P3_ADD_318_U64 & P3_SUB_320_U23); 
assign P3_ADD_318_U19 = ~(P3_ADD_318_U99 & P3_PHYADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_318_U126 = ~(P3_ADD_318_U99 & P3_ADD_318_U17); 
assign P3_SUB_370_U6 = ~(P3_SUB_370_U45 & P3_SUB_370_U44); 
assign P3_SUB_370_U19 = ~(P3_SUB_370_U51 & P3_SUB_370_U50); 
assign P3_ADD_315_U18 = ~(P3_ADD_315_U96 & P3_PHYADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_315_U120 = ~(P3_ADD_315_U96 & P3_ADD_315_U16); 
assign P3_ADD_360_1242_U28 = ~P3_ADD_360_U4; 
assign P3_ADD_360_1242_U124 = ~P3_ADD_360_1242_U27; 
assign P3_ADD_360_1242_U244 = ~(P3_ADD_360_1242_U27 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_360_1242_U247 = ~(P3_ADD_360_1242_U27 & P3_ADD_360_1242_U26 & P3_ADD_360_U4); 
assign P3_ADD_360_1242_U257 = ~(P3_ADD_360_1242_U24 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_ADD_467_U19 = ~(P3_ADD_467_U99 & P3_REIP_REG_8__SCAN_IN); 
assign P3_ADD_467_U126 = ~(P3_ADD_467_U99 & P3_ADD_467_U17); 
assign P3_ADD_430_U19 = ~(P3_ADD_430_U99 & P3_REIP_REG_8__SCAN_IN); 
assign P3_ADD_430_U126 = ~(P3_ADD_430_U99 & P3_ADD_430_U17); 
assign P3_ADD_380_U19 = ~(P3_ADD_380_U103 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_380_U133 = ~(P3_ADD_380_U103 & P3_ADD_380_U18); 
assign P3_ADD_344_U19 = ~(P3_ADD_344_U103 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_344_U133 = ~(P3_ADD_344_U103 & P3_ADD_344_U18); 
assign P3_ADD_339_U19 = ~(P3_ADD_339_U99 & P3_PHYADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_339_U126 = ~(P3_ADD_339_U99 & P3_ADD_339_U17); 
assign P3_ADD_360_U24 = ~P3_ADD_360_U7; 
assign P3_ADD_360_U37 = ~(P3_U2624 & P3_ADD_360_U7); 
assign P3_ADD_360_U39 = ~(P3_U2623 & P3_ADD_360_U4); 
assign P3_ADD_360_U40 = ~(P3_U2622 & P3_ADD_360_U6); 
assign P3_ADD_541_U19 = ~(P3_ADD_541_U99 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_541_U126 = ~(P3_ADD_541_U99 & P3_ADD_541_U17); 
assign P3_SUB_355_U6 = ~(P3_SUB_355_U45 & P3_SUB_355_U44); 
assign P3_SUB_355_U19 = ~(P3_SUB_355_U51 & P3_SUB_355_U50); 
assign P3_SUB_450_U6 = ~(P3_SUB_450_U43 & P3_SUB_450_U42); 
assign P3_SUB_450_U16 = ~(P3_SUB_450_U48 & P3_SUB_450_U47); 
assign P3_SUB_357_1258_U31 = ~P3_SUB_357_U7; 
assign P3_SUB_357_1258_U271 = ~(P3_SUB_357_U7 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_SUB_485_U6 = ~(P3_SUB_485_U43 & P3_SUB_485_U42); 
assign P3_SUB_485_U16 = ~(P3_SUB_485_U48 & P3_SUB_485_U47); 
assign P3_ADD_515_U19 = ~(P3_ADD_515_U99 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_515_U126 = ~(P3_ADD_515_U99 & P3_ADD_515_U17); 
assign P3_ADD_394_U19 = ~(P3_ADD_394_U102 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_394_U130 = ~(P3_ADD_394_U102 & P3_ADD_394_U17); 
assign P3_SUB_414_U7 = P3_SUB_414_U124 & P3_SUB_414_U29; 
assign P3_SUB_414_U30 = ~(P3_SUB_414_U47 & P3_SUB_414_U79 & P3_SUB_414_U94); 
assign P3_SUB_414_U121 = ~(P3_SUB_414_U94 & P3_SUB_414_U79); 
assign P3_SUB_414_U157 = ~(P3_SUB_414_U94 & P3_SUB_414_U79); 
assign P3_ADD_441_U19 = ~(P3_ADD_441_U99 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_441_U126 = ~(P3_ADD_441_U99 & P3_ADD_441_U17); 
assign P3_ADD_349_U19 = ~(P3_ADD_349_U103 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_349_U133 = ~(P3_ADD_349_U103 & P3_ADD_349_U18); 
assign P3_ADD_405_U19 = ~(P3_ADD_405_U102 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_405_U130 = ~(P3_ADD_405_U102 & P3_ADD_405_U17); 
assign P3_ADD_553_U19 = ~(P3_ADD_553_U103 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_553_U133 = ~(P3_ADD_553_U103 & P3_ADD_553_U18); 
assign P3_ADD_558_U19 = ~(P3_ADD_558_U103 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_558_U133 = ~(P3_ADD_558_U103 & P3_ADD_558_U18); 
assign P3_ADD_385_U19 = ~(P3_ADD_385_U103 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_385_U133 = ~(P3_ADD_385_U103 & P3_ADD_385_U18); 
assign P3_ADD_357_U10 = ~P3_SUB_357_U10; 
assign P3_ADD_357_U11 = P3_SUB_357_U7 | P3_SUB_357_U12 | P3_SUB_357_U11; 
assign P3_ADD_357_U14 = ~(P3_SUB_357_U13 | P3_SUB_357_U9); 
assign P3_ADD_357_U15 = ~(P3_SUB_357_U6 | P3_SUB_357_U8); 
assign P3_ADD_357_U16 = ~P3_SUB_357_U6; 
assign P3_ADD_357_U18 = ~P3_SUB_357_U13; 
assign P3_ADD_357_U20 = ~P3_SUB_357_U7; 
assign P3_ADD_357_U21 = ~P3_SUB_357_U12; 
assign P3_ADD_357_U28 = P3_SUB_357_U7 | P3_SUB_357_U12; 
assign P3_ADD_547_U19 = ~(P3_ADD_547_U103 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_547_U133 = ~(P3_ADD_547_U103 & P3_ADD_547_U18); 
assign P3_SUB_412_U6 = ~(P3_SUB_412_U43 & P3_SUB_412_U42); 
assign P3_SUB_412_U16 = ~(P3_SUB_412_U48 & P3_SUB_412_U47); 
assign P3_ADD_371_1212_U31 = ~P3_ADD_371_U4; 
assign P3_ADD_371_1212_U34 = ~(P3_ADD_371_U4 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_ADD_371_1212_U265 = ~(P3_ADD_371_U4 & P3_ADD_371_1212_U32); 
assign P3_SUB_504_U6 = ~(P3_SUB_504_U43 & P3_SUB_504_U42); 
assign P3_SUB_504_U16 = ~(P3_SUB_504_U48 & P3_SUB_504_U47); 
assign P3_SUB_401_U6 = ~(P3_SUB_401_U45 & P3_SUB_401_U44); 
assign P3_SUB_401_U19 = ~(P3_SUB_401_U51 & P3_SUB_401_U50); 
assign P3_ADD_371_U24 = ~(P3_ADD_371_U16 & P3_ADD_371_U26); 
assign P3_ADD_371_U43 = ~(P3_U2622 & P3_ADD_371_U4); 
assign P3_ADD_371_U44 = ~(P3_U2621 & P3_ADD_371_U7); 
assign P3_SUB_390_U6 = ~(P3_SUB_390_U45 & P3_SUB_390_U44); 
assign P3_SUB_390_U19 = ~(P3_SUB_390_U51 & P3_SUB_390_U50); 
assign P3_ADD_494_U19 = ~(P3_ADD_494_U99 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_494_U126 = ~(P3_ADD_494_U99 & P3_ADD_494_U17); 
assign P3_ADD_536_U19 = ~(P3_ADD_536_U99 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_536_U126 = ~(P3_ADD_536_U99 & P3_ADD_536_U17); 
assign P3_ADD_402_1132_U28 = ~P3_ADD_402_1132_U6; 
assign P3_ADD_402_1132_U47 = ~(P3_U2614 & P3_ADD_402_1132_U6); 
assign P3_ADD_402_1132_U50 = ~(P3_U2613 & P3_ADD_402_1132_U5); 
assign P2_ADD_402_1132_U28 = ~P2_ADD_402_1132_U6; 
assign P2_ADD_402_1132_U39 = ~(P2_U2592 & P2_ADD_402_1132_U6); 
assign P2_ADD_402_1132_U45 = ~(P2_U2591 & P2_ADD_402_1132_U4); 
assign P2_R2182_U50 = ~P2_U2698; 
assign P2_R2182_U133 = P2_U2698 | P2_U2677; 
assign P2_R2182_U135 = ~(P2_U2677 & P2_U2698); 
assign P2_R2182_U204 = ~(P2_U2698 & P2_R2182_U51); 
assign P2_R2182_U206 = ~(P2_U2698 & P2_R2182_U51); 
assign P2_R2027_U19 = ~(P2_R2027_U103 & P2_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P2_R2027_U133 = ~(P2_R2027_U103 & P2_R2027_U18); 
assign P2_R2337_U19 = ~(P2_R2337_U100 & P2_PHYADDRPOINTER_REG_9__SCAN_IN); 
assign P2_R2337_U124 = ~(P2_R2337_U100 & P2_R2337_U17); 
assign P2_R2219_U60 = ~(P2_U4428 & P2_R2219_U20); 
assign P2_R2219_U64 = ~(P2_U4428 & P2_R2219_U21); 
assign P2_R2219_U66 = ~(P2_U4428 & P2_R2219_U22); 
assign P2_R2219_U83 = ~(P2_U4428 & P2_R2219_U22); 
assign P2_R2219_U88 = ~(P2_U4428 & P2_R2219_U21); 
assign P2_R2219_U93 = ~(P2_U4428 & P2_R2219_U20); 
assign P2_R2096_U52 = ~P2_U2657; 
assign P2_R2096_U55 = ~P2_U2656; 
assign P2_R2096_U56 = ~P2_U2655; 
assign P2_R2096_U58 = ~P2_U2654; 
assign P2_R2238_U6 = ~(P2_R2238_U45 & P2_R2238_U44); 
assign P2_R2238_U19 = ~(P2_R2238_U51 & P2_R2238_U50); 
assign P2_R1957_U19 = P2_R1957_U90 & P2_R1957_U23; 
assign P2_R1957_U54 = ~P2_U3655; 
assign P2_R1957_U85 = ~P2_R1957_U23; 
assign P2_R1957_U130 = ~(P2_U3655 & P2_R1957_U23); 
assign P2_SUB_450_U6 = ~(P2_SUB_450_U43 & P2_SUB_450_U42); 
assign P2_SUB_450_U17 = ~(P2_SUB_450_U48 & P2_SUB_450_U47); 
assign P2_ADD_394_U18 = ~(P2_ADD_394_U102 & P2_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P2_ADD_394_U162 = ~(P2_ADD_394_U102 & P2_ADD_394_U17); 
assign P1_R2027_U27 = ~(P1_R2027_U87 & P1_R2027_U119); 
assign P1_R2027_U108 = ~(P1_R2027_U119 & P1_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P1_R2027_U195 = ~(P1_R2027_U119 & P1_R2027_U24); 
assign P1_R2027_U198 = ~(P1_R2027_U139 & P1_R2027_U20); 
assign P1_R2182_U12 = ~P1_U2740; 
assign P1_R2144_U13 = ~P1_U2750; 
assign P1_R2144_U15 = ~P1_U2752; 
assign P1_R2144_U16 = ~P1_U2749; 
assign P1_R2144_U17 = ~P1_U2745; 
assign P1_R2144_U18 = ~P1_U2748; 
assign P1_R2144_U20 = ~P1_U2747; 
assign P1_R2144_U22 = ~P1_U2746; 
assign P1_R2144_U76 = ~P1_U2760; 
assign P1_R2144_U77 = ~P1_U2759; 
assign P1_R2144_U85 = ~P1_U2754; 
assign P1_R2144_U86 = ~P1_U2753; 
assign P1_R2144_U87 = ~P1_U2755; 
assign P1_R2144_U88 = ~P1_U2756; 
assign P1_R2144_U89 = ~P1_U2757; 
assign P1_R2144_U90 = ~P1_U2758; 
assign P1_R2144_U203 = ~(P1_U2760 & P1_R2144_U12); 
assign P1_R2144_U206 = ~(P1_U2759 & P1_R2144_U12); 
assign P1_R2144_U221 = ~(P1_U2754 & P1_R2144_U12); 
assign P1_R2144_U224 = ~(P1_U2753 & P1_R2144_U12); 
assign P1_R2144_U227 = ~(P1_U2755 & P1_R2144_U12); 
assign P1_R2144_U230 = ~(P1_U2756 & P1_R2144_U12); 
assign P1_R2144_U233 = ~(P1_U2757 & P1_R2144_U12); 
assign P1_R2144_U236 = ~(P1_U2758 & P1_R2144_U12); 
assign P1_R2099_U182 = ~(P1_U4190 & P1_R2099_U99); 
assign P1_R2099_U185 = ~(P1_U4190 & P1_R2099_U100); 
assign P1_R2099_U188 = ~(P1_U4190 & P1_R2099_U101); 
assign P1_R2099_U191 = ~(P1_U4190 & P1_R2099_U102); 
assign P1_R2099_U194 = ~(P1_U4190 & P1_R2099_U103); 
assign P1_R2099_U197 = ~(P1_U4190 & P1_R2099_U104); 
assign P1_R2099_U200 = ~(P1_U4190 & P1_R2099_U105); 
assign P1_R2099_U203 = ~(P1_U4190 & P1_R2099_U106); 
assign P1_R2099_U206 = ~(P1_U4190 & P1_R2099_U107); 
assign P1_R2099_U209 = ~(P1_U4190 & P1_R2099_U108); 
assign P1_R2099_U226 = ~(P1_U4190 & P1_R2099_U113); 
assign P1_R2099_U229 = ~(P1_U4190 & P1_R2099_U114); 
assign P1_R2099_U232 = ~(P1_U4190 & P1_R2099_U115); 
assign P1_R2099_U235 = ~(P1_U4190 & P1_R2099_U116); 
assign P1_R2099_U238 = ~(P1_U4190 & P1_R2099_U117); 
assign P1_R2099_U241 = ~(P1_U4190 & P1_R2099_U118); 
assign P1_R2099_U244 = ~(P1_U4190 & P1_R2099_U119); 
assign P1_R2099_U247 = ~(P1_U4190 & P1_R2099_U120); 
assign P1_R2099_U250 = ~(P1_U4190 & P1_R2099_U121); 
assign P1_R2099_U253 = ~(P1_U4190 & P1_R2099_U122); 
assign P1_R2099_U256 = ~(P1_U4190 & P1_R2099_U123); 
assign P1_R2099_U259 = ~(P1_U4190 & P1_R2099_U124); 
assign P1_R2099_U262 = ~(P1_U4190 & P1_R2099_U125); 
assign P1_R2099_U265 = ~(P1_U4190 & P1_R2099_U126); 
assign P1_R2099_U268 = ~(P1_U4190 & P1_R2099_U127); 
assign P1_R2099_U271 = ~(P1_U4190 & P1_R2099_U128); 
assign P1_R2099_U274 = ~(P1_U4190 & P1_R2099_U129); 
assign P1_R2099_U277 = ~(P1_U4190 & P1_R2099_U130); 
assign P1_R2099_U280 = ~(P1_U4190 & P1_R2099_U131); 
assign P1_R2099_U283 = ~(P1_U4190 & P1_R2099_U132); 
assign P1_R2099_U286 = ~(P1_U4190 & P1_R2099_U133); 
assign P1_R2099_U289 = ~(P1_U4190 & P1_R2099_U134); 
assign P1_R2099_U347 = ~P1_R2099_U98; 
assign P1_R2337_U19 = ~(P1_R2337_U99 & P1_PHYADDRPOINTER_REG_8__SCAN_IN); 
assign P1_R2337_U126 = ~(P1_R2337_U99 & P1_R2337_U17); 
assign P1_R2096_U19 = ~(P1_R2096_U99 & P1_REIP_REG_8__SCAN_IN); 
assign P1_R2096_U126 = ~(P1_R2096_U99 & P1_R2096_U17); 
assign P1_R2238_U6 = ~(P1_R2238_U45 & P1_R2238_U44); 
assign P1_R2238_U19 = ~(P1_R2238_U51 & P1_R2238_U50); 
assign P1_SUB_450_U6 = ~(P1_SUB_450_U45 & P1_SUB_450_U44); 
assign P1_SUB_450_U19 = ~(P1_SUB_450_U51 & P1_SUB_450_U50); 
assign P1_ADD_371_U5 = ~(P1_ADD_371_U23 & P1_ADD_371_U31); 
assign P1_ADD_371_U9 = ~(P1_U3230 & P1_ADD_371_U23); 
assign P1_ADD_371_U20 = ~(P1_ADD_371_U42 & P1_ADD_371_U41); 
assign P1_ADD_371_U27 = ~P1_ADD_371_U23; 
assign P1_ADD_371_U39 = ~(P1_U3230 & P1_ADD_371_U23); 
assign P1_ADD_405_U18 = ~(P1_ADD_405_U102 & P1_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P1_ADD_405_U162 = ~(P1_ADD_405_U102 & P1_ADD_405_U17); 
assign P1_ADD_515_U18 = ~(P1_ADD_515_U99 & P1_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P1_ADD_515_U160 = ~(P1_ADD_515_U99 & P1_ADD_515_U17); 
assign P3_U2358 = P3_U3690 & P3_U4341; 
assign P3_U2362 = P3_U3691 & P3_U4341; 
assign P3_U2393 = P3_U2628 & P3_U2361; 
assign P3_U2395 = P3_U2361 & P3_U3241; 
assign P3_U2517 = P3_U3246 & P3_U5526; 
assign P3_U3182 = ~(P3_U3368 & P3_U3181); 
assign P3_U3233 = ~(P3_U4330 & P3_U3127 & P3_U5578); 
assign P3_U3283 = P3_U3652 & P3_U2356; 
assign P3_U3303 = P3_ADD_495_U8 & P3_U2356; 
assign P3_U3370 = P3_U4676 & P3_U4675; 
assign P3_U3372 = P3_U4681 & P3_U4680; 
assign P3_U3374 = P3_U4686 & P3_U4685; 
assign P3_U3376 = P3_U4691 & P3_U4690; 
assign P3_U3378 = P3_U4696 & P3_U4695; 
assign P3_U3380 = P3_U4701 & P3_U4700; 
assign P3_U3382 = P3_U4706 & P3_U4705; 
assign P3_U3384 = P3_U4711 & P3_U4710; 
assign P3_U3388 = P3_U4728 & P3_U4727; 
assign P3_U3390 = P3_U4733 & P3_U4732; 
assign P3_U3392 = P3_U4738 & P3_U4737; 
assign P3_U3394 = P3_U4743 & P3_U4742; 
assign P3_U3396 = P3_U4748 & P3_U4747; 
assign P3_U3398 = P3_U4753 & P3_U4752; 
assign P3_U3400 = P3_U4758 & P3_U4757; 
assign P3_U3402 = P3_U4763 & P3_U4762; 
assign P3_U3406 = P3_U4780 & P3_U4779; 
assign P3_U3408 = P3_U4785 & P3_U4784; 
assign P3_U3410 = P3_U4790 & P3_U4789; 
assign P3_U3412 = P3_U4795 & P3_U4794; 
assign P3_U3414 = P3_U4800 & P3_U4799; 
assign P3_U3416 = P3_U4805 & P3_U4804; 
assign P3_U3418 = P3_U4810 & P3_U4809; 
assign P3_U3420 = P3_U4815 & P3_U4814; 
assign P3_U3424 = P3_U4831 & P3_U4830; 
assign P3_U3426 = P3_U4836 & P3_U4835; 
assign P3_U3428 = P3_U4841 & P3_U4840; 
assign P3_U3430 = P3_U4846 & P3_U4845; 
assign P3_U3432 = P3_U4851 & P3_U4850; 
assign P3_U3434 = P3_U4856 & P3_U4855; 
assign P3_U3436 = P3_U4861 & P3_U4860; 
assign P3_U3438 = P3_U4866 & P3_U4865; 
assign P3_U3667 = P3_U7978 & P3_U7977 & P3_U5521 & P3_U3666; 
assign P3_U3671 = P3_U3116 & P3_U3117 & P3_U3119; 
assign P3_U3674 = P3_U5533 & P3_U5532; 
assign P3_U4298 = ~P3_U3242; 
assign P3_U4302 = ~P3_U3119; 
assign P3_U4305 = ~P3_U3115; 
assign P3_U4306 = ~P3_U3246; 
assign P3_U4314 = ~P3_U3217; 
assign P3_U4326 = ~P3_U3181; 
assign P3_U4337 = ~(P3_U2453 & P3_U3232); 
assign P3_U4619 = ~P3_U3109; 
assign P3_U4626 = ~(P3_U3353 & P3_U4303); 
assign P3_U4883 = ~(P3_U2499 & P3_U2436); 
assign P3_U4888 = ~(P3_U2499 & P3_U2434); 
assign P3_U4893 = ~(P3_U2499 & P3_U2432); 
assign P3_U4898 = ~(P3_U2499 & P3_U2430); 
assign P3_U4903 = ~(P3_U2499 & P3_U2428); 
assign P3_U4908 = ~(P3_U2499 & P3_U2426); 
assign P3_U4913 = ~(P3_U2499 & P3_U2424); 
assign P3_U4918 = ~(P3_U2499 & P3_U2422); 
assign P3_U4935 = ~(P3_U2500 & P3_U2436); 
assign P3_U4940 = ~(P3_U2500 & P3_U2434); 
assign P3_U4945 = ~(P3_U2500 & P3_U2432); 
assign P3_U4950 = ~(P3_U2500 & P3_U2430); 
assign P3_U4955 = ~(P3_U2500 & P3_U2428); 
assign P3_U4960 = ~(P3_U2500 & P3_U2426); 
assign P3_U4965 = ~(P3_U2500 & P3_U2424); 
assign P3_U4970 = ~(P3_U2500 & P3_U2422); 
assign P3_U4987 = ~(P3_U2502 & P3_U2436); 
assign P3_U4992 = ~(P3_U2502 & P3_U2434); 
assign P3_U4997 = ~(P3_U2502 & P3_U2432); 
assign P3_U5002 = ~(P3_U2502 & P3_U2430); 
assign P3_U5007 = ~(P3_U2502 & P3_U2428); 
assign P3_U5012 = ~(P3_U2502 & P3_U2426); 
assign P3_U5017 = ~(P3_U2502 & P3_U2424); 
assign P3_U5022 = ~(P3_U2502 & P3_U2422); 
assign P3_U5038 = ~(P3_U2503 & P3_U2436); 
assign P3_U5043 = ~(P3_U2503 & P3_U2434); 
assign P3_U5048 = ~(P3_U2503 & P3_U2432); 
assign P3_U5053 = ~(P3_U2503 & P3_U2430); 
assign P3_U5058 = ~(P3_U2503 & P3_U2428); 
assign P3_U5063 = ~(P3_U2503 & P3_U2426); 
assign P3_U5068 = ~(P3_U2503 & P3_U2424); 
assign P3_U5073 = ~(P3_U2503 & P3_U2422); 
assign P3_U5139 = ~(P3_U2505 & P3_U2436); 
assign P3_U5144 = ~(P3_U2505 & P3_U2434); 
assign P3_U5149 = ~(P3_U2505 & P3_U2432); 
assign P3_U5154 = ~(P3_U2505 & P3_U2430); 
assign P3_U5159 = ~(P3_U2505 & P3_U2428); 
assign P3_U5164 = ~(P3_U2505 & P3_U2426); 
assign P3_U5169 = ~(P3_U2505 & P3_U2424); 
assign P3_U5174 = ~(P3_U2505 & P3_U2422); 
assign P3_U5191 = ~(P3_U2506 & P3_U2436); 
assign P3_U5196 = ~(P3_U2506 & P3_U2434); 
assign P3_U5201 = ~(P3_U2506 & P3_U2432); 
assign P3_U5206 = ~(P3_U2506 & P3_U2430); 
assign P3_U5211 = ~(P3_U2506 & P3_U2428); 
assign P3_U5216 = ~(P3_U2506 & P3_U2426); 
assign P3_U5221 = ~(P3_U2506 & P3_U2424); 
assign P3_U5226 = ~(P3_U2506 & P3_U2422); 
assign P3_U5241 = ~(P3_U2507 & P3_U2436); 
assign P3_U5246 = ~(P3_U2507 & P3_U2434); 
assign P3_U5251 = ~(P3_U2507 & P3_U2432); 
assign P3_U5256 = ~(P3_U2507 & P3_U2430); 
assign P3_U5261 = ~(P3_U2507 & P3_U2428); 
assign P3_U5266 = ~(P3_U2507 & P3_U2426); 
assign P3_U5271 = ~(P3_U2507 & P3_U2424); 
assign P3_U5276 = ~(P3_U2507 & P3_U2422); 
assign P3_U5292 = ~(P3_U2510 & P3_U2436); 
assign P3_U5297 = ~(P3_U2510 & P3_U2434); 
assign P3_U5302 = ~(P3_U2510 & P3_U2432); 
assign P3_U5307 = ~(P3_U2510 & P3_U2430); 
assign P3_U5312 = ~(P3_U2510 & P3_U2428); 
assign P3_U5317 = ~(P3_U2510 & P3_U2426); 
assign P3_U5322 = ~(P3_U2510 & P3_U2424); 
assign P3_U5327 = ~(P3_U2510 & P3_U2422); 
assign P3_U5343 = ~(P3_U2511 & P3_U2436); 
assign P3_U5348 = ~(P3_U2511 & P3_U2434); 
assign P3_U5353 = ~(P3_U2511 & P3_U2432); 
assign P3_U5358 = ~(P3_U2511 & P3_U2430); 
assign P3_U5363 = ~(P3_U2511 & P3_U2428); 
assign P3_U5368 = ~(P3_U2511 & P3_U2426); 
assign P3_U5373 = ~(P3_U2511 & P3_U2424); 
assign P3_U5378 = ~(P3_U2511 & P3_U2422); 
assign P3_U5394 = ~(P3_U2512 & P3_U2436); 
assign P3_U5399 = ~(P3_U2512 & P3_U2434); 
assign P3_U5404 = ~(P3_U2512 & P3_U2432); 
assign P3_U5409 = ~(P3_U2512 & P3_U2430); 
assign P3_U5414 = ~(P3_U2512 & P3_U2428); 
assign P3_U5419 = ~(P3_U2512 & P3_U2426); 
assign P3_U5424 = ~(P3_U2512 & P3_U2424); 
assign P3_U5429 = ~(P3_U2512 & P3_U2422); 
assign P3_U5444 = ~(P3_U2513 & P3_U2436); 
assign P3_U5449 = ~(P3_U2513 & P3_U2434); 
assign P3_U5454 = ~(P3_U2513 & P3_U2432); 
assign P3_U5459 = ~(P3_U2513 & P3_U2430); 
assign P3_U5464 = ~(P3_U2513 & P3_U2428); 
assign P3_U5469 = ~(P3_U2513 & P3_U2426); 
assign P3_U5474 = ~(P3_U2513 & P3_U2424); 
assign P3_U5479 = ~(P3_U2513 & P3_U2422); 
assign P3_U5507 = ~(P3_U5484 & P3_U3107); 
assign P3_U5528 = ~(P3_U2456 & P3_U5527); 
assign P3_U5541 = ~(P3_ADD_495_U9 & P3_U2356); 
assign P3_U5552 = ~(P3_ADD_495_U10 & P3_U2356); 
assign P3_U5559 = ~(P3_U4341 & P3_U4608); 
assign P3_U5565 = ~(P3_ADD_495_U4 & P3_U2356); 
assign P3_U5572 = ~(P3_U2356 & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P3_U5593 = ~(P3_U4322 & P3_U7999); 
assign P3_U5639 = ~(P3_U2354 & P3_ADD_531_U5); 
assign P3_U5640 = ~(P3_U2355 & P3_ADD_526_U5); 
assign P3_U5642 = ~(P3_U2356 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_U5643 = ~(P3_U4303 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_U5644 = ~(P3_U4304 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_U5646 = ~(P3_ADD_394_U4 & P3_U2357); 
assign P3_U5648 = ~(P3_U2359 & P3_ADD_380_U5); 
assign P3_U5663 = ~(P3_ADD_531_U85 & P3_U2354); 
assign P3_U5664 = ~(P3_ADD_526_U71 & P3_U2355); 
assign P3_U5666 = ~(P3_ADD_494_U4 & P3_U2356); 
assign P3_U5667 = ~(P3_ADD_476_U4 & P3_U4303); 
assign P3_U5668 = ~(P3_ADD_441_U4 & P3_U4304); 
assign P3_U5670 = ~(P3_ADD_394_U81 & P3_U2357); 
assign P3_U5672 = ~(P3_ADD_380_U85 & P3_U2359); 
assign P3_U5687 = ~(P3_ADD_531_U74 & P3_U2354); 
assign P3_U5688 = ~(P3_ADD_526_U60 & P3_U2355); 
assign P3_U5690 = ~(P3_ADD_494_U71 & P3_U2356); 
assign P3_U5691 = ~(P3_ADD_476_U71 & P3_U4303); 
assign P3_U5692 = ~(P3_ADD_441_U71 & P3_U4304); 
assign P3_U5694 = ~(P3_ADD_394_U5 & P3_U2357); 
assign P3_U5696 = ~(P3_ADD_380_U74 & P3_U2359); 
assign P3_U5711 = ~(P3_ADD_531_U71 & P3_U2354); 
assign P3_U5712 = ~(P3_ADD_526_U57 & P3_U2355); 
assign P3_U5714 = ~(P3_ADD_494_U68 & P3_U2356); 
assign P3_U5715 = ~(P3_ADD_476_U68 & P3_U4303); 
assign P3_U5716 = ~(P3_ADD_441_U68 & P3_U4304); 
assign P3_U5718 = ~(P3_ADD_394_U93 & P3_U2357); 
assign P3_U5720 = ~(P3_ADD_380_U71 & P3_U2359); 
assign P3_U5735 = ~(P3_ADD_531_U70 & P3_U2354); 
assign P3_U5736 = ~(P3_ADD_526_U56 & P3_U2355); 
assign P3_U5738 = ~(P3_ADD_494_U67 & P3_U2356); 
assign P3_U5739 = ~(P3_ADD_476_U67 & P3_U4303); 
assign P3_U5740 = ~(P3_ADD_441_U67 & P3_U4304); 
assign P3_U5742 = ~(P3_ADD_394_U68 & P3_U2357); 
assign P3_U5744 = ~(P3_ADD_380_U70 & P3_U2359); 
assign P3_U5759 = ~(P3_ADD_531_U69 & P3_U2354); 
assign P3_U5760 = ~(P3_ADD_526_U55 & P3_U2355); 
assign P3_U5762 = ~(P3_ADD_494_U66 & P3_U2356); 
assign P3_U5763 = ~(P3_ADD_476_U66 & P3_U4303); 
assign P3_U5764 = ~(P3_ADD_441_U66 & P3_U4304); 
assign P3_U5766 = ~(P3_ADD_394_U67 & P3_U2357); 
assign P3_U5768 = ~(P3_ADD_380_U69 & P3_U2359); 
assign P3_U5783 = ~(P3_ADD_531_U68 & P3_U2354); 
assign P3_U5784 = ~(P3_ADD_526_U54 & P3_U2355); 
assign P3_U5786 = ~(P3_ADD_494_U65 & P3_U2356); 
assign P3_U5787 = ~(P3_ADD_476_U65 & P3_U4303); 
assign P3_U5788 = ~(P3_ADD_441_U65 & P3_U4304); 
assign P3_U5790 = ~(P3_ADD_394_U66 & P3_U2357); 
assign P3_U5792 = ~(P3_ADD_380_U68 & P3_U2359); 
assign P3_U5808 = ~(P3_ADD_526_U53 & P3_U2355); 
assign P3_U5810 = ~(P3_ADD_494_U64 & P3_U2356); 
assign P3_U5811 = ~(P3_ADD_476_U64 & P3_U4303); 
assign P3_U5812 = ~(P3_ADD_441_U64 & P3_U4304); 
assign P3_U5814 = ~(P3_ADD_394_U65 & P3_U2357); 
assign P3_U5832 = ~(P3_ADD_526_U52 & P3_U2355); 
assign P3_U5856 = ~(P3_ADD_526_U51 & P3_U2355); 
assign P3_U5880 = ~(P3_ADD_526_U81 & P3_U2355); 
assign P3_U5904 = ~(P3_ADD_526_U80 & P3_U2355); 
assign P3_U7377 = ~(P3_U7919 & P3_U4150 & P3_STATE2_REG_2__SCAN_IN); 
assign P3_U7969 = ~(P3_U3109 & P3_U3101); 
assign P3_U7970 = ~(P3_U4539 & P3_U5483); 
assign P2_U2361 = P2_R2238_U6 & P2_U2356; 
assign P2_U2514 = P2_U3881 & P2_U7896 & P2_U3882; 
assign P2_U3594 = P2_U3866 & P2_U4434; 
assign P2_U3616 = P2_U4434 & P2_R2147_U7; 
assign P2_U3654 = ~(P2_U8364 & P2_U8363); 
assign P2_U3883 = P2_U5608 & P2_U5607; 
assign P2_U4379 = P2_U7579 & P2_U7580 & P2_U7578; 
assign P2_U4384 = P2_U4383 & P2_U7578; 
assign P2_U4396 = P2_U8092 & P2_U8091; 
assign P2_U4618 = ~(P2_U3711 & P2_U4425); 
assign P2_U5609 = ~(P2_R2147_U8 & P2_U5604); 
assign P2_U5617 = ~(P2_R2147_U9 & P2_U5604); 
assign P2_U5626 = ~(P2_U3887 & P2_U8097); 
assign P2_U5627 = ~(P2_R2147_U4 & P2_U5604); 
assign P2_U5634 = ~(P2_U3889 & P2_U8097); 
assign P2_U5635 = ~(P2_U5604 & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P2_U6852 = ~(P2_U6851 & P2_U6850 & P2_U4186); 
assign P2_U7139 = ~(P2_U7137 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7150 = ~(P2_U7137 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P2_U7161 = ~(P2_U7137 & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P2_U7164 = ~(P2_U7137 & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P2_U7593 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P2_U7595 = ~(P2_U4423 & P2_REIP_REG_9__SCAN_IN); 
assign P2_U7596 = ~(P2_U2358 & P2_EBX_REG_9__SCAN_IN); 
assign P2_U7597 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P2_U7599 = ~(P2_U4423 & P2_REIP_REG_8__SCAN_IN); 
assign P2_U7600 = ~(P2_U2358 & P2_EBX_REG_8__SCAN_IN); 
assign P2_U7601 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P2_U7603 = ~(P2_U4423 & P2_REIP_REG_7__SCAN_IN); 
assign P2_U7604 = ~(P2_U2358 & P2_EBX_REG_7__SCAN_IN); 
assign P2_U7605 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P2_U7607 = ~(P2_U4423 & P2_REIP_REG_6__SCAN_IN); 
assign P2_U7608 = ~(P2_U2358 & P2_EBX_REG_6__SCAN_IN); 
assign P2_U7609 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P2_U7611 = ~(P2_U4423 & P2_REIP_REG_5__SCAN_IN); 
assign P2_U7612 = ~(P2_U2358 & P2_EBX_REG_5__SCAN_IN); 
assign P2_U7613 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P2_U7615 = ~(P2_U4423 & P2_REIP_REG_4__SCAN_IN); 
assign P2_U7616 = ~(P2_U2358 & P2_EBX_REG_4__SCAN_IN); 
assign P2_U7617 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P2_U7619 = ~(P2_U4423 & P2_REIP_REG_31__SCAN_IN); 
assign P2_U7620 = ~(P2_U2358 & P2_EBX_REG_31__SCAN_IN); 
assign P2_U7621 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P2_U7623 = ~(P2_U4423 & P2_REIP_REG_30__SCAN_IN); 
assign P2_U7624 = ~(P2_U2358 & P2_EBX_REG_30__SCAN_IN); 
assign P2_U7625 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P2_U7627 = ~(P2_U4423 & P2_REIP_REG_3__SCAN_IN); 
assign P2_U7628 = ~(P2_U2358 & P2_EBX_REG_3__SCAN_IN); 
assign P2_U7629 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P2_U7631 = ~(P2_U4423 & P2_REIP_REG_29__SCAN_IN); 
assign P2_U7632 = ~(P2_U2358 & P2_EBX_REG_29__SCAN_IN); 
assign P2_U7633 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P2_U7635 = ~(P2_U4423 & P2_REIP_REG_28__SCAN_IN); 
assign P2_U7636 = ~(P2_U2358 & P2_EBX_REG_28__SCAN_IN); 
assign P2_U7637 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P2_U7639 = ~(P2_U4423 & P2_REIP_REG_27__SCAN_IN); 
assign P2_U7640 = ~(P2_U2358 & P2_EBX_REG_27__SCAN_IN); 
assign P2_U7641 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P2_U7643 = ~(P2_U4423 & P2_REIP_REG_26__SCAN_IN); 
assign P2_U7644 = ~(P2_U2358 & P2_EBX_REG_26__SCAN_IN); 
assign P2_U7645 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P2_U7647 = ~(P2_U4423 & P2_REIP_REG_25__SCAN_IN); 
assign P2_U7648 = ~(P2_U2358 & P2_EBX_REG_25__SCAN_IN); 
assign P2_U7649 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P2_U7651 = ~(P2_U4423 & P2_REIP_REG_24__SCAN_IN); 
assign P2_U7652 = ~(P2_U2358 & P2_EBX_REG_24__SCAN_IN); 
assign P2_U7653 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P2_U7655 = ~(P2_U4423 & P2_REIP_REG_23__SCAN_IN); 
assign P2_U7656 = ~(P2_U2358 & P2_EBX_REG_23__SCAN_IN); 
assign P2_U7657 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P2_U7659 = ~(P2_U4423 & P2_REIP_REG_22__SCAN_IN); 
assign P2_U7660 = ~(P2_U2358 & P2_EBX_REG_22__SCAN_IN); 
assign P2_U7661 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P2_U7663 = ~(P2_U4423 & P2_REIP_REG_21__SCAN_IN); 
assign P2_U7664 = ~(P2_U2358 & P2_EBX_REG_21__SCAN_IN); 
assign P2_U7665 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P2_U7667 = ~(P2_U4423 & P2_REIP_REG_20__SCAN_IN); 
assign P2_U7668 = ~(P2_U2358 & P2_EBX_REG_20__SCAN_IN); 
assign P2_U7669 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P2_U7671 = ~(P2_U4423 & P2_REIP_REG_2__SCAN_IN); 
assign P2_U7672 = ~(P2_U2358 & P2_EBX_REG_2__SCAN_IN); 
assign P2_U7673 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P2_U7675 = ~(P2_U4423 & P2_REIP_REG_19__SCAN_IN); 
assign P2_U7676 = ~(P2_U2358 & P2_EBX_REG_19__SCAN_IN); 
assign P2_U7677 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P2_U7679 = ~(P2_U4423 & P2_REIP_REG_18__SCAN_IN); 
assign P2_U7680 = ~(P2_U2358 & P2_EBX_REG_18__SCAN_IN); 
assign P2_U7681 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P2_U7683 = ~(P2_U4423 & P2_REIP_REG_17__SCAN_IN); 
assign P2_U7684 = ~(P2_U2358 & P2_EBX_REG_17__SCAN_IN); 
assign P2_U7685 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P2_U7687 = ~(P2_U4423 & P2_REIP_REG_16__SCAN_IN); 
assign P2_U7688 = ~(P2_U2358 & P2_EBX_REG_16__SCAN_IN); 
assign P2_U7689 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P2_U7691 = ~(P2_U4423 & P2_REIP_REG_15__SCAN_IN); 
assign P2_U7692 = ~(P2_U2358 & P2_EBX_REG_15__SCAN_IN); 
assign P2_U7693 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P2_U7695 = ~(P2_U4423 & P2_REIP_REG_14__SCAN_IN); 
assign P2_U7696 = ~(P2_U2358 & P2_EBX_REG_14__SCAN_IN); 
assign P2_U7697 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P2_U7699 = ~(P2_U4423 & P2_REIP_REG_13__SCAN_IN); 
assign P2_U7700 = ~(P2_U2358 & P2_EBX_REG_13__SCAN_IN); 
assign P2_U7701 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P2_U7703 = ~(P2_U4423 & P2_REIP_REG_12__SCAN_IN); 
assign P2_U7704 = ~(P2_U2358 & P2_EBX_REG_12__SCAN_IN); 
assign P2_U7705 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P2_U7707 = ~(P2_U4423 & P2_REIP_REG_11__SCAN_IN); 
assign P2_U7708 = ~(P2_U2358 & P2_EBX_REG_11__SCAN_IN); 
assign P2_U7709 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P2_U7711 = ~(P2_U4423 & P2_REIP_REG_10__SCAN_IN); 
assign P2_U7712 = ~(P2_U2358 & P2_EBX_REG_10__SCAN_IN); 
assign P2_U7713 = ~(P2_U7592 & P2_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P2_U7715 = ~(P2_U4423 & P2_REIP_REG_1__SCAN_IN); 
assign P2_U7716 = ~(P2_U2358 & P2_EBX_REG_1__SCAN_IN); 
assign P2_U7718 = ~(P2_U7739 & P2_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P2_U7720 = ~(P2_U4423 & P2_REIP_REG_0__SCAN_IN); 
assign P2_U7721 = ~(P2_U2358 & P2_EBX_REG_0__SCAN_IN); 
assign P2_U7726 = ~(P2_R2238_U19 & P2_U2356); 
assign P2_U8351 = ~(P2_R2238_U6 & P2_U3283); 
assign P2_U8352 = ~(P2_SUB_450_U6 & P2_U4417); 
assign P2_U8353 = ~(P2_R2238_U19 & P2_U3283); 
assign P2_U8354 = ~(P2_SUB_450_U17 & P2_U4417); 
assign P2_U8423 = ~(P2_R2238_U6 & P2_U3269); 
assign P2_U8425 = ~(P2_R2238_U19 & P2_U3269); 
assign P1_U2356 = P1_R2238_U6 & P1_U4192; 
assign P1_U2718 = ~(P1_U4161 & P1_U7368); 
assign P1_U2731 = ~(P1_U2606 & P1_U7354); 
assign P1_U2751 = ~(P1_U4061 & P1_U7058); 
assign P1_U3747 = P1_U3748 & P1_U5502; 
assign P1_U3749 = P1_U7717 & P1_U7716 & P1_U5513; 
assign P1_U3750 = P1_U5524 & P1_U5522; 
assign P1_U3758 = P1_U2520 & P1_U5568 & P1_U3757; 
assign P1_U3762 = P1_U7508 & P1_STATE2_REG_2__SCAN_IN; 
assign P1_U4004 = P1_U6755 & P1_U6754; 
assign P1_U4075 = P1_U7472 & P1_U3434 & P1_U7473; 
assign P1_U4077 = P1_U2606 & P1_U7477 & P1_U4076; 
assign P1_U4113 = P1_U4112 & P1_U7472 & P1_U7473; 
assign P1_U4118 = P1_U7472 & P1_U3434 & P1_U7473; 
assign P1_U4120 = P1_U2608 & P1_U7477 & P1_U2606 & P1_U4119; 
assign P1_U4175 = P1_U7726 & P1_U7725; 
assign P1_U4198 = ~P1_U3425; 
assign P1_U6609 = ~(P1_U3965 & P1_U6607); 
assign P1_U6884 = ~(P1_ADD_371_U5 & P1_U4208); 
assign P1_U6887 = ~(P1_ADD_371_U20 & P1_U4208); 
assign P1_U6927 = ~(P1_U4207 & P1_U3234); 
assign P1_U6929 = ~(P1_U4207 & P1_U3233); 
assign P1_U6931 = ~(P1_U4207 & P1_U3232); 
assign P1_U6933 = ~(P1_U4207 & P1_U3231); 
assign P1_U6935 = ~(P1_U4207 & P1_U3230); 
assign P1_U6938 = ~(P1_U4207 & P1_U3229); 
assign P1_U7041 = ~(P1_U4207 & P1_U3228); 
assign P1_U7044 = ~(P1_U4207 & P1_U3227); 
assign P1_U7083 = ~(P1_U3425 & P1_U3421); 
assign P1_U7093 = ~(P1_U4194 & P1_U7092); 
assign P1_U7359 = ~(P1_U7355 & P1_U3271); 
assign P1_U7364 = ~(P1_R2238_U6 & P1_U7363); 
assign P1_U7365 = ~(P1_SUB_450_U6 & P1_U2354); 
assign P1_U7366 = ~(P1_R2238_U19 & P1_U7363); 
assign P1_U7367 = ~(P1_SUB_450_U19 & P1_U2354); 
assign P1_U7376 = ~(P1_R2238_U19 & P1_U4192); 
assign P1_U7487 = ~(P1_U7091 & P1_U4194); 
assign P1_U7707 = ~(P1_U7706 & P1_U7705); 
assign P3_ADD_526_U78 = ~(P3_ADD_526_U196 & P3_ADD_526_U195); 
assign P3_ADD_526_U79 = ~(P3_ADD_526_U198 & P3_ADD_526_U197); 
assign P3_ADD_526_U124 = ~P3_ADD_526_U27; 
assign P3_ADD_526_U138 = ~P3_ADD_526_U108; 
assign P3_ADD_526_U192 = ~(P3_ADD_526_U27 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_526_U193 = ~(P3_ADD_526_U108 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_552_U78 = ~(P3_ADD_552_U196 & P3_ADD_552_U195); 
assign P3_ADD_552_U79 = ~(P3_ADD_552_U198 & P3_ADD_552_U197); 
assign P3_ADD_552_U124 = ~P3_ADD_552_U27; 
assign P3_ADD_552_U138 = ~P3_ADD_552_U108; 
assign P3_ADD_552_U192 = ~(P3_ADD_552_U27 & P3_EBX_REG_15__SCAN_IN); 
assign P3_ADD_552_U193 = ~(P3_ADD_552_U108 & P3_EBX_REG_14__SCAN_IN); 
assign P3_ADD_546_U78 = ~(P3_ADD_546_U196 & P3_ADD_546_U195); 
assign P3_ADD_546_U79 = ~(P3_ADD_546_U198 & P3_ADD_546_U197); 
assign P3_ADD_546_U124 = ~P3_ADD_546_U27; 
assign P3_ADD_546_U138 = ~P3_ADD_546_U108; 
assign P3_ADD_546_U192 = ~(P3_ADD_546_U27 & P3_EAX_REG_15__SCAN_IN); 
assign P3_ADD_546_U193 = ~(P3_ADD_546_U108 & P3_EAX_REG_14__SCAN_IN); 
assign P3_GTE_401_U8 = ~(P3_SUB_401_U19 | P3_SUB_401_U20 | P3_GTE_401_U7); 
assign P3_ADD_391_1180_U8 = ~(P3_U2614 & P3_ADD_391_1180_U28); 
assign P3_ADD_391_1180_U25 = ~(P3_ADD_391_1180_U50 & P3_ADD_391_1180_U49); 
assign P3_ADD_391_1180_U48 = ~(P3_ADD_391_1180_U28 & P3_ADD_391_1180_U7); 
assign P3_ADD_476_U63 = ~(P3_ADD_476_U126 & P3_ADD_476_U125); 
assign P3_ADD_476_U100 = ~P3_ADD_476_U19; 
assign P3_ADD_476_U123 = ~(P3_ADD_476_U19 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_GTE_390_U8 = ~(P3_SUB_390_U19 | P3_SUB_390_U20 | P3_GTE_390_U7); 
assign P3_ADD_531_U67 = ~(P3_ADD_531_U133 & P3_ADD_531_U132); 
assign P3_ADD_531_U104 = ~P3_ADD_531_U19; 
assign P3_ADD_531_U130 = ~(P3_ADD_531_U19 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_SUB_320_U87 = ~(P3_SUB_320_U85 & P3_SUB_320_U54); 
assign P3_SUB_320_U131 = ~(P3_SUB_320_U85 & P3_SUB_320_U54); 
assign P3_GTE_485_U7 = ~(P3_SUB_485_U16 | P3_SUB_485_U17 | P3_SUB_485_U19 | P3_SUB_485_U18); 
assign P3_ADD_318_U63 = ~(P3_ADD_318_U126 & P3_ADD_318_U125); 
assign P3_ADD_318_U100 = ~P3_ADD_318_U19; 
assign P3_ADD_318_U123 = ~(P3_ADD_318_U19 & P3_PHYADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_315_U60 = ~(P3_ADD_315_U120 & P3_ADD_315_U119); 
assign P3_ADD_315_U97 = ~P3_ADD_315_U18; 
assign P3_ADD_315_U175 = ~(P3_ADD_315_U18 & P3_PHYADDRPOINTER_REG_10__SCAN_IN); 
assign P3_GTE_355_U8 = ~(P3_SUB_355_U19 | P3_SUB_355_U20 | P3_GTE_355_U7 | P3_SUB_355_U21); 
assign P3_ADD_360_1242_U75 = ~(P3_ADD_360_U4 & P3_ADD_360_1242_U124); 
assign P3_ADD_360_1242_U85 = ~(P3_ADD_360_1242_U258 & P3_ADD_360_1242_U257); 
assign P3_ADD_360_1242_U126 = ~(P3_ADD_360_1242_U28 & P3_ADD_360_1242_U27); 
assign P3_ADD_360_1242_U245 = ~(P3_ADD_360_1242_U124 & P3_ADD_360_1242_U26); 
assign P3_ADD_467_U63 = ~(P3_ADD_467_U126 & P3_ADD_467_U125); 
assign P3_ADD_467_U100 = ~P3_ADD_467_U19; 
assign P3_ADD_467_U123 = ~(P3_ADD_467_U19 & P3_REIP_REG_9__SCAN_IN); 
assign P3_ADD_430_U63 = ~(P3_ADD_430_U126 & P3_ADD_430_U125); 
assign P3_ADD_430_U100 = ~P3_ADD_430_U19; 
assign P3_ADD_430_U123 = ~(P3_ADD_430_U19 & P3_REIP_REG_9__SCAN_IN); 
assign P3_ADD_380_U67 = ~(P3_ADD_380_U133 & P3_ADD_380_U132); 
assign P3_ADD_380_U104 = ~P3_ADD_380_U19; 
assign P3_ADD_380_U130 = ~(P3_ADD_380_U19 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_GTE_370_U8 = ~(P3_SUB_370_U19 | P3_GTE_370_U7 | P3_SUB_370_U20); 
assign P3_ADD_344_U67 = ~(P3_ADD_344_U133 & P3_ADD_344_U132); 
assign P3_ADD_344_U104 = ~P3_ADD_344_U19; 
assign P3_ADD_344_U130 = ~(P3_ADD_344_U19 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_339_U63 = ~(P3_ADD_339_U126 & P3_ADD_339_U125); 
assign P3_ADD_339_U100 = ~P3_ADD_339_U19; 
assign P3_ADD_339_U123 = ~(P3_ADD_339_U19 & P3_PHYADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_360_U9 = ~(P3_U2624 & P3_ADD_360_U24); 
assign P3_ADD_360_U21 = ~(P3_ADD_360_U40 & P3_ADD_360_U39); 
assign P3_ADD_360_U38 = ~(P3_ADD_360_U24 & P3_ADD_360_U8); 
assign P3_ADD_541_U63 = ~(P3_ADD_541_U126 & P3_ADD_541_U125); 
assign P3_ADD_541_U100 = ~P3_ADD_541_U19; 
assign P3_ADD_541_U123 = ~(P3_ADD_541_U19 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_SUB_357_1258_U28 = ~P3_ADD_357_U10; 
assign P3_SUB_357_1258_U30 = ~(P3_ADD_357_U10 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_SUB_357_1258_U484 = ~(P3_ADD_357_U10 & P3_SUB_357_1258_U29); 
assign P3_ADD_515_U63 = ~(P3_ADD_515_U126 & P3_ADD_515_U125); 
assign P3_ADD_515_U100 = ~P3_ADD_515_U19; 
assign P3_ADD_515_U123 = ~(P3_ADD_515_U19 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_394_U64 = ~(P3_ADD_394_U130 & P3_ADD_394_U129); 
assign P3_ADD_394_U103 = ~P3_ADD_394_U19; 
assign P3_ADD_394_U127 = ~(P3_ADD_394_U19 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_GTE_450_U7 = ~(P3_SUB_450_U16 | P3_SUB_450_U17 | P3_SUB_450_U19 | P3_SUB_450_U18); 
assign P3_SUB_414_U80 = P3_SUB_414_U157 & P3_SUB_414_U156; 
assign P3_SUB_414_U95 = ~P3_SUB_414_U30; 
assign P3_SUB_414_U122 = ~(P3_SUB_414_U121 & P3_EBX_REG_14__SCAN_IN); 
assign P3_SUB_414_U154 = ~(P3_SUB_414_U30 & P3_EBX_REG_15__SCAN_IN); 
assign P3_ADD_441_U63 = ~(P3_ADD_441_U126 & P3_ADD_441_U125); 
assign P3_ADD_441_U100 = ~P3_ADD_441_U19; 
assign P3_ADD_441_U123 = ~(P3_ADD_441_U19 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_349_U67 = ~(P3_ADD_349_U133 & P3_ADD_349_U132); 
assign P3_ADD_349_U104 = ~P3_ADD_349_U19; 
assign P3_ADD_349_U130 = ~(P3_ADD_349_U19 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_405_U64 = ~(P3_ADD_405_U130 & P3_ADD_405_U129); 
assign P3_ADD_405_U103 = ~P3_ADD_405_U19; 
assign P3_ADD_405_U127 = ~(P3_ADD_405_U19 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_553_U67 = ~(P3_ADD_553_U133 & P3_ADD_553_U132); 
assign P3_ADD_553_U104 = ~P3_ADD_553_U19; 
assign P3_ADD_553_U130 = ~(P3_ADD_553_U19 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_558_U67 = ~(P3_ADD_558_U133 & P3_ADD_558_U132); 
assign P3_ADD_558_U104 = ~P3_ADD_558_U19; 
assign P3_ADD_558_U130 = ~(P3_ADD_558_U19 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_385_U67 = ~(P3_ADD_385_U133 & P3_ADD_385_U132); 
assign P3_ADD_385_U104 = ~P3_ADD_385_U19; 
assign P3_ADD_385_U130 = ~(P3_ADD_385_U19 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_357_U22 = ~P3_ADD_357_U11; 
assign P3_ADD_357_U29 = ~(P3_SUB_357_U11 & P3_ADD_357_U28); 
assign P3_ADD_357_U32 = ~(P3_SUB_357_U13 & P3_ADD_357_U11); 
assign P3_ADD_357_U34 = ~(P3_SUB_357_U7 & P3_ADD_357_U21); 
assign P3_ADD_357_U35 = ~(P3_SUB_357_U12 & P3_ADD_357_U20); 
assign P3_ADD_547_U67 = ~(P3_ADD_547_U133 & P3_ADD_547_U132); 
assign P3_ADD_547_U104 = ~P3_ADD_547_U19; 
assign P3_ADD_547_U130 = ~(P3_ADD_547_U19 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_371_1212_U121 = ~P3_ADD_371_1212_U34; 
assign P3_ADD_371_1212_U251 = ~(P3_ADD_371_1212_U34 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_371_1212_U264 = ~(P3_ADD_371_1212_U31 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_ADD_371_U5 = ~(P3_ADD_371_U24 & P3_ADD_371_U32); 
assign P3_ADD_371_U9 = ~(P3_U2624 & P3_ADD_371_U24); 
assign P3_ADD_371_U21 = ~(P3_ADD_371_U44 & P3_ADD_371_U43); 
assign P3_ADD_371_U27 = ~P3_ADD_371_U24; 
assign P3_ADD_371_U41 = ~(P3_U2624 & P3_ADD_371_U24); 
assign P3_GTE_412_U7 = ~(P3_SUB_412_U16 | P3_SUB_412_U17 | P3_SUB_412_U19 | P3_SUB_412_U18); 
assign P3_GTE_504_U7 = ~(P3_SUB_504_U16 | P3_SUB_504_U17 | P3_SUB_504_U19 | P3_SUB_504_U18); 
assign P3_ADD_494_U63 = ~(P3_ADD_494_U126 & P3_ADD_494_U125); 
assign P3_ADD_494_U100 = ~P3_ADD_494_U19; 
assign P3_ADD_494_U123 = ~(P3_ADD_494_U19 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_536_U63 = ~(P3_ADD_536_U126 & P3_ADD_536_U125); 
assign P3_ADD_536_U100 = ~P3_ADD_536_U19; 
assign P3_ADD_536_U123 = ~(P3_ADD_536_U19 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_402_1132_U8 = ~(P3_U2614 & P3_ADD_402_1132_U28); 
assign P3_ADD_402_1132_U25 = ~(P3_ADD_402_1132_U50 & P3_ADD_402_1132_U49); 
assign P3_ADD_402_1132_U48 = ~(P3_ADD_402_1132_U28 & P3_ADD_402_1132_U7); 
assign P2_ADD_402_1132_U8 = ~(P2_U2592 & P2_ADD_402_1132_U28); 
assign P2_ADD_402_1132_U23 = ~(P2_ADD_402_1132_U46 & P2_ADD_402_1132_U45); 
assign P2_ADD_402_1132_U40 = ~(P2_ADD_402_1132_U28 & P2_ADD_402_1132_U7); 
assign P2_R2182_U27 = ~P2_U2696; 
assign P2_R2182_U28 = ~P2_U2695; 
assign P2_R2182_U29 = ~P2_U2694; 
assign P2_R2182_U30 = ~P2_U2693; 
assign P2_R2182_U31 = ~P2_U2692; 
assign P2_R2182_U32 = ~P2_U2691; 
assign P2_R2182_U37 = ~P2_U2690; 
assign P2_R2182_U203 = ~(P2_U2677 & P2_R2182_U50); 
assign P2_R2182_U205 = ~(P2_U2677 & P2_R2182_U50); 
assign P2_R2167_U11 = ~P2_U2704; 
assign P2_R2027_U67 = ~(P2_R2027_U133 & P2_R2027_U132); 
assign P2_R2027_U104 = ~P2_R2027_U19; 
assign P2_R2027_U130 = ~(P2_R2027_U19 & P2_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P2_R2337_U61 = ~(P2_R2337_U124 & P2_R2337_U123); 
assign P2_R2337_U101 = ~P2_R2337_U19; 
assign P2_R2337_U181 = ~(P2_R2337_U19 & P2_PHYADDRPOINTER_REG_10__SCAN_IN); 
assign P2_R2219_U10 = ~P2_U2753; 
assign P2_R2219_U11 = ~P2_U2761; 
assign P2_R2219_U12 = ~P2_U2763; 
assign P2_R2219_U13 = ~P2_U2762; 
assign P2_R2219_U14 = ~P2_U2756; 
assign P2_R2219_U15 = ~P2_U2765; 
assign P2_R2219_U16 = ~P2_U2764; 
assign P2_R2219_U17 = ~P2_U2755; 
assign P2_R2219_U18 = ~P2_U2754; 
assign P2_R2219_U23 = ~P2_U2757; 
assign P2_R2219_U32 = ~(P2_R2219_U83 & P2_R2219_U82); 
assign P2_R2219_U33 = ~(P2_R2219_U88 & P2_R2219_U87); 
assign P2_R2219_U34 = ~(P2_R2219_U93 & P2_R2219_U92); 
assign P2_R2096_U26 = ~P2_U2631; 
assign P2_R2096_U27 = ~P2_U2638; 
assign P2_R2096_U28 = ~P2_U2640; 
assign P2_R2096_U29 = ~P2_U2618; 
assign P2_R2096_U30 = ~P2_U2619; 
assign P2_R2096_U31 = ~P2_U2635; 
assign P2_R2096_U32 = ~P2_U2636; 
assign P2_R2096_U33 = ~P2_U2637; 
assign P2_R2096_U34 = ~P2_U2633; 
assign P2_R2096_U35 = ~P2_U2634; 
assign P2_R2096_U36 = ~P2_U2629; 
assign P2_R2096_U37 = ~P2_U2641; 
assign P2_R2096_U38 = ~P2_U2622; 
assign P2_R2096_U39 = ~P2_U2627; 
assign P2_R2096_U40 = ~P2_U2620; 
assign P2_R2096_U41 = ~P2_U2621; 
assign P2_R2096_U42 = ~P2_U2623; 
assign P2_R2096_U43 = ~P2_U2624; 
assign P2_R2096_U44 = ~P2_U2625; 
assign P2_R2096_U45 = ~P2_U2626; 
assign P2_R2096_U46 = ~P2_U2628; 
assign P2_R2096_U47 = ~P2_U2630; 
assign P2_R2096_U48 = ~P2_U2632; 
assign P2_R2096_U49 = ~P2_U2639; 
assign P2_R2096_U53 = ~P2_U2649; 
assign P2_R2096_U54 = ~P2_U2648; 
assign P2_R2096_U57 = ~P2_U2647; 
assign P2_R2096_U59 = ~P2_U2646; 
assign P2_R2096_U61 = ~P2_U2645; 
assign P2_R2096_U63 = ~P2_U2644; 
assign P2_R2096_U65 = ~P2_U2643; 
assign P2_R2096_U67 = ~P2_U2642; 
assign P2_R2096_U98 = P2_U2619 & P2_U2618; 
assign P2_R2096_U112 = ~(P2_U2649 & P2_U2657); 
assign P2_R2096_U113 = ~(P2_U2649 & P2_U2657 & P2_U2656); 
assign P2_R2096_U116 = ~(P2_U2649 & P2_U2657); 
assign P2_R2096_U120 = P2_U2655 | P2_U2647; 
assign P2_R2096_U122 = ~(P2_U2647 & P2_U2655); 
assign P2_R2096_U124 = P2_U2654 | P2_U2646; 
assign P2_R2096_U126 = ~(P2_U2646 & P2_U2654); 
assign P2_R2096_U128 = P2_U2653 | P2_U2645; 
assign P2_R2096_U130 = ~(P2_U2645 & P2_U2653); 
assign P2_R2096_U132 = P2_U2652 | P2_U2644; 
assign P2_R2096_U134 = ~(P2_U2644 & P2_U2652); 
assign P2_R2096_U136 = P2_U2651 | P2_U2643; 
assign P2_R2096_U138 = ~(P2_U2643 & P2_U2651); 
assign P2_R2096_U140 = P2_U2650 | P2_U2642; 
assign P2_R2096_U142 = ~(P2_U2642 & P2_U2650); 
assign P2_R2096_U175 = ~(P2_U2642 & P2_R2096_U66); 
assign P2_R2096_U177 = ~(P2_U2642 & P2_R2096_U66); 
assign P2_R2096_U182 = ~(P2_U2643 & P2_R2096_U64); 
assign P2_R2096_U184 = ~(P2_U2643 & P2_R2096_U64); 
assign P2_R2096_U189 = ~(P2_U2644 & P2_R2096_U62); 
assign P2_R2096_U191 = ~(P2_U2644 & P2_R2096_U62); 
assign P2_R2096_U196 = ~(P2_U2645 & P2_R2096_U60); 
assign P2_R2096_U198 = ~(P2_U2645 & P2_R2096_U60); 
assign P2_R2096_U203 = ~(P2_U2646 & P2_R2096_U58); 
assign P2_R2096_U205 = ~(P2_U2646 & P2_R2096_U58); 
assign P2_R2096_U212 = ~(P2_U2647 & P2_R2096_U56); 
assign P2_R2096_U214 = ~(P2_U2647 & P2_R2096_U56); 
assign P2_R2096_U264 = ~(P2_U2649 & P2_R2096_U52); 
assign P2_R1957_U87 = ~(P2_R1957_U85 & P2_R1957_U54); 
assign P2_R1957_U131 = ~(P2_R1957_U85 & P2_R1957_U54); 
assign P2_ADD_394_U80 = ~(P2_ADD_394_U162 & P2_ADD_394_U161); 
assign P2_ADD_394_U103 = ~P2_ADD_394_U18; 
assign P2_ADD_394_U141 = ~(P2_ADD_394_U18 & P2_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P1_R2027_U78 = ~(P1_R2027_U196 & P1_R2027_U195); 
assign P1_R2027_U79 = ~(P1_R2027_U198 & P1_R2027_U197); 
assign P1_R2027_U124 = ~P1_R2027_U27; 
assign P1_R2027_U138 = ~P1_R2027_U108; 
assign P1_R2027_U192 = ~(P1_R2027_U27 & P1_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P1_R2027_U193 = ~(P1_R2027_U108 & P1_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P1_R2144_U202 = ~(P1_U2355 & P1_R2144_U76); 
assign P1_R2144_U205 = ~(P1_U2355 & P1_R2144_U77); 
assign P1_R2144_U220 = ~(P1_U2355 & P1_R2144_U85); 
assign P1_R2144_U223 = ~(P1_U2355 & P1_R2144_U86); 
assign P1_R2144_U226 = ~(P1_U2355 & P1_R2144_U87); 
assign P1_R2144_U229 = ~(P1_U2355 & P1_R2144_U88); 
assign P1_R2144_U232 = ~(P1_U2355 & P1_R2144_U89); 
assign P1_R2144_U235 = ~(P1_U2355 & P1_R2144_U90); 
assign P1_R2358_U145 = ~P1_U2614; 
assign P1_R2358_U407 = ~(P1_U2614 & P1_R2358_U23); 
assign P1_R2358_U418 = ~(P1_U2614 & P1_R2358_U23); 
assign P1_R2099_U26 = ~(P1_R2099_U210 & P1_R2099_U209); 
assign P1_R2099_U27 = ~(P1_R2099_U183 & P1_R2099_U182); 
assign P1_R2099_U28 = ~(P1_R2099_U204 & P1_R2099_U203); 
assign P1_R2099_U29 = ~(P1_R2099_U207 & P1_R2099_U206); 
assign P1_R2099_U30 = ~(P1_R2099_U198 & P1_R2099_U197); 
assign P1_R2099_U31 = ~(P1_R2099_U201 & P1_R2099_U200); 
assign P1_R2099_U32 = ~(P1_R2099_U186 & P1_R2099_U185); 
assign P1_R2099_U33 = ~(P1_R2099_U189 & P1_R2099_U188); 
assign P1_R2099_U34 = ~(P1_R2099_U195 & P1_R2099_U194); 
assign P1_R2099_U35 = ~(P1_R2099_U192 & P1_R2099_U191); 
assign P1_R2099_U43 = ~(P1_R2099_U284 & P1_R2099_U283); 
assign P1_R2099_U44 = ~(P1_R2099_U287 & P1_R2099_U286); 
assign P1_R2099_U45 = ~(P1_R2099_U227 & P1_R2099_U226); 
assign P1_R2099_U46 = ~(P1_R2099_U230 & P1_R2099_U229); 
assign P1_R2099_U47 = ~(P1_R2099_U233 & P1_R2099_U232); 
assign P1_R2099_U48 = ~(P1_R2099_U236 & P1_R2099_U235); 
assign P1_R2099_U49 = ~(P1_R2099_U239 & P1_R2099_U238); 
assign P1_R2099_U50 = ~(P1_R2099_U242 & P1_R2099_U241); 
assign P1_R2099_U51 = ~(P1_R2099_U245 & P1_R2099_U244); 
assign P1_R2099_U52 = ~(P1_R2099_U248 & P1_R2099_U247); 
assign P1_R2099_U53 = ~(P1_R2099_U251 & P1_R2099_U250); 
assign P1_R2099_U54 = ~(P1_R2099_U254 & P1_R2099_U253); 
assign P1_R2099_U55 = ~(P1_R2099_U257 & P1_R2099_U256); 
assign P1_R2099_U56 = ~(P1_R2099_U278 & P1_R2099_U277); 
assign P1_R2099_U57 = ~(P1_R2099_U281 & P1_R2099_U280); 
assign P1_R2099_U58 = ~(P1_R2099_U272 & P1_R2099_U271); 
assign P1_R2099_U59 = ~(P1_R2099_U275 & P1_R2099_U274); 
assign P1_R2099_U60 = ~(P1_R2099_U266 & P1_R2099_U265); 
assign P1_R2099_U61 = ~(P1_R2099_U269 & P1_R2099_U268); 
assign P1_R2099_U62 = ~(P1_R2099_U260 & P1_R2099_U259); 
assign P1_R2099_U63 = ~(P1_R2099_U263 & P1_R2099_U262); 
assign P1_R2099_U97 = ~(P1_R2099_U290 & P1_R2099_U289); 
assign P1_R2167_U8 = ~P1_U2720; 
assign P1_R2167_U9 = ~P1_U2719; 
assign P1_R2167_U10 = ~P1_U2713; 
assign P1_R2167_U11 = ~P1_U2712; 
assign P1_R2167_U22 = ~P1_U2721; 
assign P1_R2167_U24 = ~(P1_U2715 & P1_R2167_U23); 
assign P1_R2167_U26 = P1_U2721 | P1_U2722; 
assign P1_R2167_U29 = ~(P1_U2720 & P1_R2167_U7); 
assign P1_R2337_U63 = ~(P1_R2337_U126 & P1_R2337_U125); 
assign P1_R2337_U100 = ~P1_R2337_U19; 
assign P1_R2337_U123 = ~(P1_R2337_U19 & P1_PHYADDRPOINTER_REG_9__SCAN_IN); 
assign P1_R2096_U63 = ~(P1_R2096_U126 & P1_R2096_U125); 
assign P1_R2096_U100 = ~P1_R2096_U19; 
assign P1_R2096_U123 = ~(P1_R2096_U19 & P1_REIP_REG_9__SCAN_IN); 
assign P1_ADD_371_U28 = ~P1_ADD_371_U9; 
assign P1_ADD_371_U35 = ~(P1_U3231 & P1_ADD_371_U9); 
assign P1_ADD_371_U40 = ~(P1_ADD_371_U27 & P1_ADD_371_U8); 
assign P1_ADD_405_U80 = ~(P1_ADD_405_U162 & P1_ADD_405_U161); 
assign P1_ADD_405_U103 = ~P1_ADD_405_U18; 
assign P1_ADD_405_U141 = ~(P1_ADD_405_U18 & P1_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P1_GTE_485_U7 = ~(P1_R2238_U19 | P1_R2238_U20 | P1_R2238_U22 | P1_R2238_U21); 
assign P1_ADD_515_U80 = ~(P1_ADD_515_U160 & P1_ADD_515_U159); 
assign P1_ADD_515_U100 = ~P1_ADD_515_U18; 
assign P1_ADD_515_U139 = ~(P1_ADD_515_U18 & P1_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_U2486 = P3_U3271 & P3_U3182; 
assign P3_U2498 = P3_U7968 & P3_U3182; 
assign P3_U2515 = P3_U7970 & P3_U7969 & P3_U5485; 
assign P3_U3222 = ~(P3_U4314 & P3_U3218); 
assign P3_U3226 = ~(P3_U3674 & P3_U2517); 
assign P3_U3231 = ~(P3_U3115 & P3_U5559); 
assign P3_U3243 = ~(P3_U2461 & P3_U4314); 
assign P3_U3362 = P3_U4626 & P3_U3089; 
assign P3_U3441 = P3_U4883 & P3_U4882; 
assign P3_U3443 = P3_U4888 & P3_U4887; 
assign P3_U3445 = P3_U4893 & P3_U4892; 
assign P3_U3447 = P3_U4898 & P3_U4897; 
assign P3_U3449 = P3_U4903 & P3_U4902; 
assign P3_U3451 = P3_U4908 & P3_U4907; 
assign P3_U3453 = P3_U4913 & P3_U4912; 
assign P3_U3455 = P3_U4918 & P3_U4917; 
assign P3_U3459 = P3_U4935 & P3_U4934; 
assign P3_U3461 = P3_U4940 & P3_U4939; 
assign P3_U3463 = P3_U4945 & P3_U4944; 
assign P3_U3465 = P3_U4950 & P3_U4949; 
assign P3_U3467 = P3_U4955 & P3_U4954; 
assign P3_U3469 = P3_U4960 & P3_U4959; 
assign P3_U3471 = P3_U4965 & P3_U4964; 
assign P3_U3473 = P3_U4970 & P3_U4969; 
assign P3_U3477 = P3_U4987 & P3_U4986; 
assign P3_U3479 = P3_U4992 & P3_U4991; 
assign P3_U3481 = P3_U4997 & P3_U4996; 
assign P3_U3483 = P3_U5002 & P3_U5001; 
assign P3_U3485 = P3_U5007 & P3_U5006; 
assign P3_U3487 = P3_U5012 & P3_U5011; 
assign P3_U3489 = P3_U5017 & P3_U5016; 
assign P3_U3491 = P3_U5022 & P3_U5021; 
assign P3_U3494 = P3_U5038 & P3_U5037; 
assign P3_U3496 = P3_U5043 & P3_U5042; 
assign P3_U3498 = P3_U5048 & P3_U5047; 
assign P3_U3500 = P3_U5053 & P3_U5052; 
assign P3_U3502 = P3_U5058 & P3_U5057; 
assign P3_U3504 = P3_U5063 & P3_U5062; 
assign P3_U3506 = P3_U5068 & P3_U5067; 
assign P3_U3508 = P3_U5073 & P3_U5072; 
assign P3_U3529 = P3_U5139 & P3_U5138; 
assign P3_U3531 = P3_U5144 & P3_U5143; 
assign P3_U3533 = P3_U5149 & P3_U5148; 
assign P3_U3535 = P3_U5154 & P3_U5153; 
assign P3_U3537 = P3_U5159 & P3_U5158; 
assign P3_U3539 = P3_U5164 & P3_U5163; 
assign P3_U3541 = P3_U5169 & P3_U5168; 
assign P3_U3543 = P3_U5174 & P3_U5173; 
assign P3_U3547 = P3_U5191 & P3_U5190; 
assign P3_U3549 = P3_U5196 & P3_U5195; 
assign P3_U3551 = P3_U5201 & P3_U5200; 
assign P3_U3553 = P3_U5206 & P3_U5205; 
assign P3_U3555 = P3_U5211 & P3_U5210; 
assign P3_U3557 = P3_U5216 & P3_U5215; 
assign P3_U3559 = P3_U5221 & P3_U5220; 
assign P3_U3561 = P3_U5226 & P3_U5225; 
assign P3_U3565 = P3_U5241 & P3_U5240 & P3_U5243; 
assign P3_U3567 = P3_U5246 & P3_U5245 & P3_U5248; 
assign P3_U3569 = P3_U5251 & P3_U5250 & P3_U5253; 
assign P3_U3571 = P3_U5256 & P3_U5255 & P3_U5258; 
assign P3_U3573 = P3_U5261 & P3_U5260 & P3_U5263; 
assign P3_U3575 = P3_U5266 & P3_U5265 & P3_U5268; 
assign P3_U3577 = P3_U5271 & P3_U5270 & P3_U5273; 
assign P3_U3579 = P3_U5276 & P3_U5275 & P3_U5278; 
assign P3_U3583 = P3_U5292 & P3_U5291 & P3_U5294; 
assign P3_U3585 = P3_U5297 & P3_U5296 & P3_U5299; 
assign P3_U3587 = P3_U5302 & P3_U5301 & P3_U5304; 
assign P3_U3589 = P3_U5307 & P3_U5306 & P3_U5309; 
assign P3_U3591 = P3_U5312 & P3_U5311 & P3_U5314; 
assign P3_U3593 = P3_U5317 & P3_U5316 & P3_U5319; 
assign P3_U3595 = P3_U5322 & P3_U5321 & P3_U5324; 
assign P3_U3597 = P3_U5327 & P3_U5326 & P3_U5329; 
assign P3_U3600 = P3_U5343 & P3_U5342 & P3_U5345; 
assign P3_U3602 = P3_U5348 & P3_U5347 & P3_U5350; 
assign P3_U3604 = P3_U5353 & P3_U5352 & P3_U5355; 
assign P3_U3606 = P3_U5358 & P3_U5357 & P3_U5360; 
assign P3_U3608 = P3_U5363 & P3_U5362 & P3_U5365; 
assign P3_U3610 = P3_U5368 & P3_U5367 & P3_U5370; 
assign P3_U3612 = P3_U5373 & P3_U5372 & P3_U5375; 
assign P3_U3614 = P3_U5378 & P3_U5377 & P3_U5380; 
assign P3_U3618 = P3_U5394 & P3_U5393 & P3_U5396; 
assign P3_U3620 = P3_U5399 & P3_U5398 & P3_U5401; 
assign P3_U3622 = P3_U5404 & P3_U5403 & P3_U5406; 
assign P3_U3624 = P3_U5409 & P3_U5408 & P3_U5411; 
assign P3_U3626 = P3_U5414 & P3_U5413 & P3_U5416; 
assign P3_U3628 = P3_U5419 & P3_U5418 & P3_U5421; 
assign P3_U3630 = P3_U5424 & P3_U5423 & P3_U5426; 
assign P3_U3632 = P3_U5429 & P3_U5428 & P3_U5431; 
assign P3_U3636 = P3_U5444 & P3_U5443 & P3_U5446; 
assign P3_U3638 = P3_U5449 & P3_U5448 & P3_U5451; 
assign P3_U3640 = P3_U5454 & P3_U5453 & P3_U5456; 
assign P3_U3642 = P3_U5459 & P3_U5458 & P3_U5461; 
assign P3_U3644 = P3_U5464 & P3_U5463 & P3_U5466; 
assign P3_U3646 = P3_U5469 & P3_U5468 & P3_U5471; 
assign P3_U3648 = P3_U5474 & P3_U5473 & P3_U5476; 
assign P3_U3650 = P3_U5479 & P3_U5478 & P3_U5481; 
assign P3_U3668 = P3_U5528 & P3_U3242 & P3_U2517; 
assign P3_U3678 = P3_U5552 & P3_U5550; 
assign P3_U3695 = P3_U5639 & P3_U5640; 
assign P3_U3702 = P3_U5663 & P3_U5664; 
assign P3_U3709 = P3_U5687 & P3_U5688; 
assign P3_U3717 = P3_U5711 & P3_U5712; 
assign P3_U3725 = P3_U5735 & P3_U5736; 
assign P3_U3733 = P3_U5759 & P3_U5760; 
assign P3_U3741 = P3_U5783 & P3_U5784; 
assign P3_U4660 = ~P3_U3182; 
assign P3_U5087 = ~(P3_U4326 & P3_U2436); 
assign P3_U5092 = ~(P3_U4326 & P3_U2434); 
assign P3_U5097 = ~(P3_U4326 & P3_U2432); 
assign P3_U5102 = ~(P3_U4326 & P3_U2430); 
assign P3_U5107 = ~(P3_U4326 & P3_U2428); 
assign P3_U5112 = ~(P3_U4326 & P3_U2426); 
assign P3_U5117 = ~(P3_U4326 & P3_U2424); 
assign P3_U5122 = ~(P3_U4326 & P3_U2422); 
assign P3_U5509 = ~(P3_U4296 & P3_U5507); 
assign P3_U5579 = ~P3_U3233; 
assign P3_U5581 = ~(P3_U3233 & P3_U5580); 
assign P3_U5584 = ~(P3_U3182 & P3_U5583); 
assign P3_U5595 = ~(P3_U3686 & P3_U5593); 
assign P3_U5597 = ~(P3_U3233 & P3_U5596); 
assign P3_U5608 = ~(P3_U3233 & P3_U5607); 
assign P3_U5610 = ~(P3_U5606 & P3_U3233); 
assign P3_U5612 = ~(P3_U5611 & P3_U3233); 
assign P3_U5614 = ~(P3_U4337 & P3_U5613); 
assign P3_U5632 = ~(P3_ADD_360_1242_U85 & P3_U2395); 
assign P3_U5635 = ~(P3_U4298 & P3_ADD_553_U5); 
assign P3_U5641 = ~(P3_U4302 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_U5645 = ~(P3_ADD_405_U4 & P3_U4305); 
assign P3_U5647 = ~(P3_U2358 & P3_ADD_385_U5); 
assign P3_U5649 = ~(P3_U4306 & P3_ADD_349_U5); 
assign P3_U5650 = ~(P3_U2362 & P3_ADD_344_U5); 
assign P3_U5659 = ~(P3_ADD_553_U85 & P3_U4298); 
assign P3_U5665 = ~(P3_ADD_515_U4 & P3_U4302); 
assign P3_U5669 = ~(P3_ADD_405_U81 & P3_U4305); 
assign P3_U5671 = ~(P3_ADD_385_U85 & P3_U2358); 
assign P3_U5673 = ~(P3_ADD_349_U85 & P3_U4306); 
assign P3_U5674 = ~(P3_ADD_344_U85 & P3_U2362); 
assign P3_U5683 = ~(P3_ADD_553_U74 & P3_U4298); 
assign P3_U5689 = ~(P3_ADD_515_U71 & P3_U4302); 
assign P3_U5693 = ~(P3_ADD_405_U5 & P3_U4305); 
assign P3_U5695 = ~(P3_ADD_385_U74 & P3_U2358); 
assign P3_U5697 = ~(P3_ADD_349_U74 & P3_U4306); 
assign P3_U5698 = ~(P3_ADD_344_U74 & P3_U2362); 
assign P3_U5707 = ~(P3_ADD_553_U71 & P3_U4298); 
assign P3_U5713 = ~(P3_ADD_515_U68 & P3_U4302); 
assign P3_U5717 = ~(P3_ADD_405_U93 & P3_U4305); 
assign P3_U5719 = ~(P3_ADD_385_U71 & P3_U2358); 
assign P3_U5721 = ~(P3_ADD_349_U71 & P3_U4306); 
assign P3_U5722 = ~(P3_ADD_344_U71 & P3_U2362); 
assign P3_U5731 = ~(P3_ADD_553_U70 & P3_U4298); 
assign P3_U5737 = ~(P3_ADD_515_U67 & P3_U4302); 
assign P3_U5741 = ~(P3_ADD_405_U68 & P3_U4305); 
assign P3_U5743 = ~(P3_ADD_385_U70 & P3_U2358); 
assign P3_U5745 = ~(P3_ADD_349_U70 & P3_U4306); 
assign P3_U5746 = ~(P3_ADD_344_U70 & P3_U2362); 
assign P3_U5755 = ~(P3_ADD_553_U69 & P3_U4298); 
assign P3_U5761 = ~(P3_ADD_515_U66 & P3_U4302); 
assign P3_U5765 = ~(P3_ADD_405_U67 & P3_U4305); 
assign P3_U5767 = ~(P3_ADD_385_U69 & P3_U2358); 
assign P3_U5769 = ~(P3_ADD_349_U69 & P3_U4306); 
assign P3_U5770 = ~(P3_ADD_344_U69 & P3_U2362); 
assign P3_U5779 = ~(P3_ADD_553_U68 & P3_U4298); 
assign P3_U5785 = ~(P3_ADD_515_U65 & P3_U4302); 
assign P3_U5789 = ~(P3_ADD_405_U66 & P3_U4305); 
assign P3_U5791 = ~(P3_ADD_385_U68 & P3_U2358); 
assign P3_U5793 = ~(P3_ADD_349_U68 & P3_U4306); 
assign P3_U5794 = ~(P3_ADD_344_U68 & P3_U2362); 
assign P3_U5803 = ~(P3_ADD_553_U67 & P3_U4298); 
assign P3_U5807 = ~(P3_ADD_531_U67 & P3_U2354); 
assign P3_U5809 = ~(P3_ADD_515_U64 & P3_U4302); 
assign P3_U5813 = ~(P3_ADD_405_U65 & P3_U4305); 
assign P3_U5815 = ~(P3_ADD_385_U67 & P3_U2358); 
assign P3_U5816 = ~(P3_ADD_380_U67 & P3_U2359); 
assign P3_U5817 = ~(P3_ADD_349_U67 & P3_U4306); 
assign P3_U5818 = ~(P3_ADD_344_U67 & P3_U2362); 
assign P3_U5833 = ~(P3_ADD_515_U63 & P3_U4302); 
assign P3_U5834 = ~(P3_ADD_494_U63 & P3_U2356); 
assign P3_U5835 = ~(P3_ADD_476_U63 & P3_U4303); 
assign P3_U5836 = ~(P3_ADD_441_U63 & P3_U4304); 
assign P3_U5837 = ~(P3_ADD_405_U64 & P3_U4305); 
assign P3_U5838 = ~(P3_ADD_394_U64 & P3_U2357); 
assign P3_U5928 = ~(P3_ADD_526_U79 & P3_U2355); 
assign P3_U5952 = ~(P3_ADD_526_U78 & P3_U2355); 
assign P3_U7378 = ~(P3_U7377 & P3_STATE2_REG_0__SCAN_IN); 
assign P2_U2703 = ~(P2_U7727 & P2_U7726); 
assign P2_U2716 = ~(P2_U7620 & P2_U7619 & P2_U7618 & P2_U7617); 
assign P2_U2717 = ~(P2_U7624 & P2_U7623 & P2_U7622 & P2_U7621); 
assign P2_U2718 = ~(P2_U7632 & P2_U7631 & P2_U7630 & P2_U7629); 
assign P2_U2719 = ~(P2_U7636 & P2_U7635 & P2_U7634 & P2_U7633); 
assign P2_U2720 = ~(P2_U7640 & P2_U7639 & P2_U7638 & P2_U7637); 
assign P2_U2721 = ~(P2_U7644 & P2_U7643 & P2_U7642 & P2_U7641); 
assign P2_U2722 = ~(P2_U7648 & P2_U7647 & P2_U7646 & P2_U7645); 
assign P2_U2723 = ~(P2_U7652 & P2_U7651 & P2_U7650 & P2_U7649); 
assign P2_U2724 = ~(P2_U7656 & P2_U7655 & P2_U7654 & P2_U7653); 
assign P2_U2725 = ~(P2_U7660 & P2_U7659 & P2_U7658 & P2_U7657); 
assign P2_U2726 = ~(P2_U7664 & P2_U7663 & P2_U7662 & P2_U7661); 
assign P2_U2727 = ~(P2_U7668 & P2_U7667 & P2_U7666 & P2_U7665); 
assign P2_U2728 = ~(P2_U7676 & P2_U7675 & P2_U7674 & P2_U7673); 
assign P2_U2729 = ~(P2_U7680 & P2_U7679 & P2_U7678 & P2_U7677); 
assign P2_U2730 = ~(P2_U7684 & P2_U7683 & P2_U7682 & P2_U7681); 
assign P2_U2731 = ~(P2_U7688 & P2_U7687 & P2_U7686 & P2_U7685); 
assign P2_U2732 = ~(P2_U7692 & P2_U7691 & P2_U7690 & P2_U7689); 
assign P2_U2733 = ~(P2_U7696 & P2_U7695 & P2_U7694 & P2_U7693); 
assign P2_U2734 = ~(P2_U7700 & P2_U7699 & P2_U7698 & P2_U7697); 
assign P2_U2735 = ~(P2_U7704 & P2_U7703 & P2_U7702 & P2_U7701); 
assign P2_U2736 = ~(P2_U7708 & P2_U7707 & P2_U7706 & P2_U7705); 
assign P2_U2737 = ~(P2_U7712 & P2_U7711 & P2_U7710 & P2_U7709); 
assign P2_U2738 = ~(P2_U7596 & P2_U7595 & P2_U7594 & P2_U7593); 
assign P2_U2739 = ~(P2_U7600 & P2_U7599 & P2_U7598 & P2_U7597); 
assign P2_U2740 = ~(P2_U7604 & P2_U7603 & P2_U7602 & P2_U7601); 
assign P2_U2741 = ~(P2_U7608 & P2_U7607 & P2_U7606 & P2_U7605); 
assign P2_U2742 = ~(P2_U7612 & P2_U7611 & P2_U7610 & P2_U7609); 
assign P2_U2743 = ~(P2_U7616 & P2_U7615 & P2_U7614 & P2_U7613); 
assign P2_U2744 = ~(P2_U7628 & P2_U7627 & P2_U7626 & P2_U7625); 
assign P2_U2745 = ~(P2_U7672 & P2_U7671 & P2_U7670 & P2_U7669); 
assign P2_U2746 = ~(P2_U7716 & P2_U7715 & P2_U7714 & P2_U7713); 
assign P2_U3648 = ~(P2_U8352 & P2_U8351); 
assign P2_U3649 = ~(P2_U8354 & P2_U8353); 
assign P2_U3684 = ~(P2_U8424 & P2_U8423); 
assign P2_U3685 = ~(P2_U8426 & P2_U8425); 
assign P2_U3715 = P2_U3714 & P2_U4618; 
assign P2_U3884 = P2_U3883 & P2_U5609; 
assign P2_U3885 = P2_U4396 & P2_U5617; 
assign P2_U3888 = P2_U5627 & P2_U5626; 
assign P2_U3890 = P2_U5635 & P2_U5634; 
assign P2_U4389 = P2_U7719 & P2_U7718; 
assign P2_U5603 = ~(P2_U2514 & P2_U3288); 
assign P2_U5675 = ~(P2_U3895 & P2_U2514); 
assign P2_U7141 = ~(P2_ADD_402_1132_U23 & P2_U2355); 
assign P2_U7722 = ~(P2_U7720 & P2_U3575); 
assign P2_U7888 = ~(P2_U4386 & P2_U7887 & P2_U2589 & P2_U4385 & P2_U4384); 
assign P2_U7890 = ~(P2_U7889 & P2_U4458 & P2_U2589 & P2_U4379); 
assign P2_U8361 = ~(P2_R2337_U61 & P2_U3284); 
assign P1_U2615 = ~(P1_U6753 & P1_U4004); 
assign P1_U2711 = ~(P1_U7377 & P1_U7376); 
assign P1_U2716 = ~(P1_U7365 & P1_U7364); 
assign P1_U2717 = ~(P1_U7367 & P1_U7366); 
assign P1_U2723 = P1_U7236 & P1_U7083; 
assign P1_U2724 = P1_U7253 & P1_U7083; 
assign P1_U2725 = P1_U7270 & P1_U7083; 
assign P1_U2726 = P1_U7620 & P1_U7083; 
assign P1_U2727 = P1_U7302 & P1_U7083; 
assign P1_U2728 = P1_U7319 & P1_U7083; 
assign P1_U2729 = P1_U7336 & P1_U7083; 
assign P1_U2730 = P1_U7353 & P1_U7083; 
assign P1_U2732 = P1_U7083 & P1_U7082; 
assign P1_U2733 = P1_U7114 & P1_U7083; 
assign P1_U2734 = P1_U7131 & P1_U7083; 
assign P1_U2735 = P1_U7618 & P1_U7083; 
assign P1_U2736 = P1_U7163 & P1_U7083; 
assign P1_U2737 = P1_U7180 & P1_U7083; 
assign P1_U2738 = P1_U7197 & P1_U7083; 
assign P1_U2739 = P1_U7214 & P1_U7083; 
assign P1_U2761 = ~(P1_U6928 & P1_U6927); 
assign P1_U2762 = ~(P1_U6930 & P1_U6929); 
assign P1_U2763 = ~(P1_U6932 & P1_U6931); 
assign P1_U2764 = ~(P1_U6934 & P1_U6933); 
assign P1_U3450 = ~(P1_U4074 & P1_U7093 & P1_U4075 & P1_U4077); 
assign P1_U4114 = P1_U7090 & P1_U3434 & P1_U4111 & P1_U4113; 
assign P1_U4116 = P1_U7505 & P1_U7489 & P1_U7488 & P1_U7487; 
assign P1_U4156 = P1_U4155 & P1_U7359; 
assign P1_U5499 = ~(P1_U4494 & P1_U7707); 
assign P1_U6752 = ~(P1_R2337_U63 & P1_U2352); 
assign P1_U7479 = ~(P1_U4117 & P1_U7093 & P1_U4118 & P1_U4120); 
assign P1_U7792 = ~(P1_U7707 & P1_U4494); 
assign P3_ADD_526_U31 = ~(P3_ADD_526_U88 & P3_ADD_526_U124); 
assign P3_ADD_526_U107 = ~(P3_ADD_526_U124 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_526_U191 = ~(P3_ADD_526_U124 & P3_ADD_526_U26); 
assign P3_ADD_526_U194 = ~(P3_ADD_526_U138 & P3_ADD_526_U23); 
assign P3_ADD_552_U31 = ~(P3_ADD_552_U88 & P3_ADD_552_U124); 
assign P3_ADD_552_U107 = ~(P3_ADD_552_U124 & P3_EBX_REG_15__SCAN_IN); 
assign P3_ADD_552_U191 = ~(P3_ADD_552_U124 & P3_ADD_552_U26); 
assign P3_ADD_552_U194 = ~(P3_ADD_552_U138 & P3_ADD_552_U23); 
assign P3_ADD_546_U31 = ~(P3_ADD_546_U88 & P3_ADD_546_U124); 
assign P3_ADD_546_U107 = ~(P3_ADD_546_U124 & P3_EAX_REG_15__SCAN_IN); 
assign P3_ADD_546_U191 = ~(P3_ADD_546_U124 & P3_ADD_546_U26); 
assign P3_ADD_546_U194 = ~(P3_ADD_546_U138 & P3_ADD_546_U23); 
assign P3_GTE_401_U6 = ~(P3_SUB_401_U6 | P3_GTE_401_U8); 
assign P3_ADD_391_1180_U24 = ~(P3_ADD_391_1180_U48 & P3_ADD_391_1180_U47); 
assign P3_ADD_391_1180_U29 = ~P3_ADD_391_1180_U8; 
assign P3_ADD_391_1180_U45 = ~(P3_U2615 & P3_ADD_391_1180_U8); 
assign P3_ADD_476_U20 = ~(P3_ADD_476_U100 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_476_U124 = ~(P3_ADD_476_U100 & P3_ADD_476_U18); 
assign P3_GTE_390_U6 = ~(P3_SUB_390_U6 | P3_GTE_390_U8); 
assign P3_ADD_531_U22 = ~(P3_ADD_531_U104 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_531_U131 = ~(P3_ADD_531_U104 & P3_ADD_531_U20); 
assign P3_SUB_320_U25 = ~P3_ADD_318_U63; 
assign P3_SUB_320_U55 = P3_SUB_320_U131 & P3_SUB_320_U130; 
assign P3_SUB_320_U88 = ~(P3_ADD_318_U63 & P3_SUB_320_U87); 
assign P3_GTE_485_U6 = ~(P3_SUB_485_U6 | P3_GTE_485_U7); 
assign P3_ADD_318_U20 = ~(P3_ADD_318_U100 & P3_PHYADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_318_U124 = ~(P3_ADD_318_U100 & P3_ADD_318_U18); 
assign P3_ADD_315_U20 = ~(P3_ADD_315_U97 & P3_PHYADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_315_U176 = ~(P3_ADD_315_U97 & P3_ADD_315_U19); 
assign P3_GTE_355_U6 = ~(P3_SUB_355_U6 | P3_GTE_355_U8); 
assign P3_ADD_360_1242_U29 = ~P3_ADD_360_U21; 
assign P3_ADD_360_1242_U122 = ~P3_ADD_360_1242_U75; 
assign P3_ADD_360_1242_U127 = ~(P3_ADD_360_1242_U126 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_360_1242_U129 = P3_ADD_360_U21 | P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_360_1242_U131 = ~(P3_ADD_360_U21 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_360_1242_U232 = ~(P3_ADD_360_U21 & P3_ADD_360_1242_U30); 
assign P3_ADD_360_1242_U234 = ~(P3_ADD_360_U21 & P3_ADD_360_1242_U30); 
assign P3_ADD_360_1242_U246 = ~(P3_ADD_360_1242_U245 & P3_ADD_360_1242_U244); 
assign P3_ADD_467_U20 = ~(P3_ADD_467_U100 & P3_REIP_REG_9__SCAN_IN); 
assign P3_ADD_467_U124 = ~(P3_ADD_467_U100 & P3_ADD_467_U18); 
assign P3_ADD_430_U20 = ~(P3_ADD_430_U100 & P3_REIP_REG_9__SCAN_IN); 
assign P3_ADD_430_U124 = ~(P3_ADD_430_U100 & P3_ADD_430_U18); 
assign P3_ADD_380_U22 = ~(P3_ADD_380_U104 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_380_U131 = ~(P3_ADD_380_U104 & P3_ADD_380_U20); 
assign P3_GTE_370_U6 = ~(P3_SUB_370_U6 | P3_GTE_370_U8); 
assign P3_ADD_344_U22 = ~(P3_ADD_344_U104 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_344_U131 = ~(P3_ADD_344_U104 & P3_ADD_344_U20); 
assign P3_ADD_339_U20 = ~(P3_ADD_339_U100 & P3_PHYADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_339_U124 = ~(P3_ADD_339_U100 & P3_ADD_339_U18); 
assign P3_ADD_360_U20 = ~(P3_ADD_360_U38 & P3_ADD_360_U37); 
assign P3_ADD_360_U25 = ~P3_ADD_360_U9; 
assign P3_ADD_360_U35 = ~(P3_U2625 & P3_ADD_360_U9); 
assign P3_ADD_541_U20 = ~(P3_ADD_541_U100 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_541_U124 = ~(P3_ADD_541_U100 & P3_ADD_541_U18); 
assign P3_SUB_357_1258_U161 = ~P3_SUB_357_1258_U30; 
assign P3_SUB_357_1258_U422 = ~(P3_SUB_357_1258_U30 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_SUB_357_1258_U425 = ~(P3_SUB_357_1258_U30 & P3_SUB_357_1258_U34 & P3_SUB_357_U7); 
assign P3_SUB_357_1258_U483 = ~(P3_SUB_357_1258_U28 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_ADD_515_U20 = ~(P3_ADD_515_U100 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_515_U124 = ~(P3_ADD_515_U100 & P3_ADD_515_U18); 
assign P3_ADD_394_U20 = ~(P3_ADD_394_U103 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_394_U128 = ~(P3_ADD_394_U103 & P3_ADD_394_U18); 
assign P3_GTE_450_U6 = ~(P3_SUB_450_U6 | P3_GTE_450_U7); 
assign P3_SUB_414_U8 = P3_SUB_414_U122 & P3_SUB_414_U30; 
assign P3_SUB_414_U31 = ~(P3_SUB_414_U46 & P3_SUB_414_U77 & P3_SUB_414_U95); 
assign P3_SUB_414_U119 = ~(P3_SUB_414_U95 & P3_SUB_414_U77); 
assign P3_SUB_414_U155 = ~(P3_SUB_414_U95 & P3_SUB_414_U77); 
assign P3_ADD_441_U20 = ~(P3_ADD_441_U100 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_441_U124 = ~(P3_ADD_441_U100 & P3_ADD_441_U18); 
assign P3_ADD_349_U22 = ~(P3_ADD_349_U104 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_349_U131 = ~(P3_ADD_349_U104 & P3_ADD_349_U20); 
assign P3_ADD_405_U20 = ~(P3_ADD_405_U103 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_405_U128 = ~(P3_ADD_405_U103 & P3_ADD_405_U18); 
assign P3_ADD_553_U22 = ~(P3_ADD_553_U104 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_553_U131 = ~(P3_ADD_553_U104 & P3_ADD_553_U20); 
assign P3_ADD_558_U22 = ~(P3_ADD_558_U104 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_558_U131 = ~(P3_ADD_558_U104 & P3_ADD_558_U20); 
assign P3_ADD_385_U22 = ~(P3_ADD_385_U104 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_385_U131 = ~(P3_ADD_385_U104 & P3_ADD_385_U20); 
assign P3_ADD_357_U7 = P3_ADD_357_U29 & P3_ADD_357_U11; 
assign P3_ADD_357_U12 = ~(P3_ADD_357_U14 & P3_ADD_357_U22); 
assign P3_ADD_357_U13 = ~(P3_ADD_357_U35 & P3_ADD_357_U34); 
assign P3_ADD_357_U26 = ~(P3_ADD_357_U22 & P3_ADD_357_U18); 
assign P3_ADD_357_U33 = ~(P3_ADD_357_U22 & P3_ADD_357_U18); 
assign P3_ADD_547_U22 = ~(P3_ADD_547_U104 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_547_U131 = ~(P3_ADD_547_U104 & P3_ADD_547_U20); 
assign P3_ADD_371_1212_U26 = ~P3_ADD_371_U5; 
assign P3_ADD_371_1212_U29 = ~(P3_ADD_371_U5 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_371_1212_U35 = ~P3_ADD_371_U21; 
assign P3_ADD_371_1212_U77 = ~(P3_ADD_371_U21 & P3_ADD_371_1212_U121); 
assign P3_ADD_371_1212_U87 = ~(P3_ADD_371_1212_U265 & P3_ADD_371_1212_U264); 
assign P3_ADD_371_1212_U125 = P3_ADD_371_U5 | P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_371_1212_U157 = P3_ADD_371_U5 | P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_371_1212_U175 = P3_ADD_371_U5 | P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_ADD_371_1212_U241 = ~(P3_ADD_371_U5 & P3_ADD_371_1212_U27); 
assign P3_ADD_371_1212_U252 = ~(P3_ADD_371_1212_U121 & P3_ADD_371_1212_U33); 
assign P3_ADD_371_1212_U254 = ~(P3_ADD_371_1212_U34 & P3_ADD_371_1212_U33 & P3_ADD_371_U21); 
assign P3_ADD_371_U28 = ~P3_ADD_371_U9; 
assign P3_ADD_371_U39 = ~(P3_U2625 & P3_ADD_371_U9); 
assign P3_ADD_371_U42 = ~(P3_ADD_371_U27 & P3_ADD_371_U8); 
assign P3_GTE_412_U6 = ~(P3_SUB_412_U6 | P3_GTE_412_U7); 
assign P3_GTE_504_U6 = ~(P3_SUB_504_U6 | P3_GTE_504_U7); 
assign P3_ADD_494_U20 = ~(P3_ADD_494_U100 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_494_U124 = ~(P3_ADD_494_U100 & P3_ADD_494_U18); 
assign P3_ADD_536_U20 = ~(P3_ADD_536_U100 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_536_U124 = ~(P3_ADD_536_U100 & P3_ADD_536_U18); 
assign P3_ADD_402_1132_U24 = ~(P3_ADD_402_1132_U48 & P3_ADD_402_1132_U47); 
assign P3_ADD_402_1132_U29 = ~P3_ADD_402_1132_U8; 
assign P3_ADD_402_1132_U45 = ~(P3_U2615 & P3_ADD_402_1132_U8); 
assign P2_ADD_402_1132_U20 = ~(P2_ADD_402_1132_U40 & P2_ADD_402_1132_U39); 
assign P2_ADD_402_1132_U29 = ~P2_ADD_402_1132_U8; 
assign P2_ADD_402_1132_U49 = ~(P2_U2593 & P2_ADD_402_1132_U8); 
assign P2_R2182_U103 = P2_R2182_U204 & P2_R2182_U203; 
assign P2_R2182_U207 = ~(P2_R2182_U206 & P2_R2182_U205); 
assign P2_R2167_U15 = ~P2_U2361; 
assign P2_R2027_U22 = ~(P2_R2027_U104 & P2_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P2_R2027_U131 = ~(P2_R2027_U104 & P2_R2027_U20); 
assign P2_R2337_U21 = ~(P2_R2337_U101 & P2_PHYADDRPOINTER_REG_10__SCAN_IN); 
assign P2_R2337_U182 = ~(P2_R2337_U101 & P2_R2337_U20); 
assign P2_R2219_U45 = ~(P2_U2765 & P2_R2219_U23); 
assign P2_R2219_U47 = ~(P2_U2764 & P2_R2219_U14); 
assign P2_R2219_U48 = ~(P2_U2763 & P2_R2219_U17); 
assign P2_R2219_U50 = ~(P2_U2755 & P2_R2219_U12); 
assign P2_R2219_U52 = ~(P2_U2762 & P2_R2219_U18); 
assign P2_R2219_U53 = ~(P2_U2754 & P2_R2219_U13); 
assign P2_R2219_U55 = ~(P2_U2761 & P2_R2219_U10); 
assign P2_R2219_U56 = ~(P2_U2753 & P2_R2219_U11); 
assign P2_R2219_U69 = ~(P2_U2757 & P2_R2219_U15); 
assign P2_R2219_U70 = ~(P2_U2756 & P2_R2219_U16); 
assign P2_R2219_U76 = ~(P2_U2762 & P2_R2219_U18); 
assign P2_R2219_U77 = ~(P2_U2764 & P2_R2219_U14); 
assign P2_R2219_U84 = ~P2_R2219_U32; 
assign P2_R2219_U89 = ~P2_R2219_U33; 
assign P2_R2219_U94 = ~P2_R2219_U34; 
assign P2_R2219_U97 = ~(P2_U2761 & P2_R2219_U10); 
assign P2_R2219_U98 = ~(P2_U2753 & P2_R2219_U11); 
assign P2_R2219_U102 = ~(P2_U2762 & P2_R2219_U18); 
assign P2_R2219_U103 = ~(P2_U2754 & P2_R2219_U13); 
assign P2_R2219_U107 = ~(P2_U2763 & P2_R2219_U17); 
assign P2_R2219_U108 = ~(P2_U2755 & P2_R2219_U12); 
assign P2_R2219_U112 = ~(P2_U2764 & P2_R2219_U14); 
assign P2_R2219_U113 = ~(P2_U2756 & P2_R2219_U16); 
assign P2_R2096_U115 = ~P2_R2096_U113; 
assign P2_R2096_U117 = ~(P2_R2096_U55 & P2_R2096_U116); 
assign P2_R2096_U169 = ~P2_R2096_U112; 
assign P2_R2096_U176 = ~(P2_U2650 & P2_R2096_U67); 
assign P2_R2096_U178 = ~(P2_U2650 & P2_R2096_U67); 
assign P2_R2096_U183 = ~(P2_U2651 & P2_R2096_U65); 
assign P2_R2096_U185 = ~(P2_U2651 & P2_R2096_U65); 
assign P2_R2096_U190 = ~(P2_U2652 & P2_R2096_U63); 
assign P2_R2096_U192 = ~(P2_U2652 & P2_R2096_U63); 
assign P2_R2096_U197 = ~(P2_U2653 & P2_R2096_U61); 
assign P2_R2096_U199 = ~(P2_U2653 & P2_R2096_U61); 
assign P2_R2096_U204 = ~(P2_U2654 & P2_R2096_U59); 
assign P2_R2096_U206 = ~(P2_U2654 & P2_R2096_U59); 
assign P2_R2096_U213 = ~(P2_U2655 & P2_R2096_U57); 
assign P2_R2096_U215 = ~(P2_U2655 & P2_R2096_U57); 
assign P2_R2096_U239 = ~(P2_U2648 & P2_R2096_U112); 
assign P2_R2096_U242 = ~(P2_U2656 & P2_R2096_U116 & P2_R2096_U54); 
assign P2_R2096_U265 = ~(P2_U2657 & P2_R2096_U53); 
assign P2_R1957_U25 = ~P2_U3654; 
assign P2_R1957_U55 = P2_R1957_U131 & P2_R1957_U130; 
assign P2_R1957_U88 = ~(P2_U3654 & P2_R1957_U87); 
assign P2_ADD_394_U20 = ~(P2_ADD_394_U103 & P2_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P2_ADD_394_U142 = ~(P2_ADD_394_U103 & P2_ADD_394_U19); 
assign P1_R2027_U31 = ~(P1_R2027_U88 & P1_R2027_U124); 
assign P1_R2027_U107 = ~(P1_R2027_U124 & P1_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P1_R2027_U191 = ~(P1_R2027_U124 & P1_R2027_U26); 
assign P1_R2027_U194 = ~(P1_R2027_U138 & P1_R2027_U23); 
assign P1_R2144_U14 = ~P1_U2751; 
assign P1_R2144_U27 = ~(P1_R2144_U206 & P1_R2144_U205); 
assign P1_R2144_U29 = ~(P1_R2144_U203 & P1_R2144_U202); 
assign P1_R2144_U31 = ~(P1_R2144_U224 & P1_R2144_U223); 
assign P1_R2144_U32 = ~(P1_R2144_U221 & P1_R2144_U220); 
assign P1_R2144_U33 = ~(P1_R2144_U227 & P1_R2144_U226); 
assign P1_R2144_U34 = ~(P1_R2144_U230 & P1_R2144_U229); 
assign P1_R2144_U35 = ~(P1_R2144_U233 & P1_R2144_U232); 
assign P1_R2144_U36 = ~(P1_R2144_U236 & P1_R2144_U235); 
assign P1_R2358_U406 = ~(P1_U2352 & P1_R2358_U145); 
assign P1_R2358_U417 = ~(P1_U2352 & P1_R2358_U145); 
assign P1_R2099_U88 = P1_R2099_U34 & P1_R2099_U35; 
assign P1_R2099_U89 = P1_R2099_U31 & P1_R2099_U30; 
assign P1_R2099_U90 = P1_R2099_U29 & P1_R2099_U28; 
assign P1_R2099_U91 = P1_R2099_U26 & P1_R2099_U27; 
assign P1_R2099_U92 = P1_R2099_U63 & P1_R2099_U62; 
assign P1_R2099_U93 = P1_R2099_U61 & P1_R2099_U60; 
assign P1_R2099_U94 = P1_R2099_U59 & P1_R2099_U58; 
assign P1_R2099_U95 = P1_R2099_U57 & P1_R2099_U56; 
assign P1_R2099_U96 = P1_R2099_U44 & P1_R2099_U43; 
assign P1_R2099_U147 = ~(P1_R2099_U32 & P1_R2099_U146); 
assign P1_R2099_U152 = ~(P1_U2678 & P1_R2099_U33); 
assign P1_R2099_U184 = ~P1_R2099_U27; 
assign P1_R2099_U187 = ~P1_R2099_U32; 
assign P1_R2099_U190 = ~P1_R2099_U33; 
assign P1_R2099_U193 = ~P1_R2099_U35; 
assign P1_R2099_U196 = ~P1_R2099_U34; 
assign P1_R2099_U199 = ~P1_R2099_U30; 
assign P1_R2099_U202 = ~P1_R2099_U31; 
assign P1_R2099_U205 = ~P1_R2099_U28; 
assign P1_R2099_U208 = ~P1_R2099_U29; 
assign P1_R2099_U211 = ~P1_R2099_U26; 
assign P1_R2099_U228 = ~P1_R2099_U45; 
assign P1_R2099_U231 = ~P1_R2099_U46; 
assign P1_R2099_U234 = ~P1_R2099_U47; 
assign P1_R2099_U237 = ~P1_R2099_U48; 
assign P1_R2099_U240 = ~P1_R2099_U49; 
assign P1_R2099_U243 = ~P1_R2099_U50; 
assign P1_R2099_U246 = ~P1_R2099_U51; 
assign P1_R2099_U249 = ~P1_R2099_U52; 
assign P1_R2099_U252 = ~P1_R2099_U53; 
assign P1_R2099_U255 = ~P1_R2099_U54; 
assign P1_R2099_U258 = ~P1_R2099_U55; 
assign P1_R2099_U261 = ~P1_R2099_U62; 
assign P1_R2099_U264 = ~P1_R2099_U63; 
assign P1_R2099_U267 = ~P1_R2099_U60; 
assign P1_R2099_U270 = ~P1_R2099_U61; 
assign P1_R2099_U273 = ~P1_R2099_U58; 
assign P1_R2099_U276 = ~P1_R2099_U59; 
assign P1_R2099_U279 = ~P1_R2099_U56; 
assign P1_R2099_U282 = ~P1_R2099_U57; 
assign P1_R2099_U285 = ~P1_R2099_U43; 
assign P1_R2099_U288 = ~P1_R2099_U44; 
assign P1_R2099_U291 = ~P1_R2099_U97; 
assign P1_R2099_U319 = ~(P1_R2099_U33 & P1_R2099_U6); 
assign P1_R2099_U321 = ~(P1_R2099_U33 & P1_R2099_U6); 
assign P1_R2099_U348 = ~(P1_R2099_U32 & P1_R2099_U347); 
assign P1_R2167_U12 = ~P1_U2718; 
assign P1_R2167_U15 = ~P1_U2356; 
assign P1_R2167_U25 = ~(P1_U2715 & P1_R2167_U22); 
assign P1_R2167_U27 = ~(P1_U2714 & P1_R2167_U8); 
assign P1_R2167_U30 = ~(P1_U2719 & P1_R2167_U10); 
assign P1_R2167_U32 = ~(P1_U2713 & P1_R2167_U9); 
assign P1_R2167_U35 = ~(P1_U2718 & P1_R2167_U11); 
assign P1_R2337_U20 = ~(P1_R2337_U100 & P1_PHYADDRPOINTER_REG_9__SCAN_IN); 
assign P1_R2337_U124 = ~(P1_R2337_U100 & P1_R2337_U18); 
assign P1_R2096_U20 = ~(P1_R2096_U100 & P1_REIP_REG_9__SCAN_IN); 
assign P1_R2096_U124 = ~(P1_R2096_U100 & P1_R2096_U18); 
assign P1_ADD_371_U11 = ~(P1_U3231 & P1_ADD_371_U28); 
assign P1_ADD_371_U24 = P1_ADD_371_U40 & P1_ADD_371_U39; 
assign P1_ADD_371_U36 = ~(P1_ADD_371_U28 & P1_ADD_371_U10); 
assign P1_ADD_405_U20 = ~(P1_ADD_405_U103 & P1_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P1_ADD_405_U142 = ~(P1_ADD_405_U103 & P1_ADD_405_U19); 
assign P1_GTE_485_U6 = ~(P1_R2238_U6 | P1_GTE_485_U7); 
assign P1_ADD_515_U20 = ~(P1_ADD_515_U100 & P1_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P1_ADD_515_U140 = ~(P1_ADD_515_U100 & P1_ADD_515_U19); 
assign P3_U2504 = P3_U4660 & P3_U3271; 
assign P3_U2508 = P3_U4660 & P3_U7968; 
assign P3_U2867 = P3_U5579 & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign P3_U3144 = ~(P3_U4647 & P3_U2486); 
assign P3_U3149 = ~(P3_U2490 & P3_U2486); 
assign P3_U3157 = ~(P3_U2493 & P3_U2486); 
assign P3_U3162 = ~(P3_U2495 & P3_U2486); 
assign P3_U3166 = ~(P3_U2498 & P3_U4647); 
assign P3_U3170 = ~(P3_U2498 & P3_U2490); 
assign P3_U3174 = ~(P3_U2498 & P3_U2493); 
assign P3_U3178 = ~(P3_U2498 & P3_U2495); 
assign P3_U3210 = ~P3_GTE_412_U6; 
assign P3_U3211 = ~P3_GTE_485_U6; 
assign P3_U3212 = ~P3_GTE_390_U6; 
assign P3_U3213 = ~P3_GTE_450_U6; 
assign P3_U3214 = ~P3_GTE_504_U6; 
assign P3_U3215 = ~P3_GTE_401_U6; 
assign P3_U3221 = ~(P3_U3222 & P3_U3119 & P3_U5524); 
assign P3_U3237 = ~P3_GTE_370_U6; 
assign P3_U3238 = ~P3_GTE_355_U6; 
assign P3_U3511 = P3_U5087 & P3_U5086; 
assign P3_U3513 = P3_U5092 & P3_U5091; 
assign P3_U3515 = P3_U5097 & P3_U5096; 
assign P3_U3517 = P3_U5102 & P3_U5101; 
assign P3_U3519 = P3_U5107 & P3_U5106; 
assign P3_U3521 = P3_U5112 & P3_U5111; 
assign P3_U3523 = P3_U5117 & P3_U5116; 
assign P3_U3525 = P3_U5122 & P3_U5121; 
assign P3_U3694 = P3_U3695 & P3_U5641; 
assign P3_U3696 = P3_U5643 & P3_U5642 & P3_U5644 & P3_U5646 & P3_U5645; 
assign P3_U3701 = P3_U3702 & P3_U5665; 
assign P3_U3703 = P3_U5667 & P3_U5666 & P3_U5668 & P3_U5670 & P3_U5669; 
assign P3_U3704 = P3_U5674 & P3_U5671 & P3_U5672 & P3_U5673; 
assign P3_U3708 = P3_U3709 & P3_U5689; 
assign P3_U3711 = P3_U5691 & P3_U5690 & P3_U5692 & P3_U5694 & P3_U5693; 
assign P3_U3712 = P3_U5698 & P3_U5695 & P3_U5696 & P3_U5697; 
assign P3_U3716 = P3_U3717 & P3_U5713; 
assign P3_U3719 = P3_U5715 & P3_U5714 & P3_U5716 & P3_U5718 & P3_U5717; 
assign P3_U3720 = P3_U5722 & P3_U5719 & P3_U5720 & P3_U5721; 
assign P3_U3724 = P3_U3725 & P3_U5737; 
assign P3_U3727 = P3_U5739 & P3_U5738 & P3_U5740 & P3_U5742 & P3_U5741; 
assign P3_U3728 = P3_U5746 & P3_U5743 & P3_U5744 & P3_U5745; 
assign P3_U3732 = P3_U3733 & P3_U5761; 
assign P3_U3735 = P3_U5763 & P3_U5762 & P3_U5764 & P3_U5766 & P3_U5765; 
assign P3_U3736 = P3_U5770 & P3_U5767 & P3_U5768 & P3_U5769; 
assign P3_U3740 = P3_U3741 & P3_U5785; 
assign P3_U3743 = P3_U5787 & P3_U5786 & P3_U5788 & P3_U5790 & P3_U5789; 
assign P3_U3744 = P3_U5794 & P3_U5791 & P3_U5792 & P3_U5793; 
assign P3_U3749 = P3_U5807 & P3_U5808; 
assign P3_U3751 = P3_U5811 & P3_U5810 & P3_U5812 & P3_U5814 & P3_U5813; 
assign P3_U3752 = P3_U5818 & P3_U5815 & P3_U5816 & P3_U5817; 
assign P3_U3758 = P3_U5835 & P3_U5834 & P3_U5836 & P3_U5838 & P3_U5837; 
assign P3_U4299 = ~P3_U3243; 
assign P3_U4352 = ~P3_U3222; 
assign P3_U5486 = ~(P3_GTE_450_U6 & P3_U4303); 
assign P3_U5487 = ~(P3_GTE_504_U6 & P3_U4302); 
assign P3_U5489 = ~(P3_GTE_412_U6 & P3_U4304); 
assign P3_U5490 = ~(P3_GTE_485_U6 & P3_U2356); 
assign P3_U5493 = ~(P3_GTE_390_U6 & P3_U2357); 
assign P3_U5495 = ~(P3_GTE_401_U6 & P3_U4305); 
assign P3_U5512 = ~(P3_U5509 & P3_U3665); 
assign P3_U5534 = ~P3_U3226; 
assign P3_U5540 = ~(P3_U5506 & P3_U3226); 
assign P3_U5560 = ~P3_U3231; 
assign P3_U5564 = ~(P3_U5558 & P3_U3231); 
assign P3_U5591 = ~(P3_U5581 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_U5598 = ~(P3_U5597 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_U5599 = ~(P3_U5595 & P3_U3233); 
assign P3_U5609 = ~(P3_U5608 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_U5615 = ~(P3_U5614 & P3_U3233); 
assign P3_U5616 = ~(P3_U5612 & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P3_U5617 = ~(P3_U2463 & P3_U4294 & P3_GTE_450_U6); 
assign P3_U5618 = ~(P3_GTE_370_U6 & P3_U4344); 
assign P3_U5620 = ~(P3_U4590 & P3_U2630 & P3_GTE_412_U6); 
assign P3_U5621 = ~(P3_GTE_355_U6 & P3_U3074); 
assign P3_U5623 = ~(P3_GTE_390_U6 & P3_U4488); 
assign P3_U5625 = ~(P3_U3102 & P3_U3108 & P3_GTE_401_U6); 
assign P3_U5626 = ~(P3_U4349 & P3_GTE_504_U6); 
assign P3_U5627 = ~(P3_U4348 & P3_GTE_485_U6); 
assign P3_U5651 = ~(P3_ADD_371_1212_U87 & P3_U2360); 
assign P3_U6399 = ~(P3_GTE_355_U6 & P3_U2361); 
assign P3_U6400 = ~(P3_GTE_370_U6 & P3_U2360); 
assign P3_U6661 = ~(P3_U4304 & P3_U2630 & P3_GTE_412_U6); 
assign P3_U6662 = ~(P3_GTE_450_U6 & P3_U4303); 
assign P3_U6996 = ~(P3_GTE_401_U6 & P3_U4305); 
assign P3_U7379 = ~(P3_U3125 & P3_U7378); 
assign P2_U2688 = P2_ADD_402_1132_U20 & P2_U2355; 
assign P2_U2689 = ~(P2_U7142 & P2_U7141); 
assign P2_U2751 = P2_U7888 & P2_U7737; 
assign P2_U3653 = ~(P2_U8362 & P2_U8361); 
assign P2_U7583 = ~(P2_U7890 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U7584 = ~(P2_U7890 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P2_U7588 = ~(P2_U7890 & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P2_U7886 = ~(P2_U7722 & P2_U5589); 
assign P1_U2519 = P1_U3744 & P1_U5499; 
assign P1_U2744 = P1_U7479 & P1_U7478; 
assign P1_U3246 = ~(P1_U7792 & P1_U7791 & P1_U4158 & P1_U4156); 
assign P1_U3388 = ~P1_GTE_485_U6; 
assign P1_U4003 = P1_U6752 & P1_U6751; 
assign P1_U5470 = ~(P1_U4215 & P1_U3257 & P1_GTE_485_U6); 
assign P1_U6149 = ~(P1_U4194 & P1_U2447 & P1_GTE_485_U6); 
assign P1_U6360 = ~(P1_U4204 & P1_GTE_485_U6); 
assign P1_U6808 = ~(P1_U2724 & P1_U6746); 
assign P1_U6812 = ~(P1_U2725 & P1_U6746); 
assign P1_U6816 = ~(P1_U2726 & P1_U6746); 
assign P1_U6825 = ~(P1_U2727 & P1_U6746); 
assign P1_U6829 = ~(P1_U2728 & P1_U6746); 
assign P1_U6833 = ~(P1_U2729 & P1_U6746); 
assign P1_U6837 = ~(P1_U2730 & P1_U6746); 
assign P1_U6882 = ~(P1_ADD_371_U24 & P1_U4208); 
assign P1_U7094 = ~P1_U3450; 
assign P1_U7096 = ~(P1_U3450 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P1_U7506 = ~(P1_U4116 & P1_U4115 & P1_U4114); 
assign P3_ADD_526_U76 = ~(P3_ADD_526_U192 & P3_ADD_526_U191); 
assign P3_ADD_526_U77 = ~(P3_ADD_526_U194 & P3_ADD_526_U193); 
assign P3_ADD_526_U117 = ~P3_ADD_526_U31; 
assign P3_ADD_526_U137 = ~P3_ADD_526_U107; 
assign P3_ADD_526_U188 = ~(P3_ADD_526_U31 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_526_U189 = ~(P3_ADD_526_U107 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_552_U76 = ~(P3_ADD_552_U192 & P3_ADD_552_U191); 
assign P3_ADD_552_U77 = ~(P3_ADD_552_U194 & P3_ADD_552_U193); 
assign P3_ADD_552_U117 = ~P3_ADD_552_U31; 
assign P3_ADD_552_U137 = ~P3_ADD_552_U107; 
assign P3_ADD_552_U188 = ~(P3_ADD_552_U31 & P3_EBX_REG_17__SCAN_IN); 
assign P3_ADD_552_U189 = ~(P3_ADD_552_U107 & P3_EBX_REG_16__SCAN_IN); 
assign P3_ADD_546_U76 = ~(P3_ADD_546_U192 & P3_ADD_546_U191); 
assign P3_ADD_546_U77 = ~(P3_ADD_546_U194 & P3_ADD_546_U193); 
assign P3_ADD_546_U117 = ~P3_ADD_546_U31; 
assign P3_ADD_546_U137 = ~P3_ADD_546_U107; 
assign P3_ADD_546_U188 = ~(P3_ADD_546_U31 & P3_EAX_REG_17__SCAN_IN); 
assign P3_ADD_546_U189 = ~(P3_ADD_546_U107 & P3_EAX_REG_16__SCAN_IN); 
assign P3_ADD_391_1180_U10 = ~(P3_U2615 & P3_ADD_391_1180_U29); 
assign P3_ADD_391_1180_U46 = ~(P3_ADD_391_1180_U29 & P3_ADD_391_1180_U9); 
assign P3_ADD_476_U62 = ~(P3_ADD_476_U124 & P3_ADD_476_U123); 
assign P3_ADD_476_U101 = ~P3_ADD_476_U20; 
assign P3_ADD_476_U181 = ~(P3_ADD_476_U20 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_531_U66 = ~(P3_ADD_531_U131 & P3_ADD_531_U130); 
assign P3_ADD_531_U105 = ~P3_ADD_531_U22; 
assign P3_ADD_531_U128 = ~(P3_ADD_531_U22 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_SUB_320_U24 = ~(P3_SUB_320_U25 & P3_SUB_320_U54 & P3_SUB_320_U85); 
assign P3_ADD_318_U62 = ~(P3_ADD_318_U124 & P3_ADD_318_U123); 
assign P3_ADD_318_U101 = ~P3_ADD_318_U20; 
assign P3_ADD_318_U181 = ~(P3_ADD_318_U20 & P3_PHYADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_315_U88 = ~(P3_ADD_315_U176 & P3_ADD_315_U175); 
assign P3_ADD_315_U98 = ~P3_ADD_315_U20; 
assign P3_ADD_315_U173 = ~(P3_ADD_315_U20 & P3_PHYADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_360_1242_U22 = ~P3_ADD_360_U20; 
assign P3_ADD_360_1242_U92 = P3_ADD_360_U20 & P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_360_1242_U118 = ~(P3_ADD_360_1242_U75 & P3_ADD_360_1242_U127); 
assign P3_ADD_360_1242_U133 = P3_ADD_360_U20 | P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_ADD_360_1242_U135 = ~(P3_ADD_360_U20 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_360_1242_U192 = ~(P3_ADD_360_1242_U122 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_360_1242_U226 = ~(P3_ADD_360_U20 & P3_ADD_360_1242_U23); 
assign P3_ADD_360_1242_U231 = ~(P3_ADD_360_1242_U29 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_360_1242_U233 = ~(P3_ADD_360_1242_U29 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_360_1242_U248 = ~(P3_ADD_360_1242_U246 & P3_ADD_360_1242_U28); 
assign P3_ADD_467_U62 = ~(P3_ADD_467_U124 & P3_ADD_467_U123); 
assign P3_ADD_467_U101 = ~P3_ADD_467_U20; 
assign P3_ADD_467_U181 = ~(P3_ADD_467_U20 & P3_REIP_REG_10__SCAN_IN); 
assign P3_ADD_430_U62 = ~(P3_ADD_430_U124 & P3_ADD_430_U123); 
assign P3_ADD_430_U101 = ~P3_ADD_430_U20; 
assign P3_ADD_430_U181 = ~(P3_ADD_430_U20 & P3_REIP_REG_10__SCAN_IN); 
assign P3_ADD_380_U66 = ~(P3_ADD_380_U131 & P3_ADD_380_U130); 
assign P3_ADD_380_U105 = ~P3_ADD_380_U22; 
assign P3_ADD_380_U128 = ~(P3_ADD_380_U22 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_344_U66 = ~(P3_ADD_344_U131 & P3_ADD_344_U130); 
assign P3_ADD_344_U105 = ~P3_ADD_344_U22; 
assign P3_ADD_344_U128 = ~(P3_ADD_344_U22 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_339_U62 = ~(P3_ADD_339_U124 & P3_ADD_339_U123); 
assign P3_ADD_339_U101 = ~P3_ADD_339_U20; 
assign P3_ADD_339_U181 = ~(P3_ADD_339_U20 & P3_PHYADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_360_U11 = ~(P3_U2625 & P3_ADD_360_U25); 
assign P3_ADD_360_U36 = ~(P3_ADD_360_U25 & P3_ADD_360_U10); 
assign P3_ADD_541_U62 = ~(P3_ADD_541_U124 & P3_ADD_541_U123); 
assign P3_ADD_541_U101 = ~P3_ADD_541_U20; 
assign P3_ADD_541_U181 = ~(P3_ADD_541_U20 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_SUB_357_1258_U32 = ~P3_ADD_357_U13; 
assign P3_SUB_357_1258_U35 = ~P3_ADD_357_U7; 
assign P3_SUB_357_1258_U66 = ~(P3_SUB_357_U7 & P3_SUB_357_1258_U161); 
assign P3_SUB_357_1258_U69 = ~(P3_SUB_357_1258_U484 & P3_SUB_357_1258_U483); 
assign P3_SUB_357_1258_U95 = P3_ADD_357_U7 & P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_SUB_357_1258_U159 = ~(P3_ADD_357_U13 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_SUB_357_1258_U163 = P3_ADD_357_U7 | P3_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P3_SUB_357_1258_U164 = P3_ADD_357_U13 | P3_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P3_SUB_357_1258_U181 = ~(P3_ADD_357_U7 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_SUB_357_1258_U185 = ~(P3_ADD_357_U7 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_SUB_357_1258_U270 = ~(P3_SUB_357_1258_U161 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_SUB_357_1258_U347 = ~(P3_ADD_357_U7 & P3_SUB_357_1258_U36); 
assign P3_SUB_357_1258_U363 = ~(P3_ADD_357_U13 & P3_SUB_357_1258_U33); 
assign P3_SUB_357_1258_U423 = ~(P3_SUB_357_1258_U161 & P3_SUB_357_1258_U34); 
assign P3_ADD_515_U62 = ~(P3_ADD_515_U124 & P3_ADD_515_U123); 
assign P3_ADD_515_U101 = ~P3_ADD_515_U20; 
assign P3_ADD_515_U181 = ~(P3_ADD_515_U20 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_394_U63 = ~(P3_ADD_394_U128 & P3_ADD_394_U127); 
assign P3_ADD_394_U104 = ~P3_ADD_394_U20; 
assign P3_ADD_394_U185 = ~(P3_ADD_394_U20 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_SUB_414_U78 = P3_SUB_414_U155 & P3_SUB_414_U154; 
assign P3_SUB_414_U96 = ~P3_SUB_414_U31; 
assign P3_SUB_414_U120 = ~(P3_SUB_414_U119 & P3_EBX_REG_16__SCAN_IN); 
assign P3_SUB_414_U152 = ~(P3_SUB_414_U31 & P3_EBX_REG_17__SCAN_IN); 
assign P3_ADD_441_U62 = ~(P3_ADD_441_U124 & P3_ADD_441_U123); 
assign P3_ADD_441_U101 = ~P3_ADD_441_U20; 
assign P3_ADD_441_U181 = ~(P3_ADD_441_U20 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_349_U66 = ~(P3_ADD_349_U131 & P3_ADD_349_U130); 
assign P3_ADD_349_U105 = ~P3_ADD_349_U22; 
assign P3_ADD_349_U128 = ~(P3_ADD_349_U22 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_405_U63 = ~(P3_ADD_405_U128 & P3_ADD_405_U127); 
assign P3_ADD_405_U104 = ~P3_ADD_405_U20; 
assign P3_ADD_405_U185 = ~(P3_ADD_405_U20 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_553_U66 = ~(P3_ADD_553_U131 & P3_ADD_553_U130); 
assign P3_ADD_553_U105 = ~P3_ADD_553_U22; 
assign P3_ADD_553_U128 = ~(P3_ADD_553_U22 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_558_U66 = ~(P3_ADD_558_U131 & P3_ADD_558_U130); 
assign P3_ADD_558_U105 = ~P3_ADD_558_U22; 
assign P3_ADD_558_U128 = ~(P3_ADD_558_U22 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_385_U66 = ~(P3_ADD_385_U131 & P3_ADD_385_U130); 
assign P3_ADD_385_U105 = ~P3_ADD_385_U22; 
assign P3_ADD_385_U128 = ~(P3_ADD_385_U22 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_357_U19 = P3_ADD_357_U33 & P3_ADD_357_U32; 
assign P3_ADD_357_U23 = ~P3_ADD_357_U12; 
assign P3_ADD_357_U27 = ~(P3_SUB_357_U9 & P3_ADD_357_U26); 
assign P3_ADD_357_U30 = ~(P3_SUB_357_U6 & P3_ADD_357_U12); 
assign P3_ADD_547_U66 = ~(P3_ADD_547_U131 & P3_ADD_547_U130); 
assign P3_ADD_547_U105 = ~P3_ADD_547_U22; 
assign P3_ADD_547_U128 = ~(P3_ADD_547_U22 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_371_1212_U120 = ~P3_ADD_371_1212_U77; 
assign P3_ADD_371_1212_U122 = ~(P3_ADD_371_1212_U35 & P3_ADD_371_1212_U34); 
assign P3_ADD_371_1212_U126 = ~P3_ADD_371_1212_U29; 
assign P3_ADD_371_1212_U199 = ~(P3_ADD_371_1212_U175 & P3_ADD_371_1212_U29); 
assign P3_ADD_371_1212_U201 = ~(P3_ADD_371_1212_U125 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_371_1212_U240 = ~(P3_ADD_371_1212_U26 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_ADD_371_1212_U253 = ~(P3_ADD_371_1212_U252 & P3_ADD_371_1212_U251); 
assign P3_ADD_371_U11 = ~(P3_U2625 & P3_ADD_371_U28); 
assign P3_ADD_371_U25 = P3_ADD_371_U42 & P3_ADD_371_U41; 
assign P3_ADD_371_U40 = ~(P3_ADD_371_U28 & P3_ADD_371_U10); 
assign P3_ADD_494_U62 = ~(P3_ADD_494_U124 & P3_ADD_494_U123); 
assign P3_ADD_494_U101 = ~P3_ADD_494_U20; 
assign P3_ADD_494_U181 = ~(P3_ADD_494_U20 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_536_U62 = ~(P3_ADD_536_U124 & P3_ADD_536_U123); 
assign P3_ADD_536_U101 = ~P3_ADD_536_U20; 
assign P3_ADD_536_U181 = ~(P3_ADD_536_U20 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_402_1132_U10 = ~(P3_U2615 & P3_ADD_402_1132_U29); 
assign P3_ADD_402_1132_U46 = ~(P3_ADD_402_1132_U29 & P3_ADD_402_1132_U9); 
assign P2_R2099_U9 = ~P2_U2746; 
assign P2_R2099_U11 = ~P2_U2745; 
assign P2_R2099_U13 = ~P2_U2744; 
assign P2_R2099_U14 = ~P2_U2743; 
assign P2_R2099_U16 = ~P2_U2742; 
assign P2_R2099_U18 = ~P2_U2741; 
assign P2_R2099_U20 = ~P2_U2740; 
assign P2_R2099_U22 = ~P2_U2739; 
assign P2_R2099_U23 = ~P2_U2738; 
assign P2_R2099_U26 = ~P2_U2737; 
assign P2_R2099_U28 = ~P2_U2736; 
assign P2_R2099_U30 = ~P2_U2735; 
assign P2_R2099_U32 = ~P2_U2734; 
assign P2_R2099_U34 = ~P2_U2733; 
assign P2_R2099_U36 = ~P2_U2732; 
assign P2_R2099_U38 = ~P2_U2731; 
assign P2_R2099_U40 = ~P2_U2730; 
assign P2_R2099_U42 = ~P2_U2729; 
assign P2_R2099_U44 = ~P2_U2728; 
assign P2_R2099_U46 = ~P2_U2727; 
assign P2_R2099_U48 = ~P2_U2726; 
assign P2_R2099_U50 = ~P2_U2725; 
assign P2_R2099_U52 = ~P2_U2724; 
assign P2_R2099_U54 = ~P2_U2723; 
assign P2_R2099_U56 = ~P2_U2722; 
assign P2_R2099_U58 = ~P2_U2721; 
assign P2_R2099_U60 = ~P2_U2720; 
assign P2_R2099_U62 = ~P2_U2719; 
assign P2_R2099_U64 = ~P2_U2718; 
assign P2_R2099_U66 = ~P2_U2717; 
assign P2_R2099_U101 = ~P2_U2716; 
assign P2_ADD_402_1132_U10 = ~(P2_U2593 & P2_ADD_402_1132_U29); 
assign P2_ADD_402_1132_U50 = ~(P2_ADD_402_1132_U29 & P2_ADD_402_1132_U9); 
assign P2_R2167_U14 = ~P2_U2703; 
assign P2_R2027_U66 = ~(P2_R2027_U131 & P2_R2027_U130); 
assign P2_R2027_U105 = ~P2_R2027_U22; 
assign P2_R2027_U128 = ~(P2_R2027_U22 & P2_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P2_R2337_U90 = ~(P2_R2337_U182 & P2_R2337_U181); 
assign P2_R2337_U102 = ~P2_R2337_U21; 
assign P2_R2337_U179 = ~(P2_R2337_U21 & P2_PHYADDRPOINTER_REG_11__SCAN_IN); 
assign P2_R2219_U6 = P2_R2219_U52 & P2_R2219_U48; 
assign P2_R2219_U8 = ~(P2_R2219_U45 & P2_R2219_U69); 
assign P2_R2219_U35 = ~(P2_R2219_U98 & P2_R2219_U97); 
assign P2_R2219_U36 = ~(P2_R2219_U103 & P2_R2219_U102); 
assign P2_R2219_U37 = ~(P2_R2219_U108 & P2_R2219_U107); 
assign P2_R2219_U38 = ~(P2_R2219_U113 & P2_R2219_U112); 
assign P2_R2219_U46 = ~P2_R2219_U45; 
assign P2_R2219_U72 = ~(P2_R2219_U53 & P2_R2219_U50); 
assign P2_R2219_U78 = ~(P2_R2219_U47 & P2_R2219_U45); 
assign P2_R2219_U80 = ~(P2_R2219_U77 & P2_R2219_U45); 
assign P2_R2096_U68 = ~(P2_R2096_U265 & P2_R2096_U264); 
assign P2_R2096_U100 = P2_R2096_U176 & P2_R2096_U175; 
assign P2_R2096_U102 = P2_R2096_U183 & P2_R2096_U182; 
assign P2_R2096_U104 = P2_R2096_U190 & P2_R2096_U189; 
assign P2_R2096_U106 = P2_R2096_U197 & P2_R2096_U196; 
assign P2_R2096_U108 = P2_R2096_U204 & P2_R2096_U203; 
assign P2_R2096_U110 = P2_R2096_U213 & P2_R2096_U212; 
assign P2_R2096_U118 = ~(P2_U2648 & P2_R2096_U117); 
assign P2_R2096_U179 = ~(P2_R2096_U178 & P2_R2096_U177); 
assign P2_R2096_U186 = ~(P2_R2096_U185 & P2_R2096_U184); 
assign P2_R2096_U193 = ~(P2_R2096_U192 & P2_R2096_U191); 
assign P2_R2096_U200 = ~(P2_R2096_U199 & P2_R2096_U198); 
assign P2_R2096_U207 = ~(P2_R2096_U206 & P2_R2096_U205); 
assign P2_R2096_U216 = ~(P2_R2096_U215 & P2_R2096_U214); 
assign P2_R2096_U240 = ~(P2_R2096_U169 & P2_R2096_U54); 
assign P2_R2096_U243 = ~(P2_R2096_U115 & P2_U2648); 
assign P2_R1957_U24 = ~(P2_R1957_U85 & P2_R1957_U54 & P2_R1957_U25); 
assign P2_R2088_U7 = ~(P2_U3648 | P2_U3649 | P2_U3650 | P2_U3652 | P2_U3651); 
assign P2_ADD_394_U70 = ~(P2_ADD_394_U142 & P2_ADD_394_U141); 
assign P2_ADD_394_U104 = ~P2_ADD_394_U20; 
assign P2_ADD_394_U167 = ~(P2_ADD_394_U20 & P2_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P1_R2027_U76 = ~(P1_R2027_U192 & P1_R2027_U191); 
assign P1_R2027_U77 = ~(P1_R2027_U194 & P1_R2027_U193); 
assign P1_R2027_U117 = ~P1_R2027_U31; 
assign P1_R2027_U137 = ~P1_R2027_U107; 
assign P1_R2027_U188 = ~(P1_R2027_U31 & P1_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P1_R2027_U189 = ~(P1_R2027_U107 & P1_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P1_R2182_U14 = ~P1_U2737; 
assign P1_R2182_U15 = ~P1_U2738; 
assign P1_R2182_U16 = ~(P1_U2723 & P1_U2739); 
assign P1_R2182_U17 = ~P1_U2736; 
assign P1_R2182_U18 = ~P1_U2735; 
assign P1_R2182_U20 = ~P1_U2734; 
assign P1_R2182_U23 = ~P1_U2733; 
assign P1_R2182_U36 = P1_U2738 & P1_U2737; 
assign P1_R2182_U37 = P1_U2735 & P1_U2736; 
assign P1_R2182_U39 = ~P1_U2732; 
assign P1_R2182_U60 = P1_U2739 | P1_U2723; 
assign P1_R2144_U6 = P1_R2144_U36 & P1_R2144_U35 & P1_R2144_U27 & P1_R2144_U29; 
assign P1_R2144_U64 = P1_R2144_U34 & P1_R2144_U33 & P1_R2144_U31 & P1_R2144_U32; 
assign P1_R2144_U65 = P1_R2144_U34 & P1_R2144_U33; 
assign P1_R2144_U66 = P1_R2144_U36 & P1_R2144_U27 & P1_R2144_U29; 
assign P1_R2144_U67 = P1_R2144_U29 & P1_R2144_U27; 
assign P1_R2144_U68 = ~P1_U2762; 
assign P1_R2144_U69 = ~P1_U2761; 
assign P1_R2144_U70 = ~P1_U2763; 
assign P1_R2144_U71 = ~P1_U2764; 
assign P1_R2144_U165 = ~(P1_U2762 & P1_R2144_U12); 
assign P1_R2144_U167 = ~(P1_U2761 & P1_R2144_U12); 
assign P1_R2144_U169 = ~(P1_U2763 & P1_R2144_U12); 
assign P1_R2144_U172 = ~(P1_U2762 & P1_R2144_U12); 
assign P1_R2144_U175 = ~(P1_U2763 & P1_R2144_U12); 
assign P1_R2144_U177 = ~(P1_U2764 & P1_R2144_U12); 
assign P1_R2144_U180 = ~(P1_U2761 & P1_R2144_U12); 
assign P1_R2144_U201 = ~(P1_U2764 & P1_R2144_U12); 
assign P1_R2144_U204 = ~P1_R2144_U29; 
assign P1_R2144_U207 = ~P1_R2144_U27; 
assign P1_R2144_U222 = ~P1_R2144_U32; 
assign P1_R2144_U225 = ~P1_R2144_U31; 
assign P1_R2144_U228 = ~P1_R2144_U33; 
assign P1_R2144_U231 = ~P1_R2144_U34; 
assign P1_R2144_U234 = ~P1_R2144_U35; 
assign P1_R2144_U237 = ~P1_R2144_U36; 
assign P1_R2358_U144 = ~P1_U2615; 
assign P1_R2358_U405 = ~(P1_U2615 & P1_R2358_U23); 
assign P1_R2358_U408 = ~(P1_R2358_U407 & P1_R2358_U406); 
assign P1_R2358_U420 = ~(P1_U2615 & P1_R2358_U23); 
assign P1_R2099_U140 = ~(P1_R2099_U148 & P1_R2099_U147); 
assign P1_R2099_U150 = ~(P1_R2099_U190 & P1_R2099_U6); 
assign P1_R2099_U318 = ~(P1_R2099_U190 & P1_U2678); 
assign P1_R2099_U320 = ~(P1_R2099_U190 & P1_U2678); 
assign P1_R2099_U349 = ~(P1_R2099_U98 & P1_R2099_U187); 
assign P1_R2167_U6 = ~P1_U2716; 
assign P1_R2167_U13 = ~P1_U2717; 
assign P1_R2167_U14 = ~P1_U2711; 
assign P1_R2167_U18 = P1_R2167_U29 & P1_R2167_U30; 
assign P1_R2167_U28 = ~(P1_R2167_U27 & P1_R2167_U26 & P1_R2167_U25 & P1_R2167_U24); 
assign P1_R2167_U33 = ~(P1_U2712 & P1_R2167_U12); 
assign P1_R2167_U41 = ~(P1_U2716 & P1_R2167_U15); 
assign P1_R2167_U43 = ~(P1_U2716 & P1_R2167_U16); 
assign P1_R2337_U62 = ~(P1_R2337_U124 & P1_R2337_U123); 
assign P1_R2337_U101 = ~P1_R2337_U20; 
assign P1_R2337_U181 = ~(P1_R2337_U20 & P1_PHYADDRPOINTER_REG_10__SCAN_IN); 
assign P1_R2096_U62 = ~(P1_R2096_U124 & P1_R2096_U123); 
assign P1_R2096_U101 = ~P1_R2096_U20; 
assign P1_R2096_U181 = ~(P1_R2096_U20 & P1_REIP_REG_10__SCAN_IN); 
assign P1_ADD_371_U18 = ~(P1_ADD_371_U36 & P1_ADD_371_U35); 
assign P1_ADD_371_U29 = ~P1_ADD_371_U11; 
assign P1_ADD_371_U37 = ~(P1_U3232 & P1_ADD_371_U11); 
assign P1_ADD_405_U70 = ~(P1_ADD_405_U142 & P1_ADD_405_U141); 
assign P1_ADD_405_U104 = ~P1_ADD_405_U20; 
assign P1_ADD_405_U167 = ~(P1_ADD_405_U20 & P1_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P1_ADD_515_U70 = ~(P1_ADD_515_U140 & P1_ADD_515_U139); 
assign P1_ADD_515_U101 = ~P1_ADD_515_U20; 
assign P1_ADD_515_U165 = ~(P1_ADD_515_U20 & P1_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_U2863 = ~(P3_U5616 & P3_U5615); 
assign P3_U2864 = ~(P3_U5610 & P3_U5609); 
assign P3_U2865 = ~(P3_U5599 & P3_U5598); 
assign P3_U3145 = ~(P3_U3144 & P3_U4667); 
assign P3_U3151 = ~(P3_U3149 & P3_U4719); 
assign P3_U3159 = ~(P3_U3157 & P3_U4771); 
assign P3_U3163 = ~(P3_U3162 & P3_U4822); 
assign P3_U3167 = ~(P3_U3166 & P3_U4874); 
assign P3_U3171 = ~(P3_U3170 & P3_U4926); 
assign P3_U3175 = ~(P3_U3174 & P3_U4978); 
assign P3_U3179 = ~(P3_U3178 & P3_U5029); 
assign P3_U3183 = ~(P3_U2504 & P3_U4647); 
assign P3_U3187 = ~(P3_U2504 & P3_U2490); 
assign P3_U3191 = ~(P3_U2504 & P3_U2493); 
assign P3_U3195 = ~(P3_U2504 & P3_U2495); 
assign P3_U3197 = ~(P3_U2508 & P3_U4647); 
assign P3_U3200 = ~(P3_U2508 & P3_U2490); 
assign P3_U3203 = ~(P3_U2508 & P3_U2493); 
assign P3_U3206 = ~(P3_U2508 & P3_U2495); 
assign P3_U3244 = ~(P3_U4352 & P3_U4522); 
assign P3_U3245 = ~(P3_U4352 & P3_U3102); 
assign P3_U3254 = ~(P3_U5490 & P3_U5489); 
assign P3_U3255 = ~(P3_U5487 & P3_U5486); 
assign P3_U3656 = P3_U5495 & P3_U4333; 
assign P3_U3677 = P3_U5540 & P3_U5541; 
assign P3_U3682 = P3_U5565 & P3_U5564; 
assign P3_U3687 = P3_U5625 & P3_U4333 & P3_U5626; 
assign P3_U3697 = P3_U5648 & P3_U5649 & P3_U5647 & P3_U5651 & P3_U5650; 
assign P3_U3748 = P3_U3749 & P3_U5809; 
assign P3_U4609 = ~(P3_U2361 & P3_U3238); 
assign P3_U4610 = ~(P3_U2360 & P3_U3237); 
assign P3_U4611 = ~(P3_U2357 & P3_U3212); 
assign P3_U4612 = ~(P3_U4305 & P3_U3215); 
assign P3_U4613 = ~(P3_U4304 & P3_U3210); 
assign P3_U4614 = ~(P3_U4303 & P3_U3213); 
assign P3_U4615 = ~(P3_U2356 & P3_U3211); 
assign P3_U4616 = ~(P3_U4302 & P3_U3214); 
assign P3_U4661 = ~P3_U3144; 
assign P3_U4715 = ~P3_U3149; 
assign P3_U4767 = ~P3_U3157; 
assign P3_U4819 = ~P3_U3162; 
assign P3_U4870 = ~P3_U3166; 
assign P3_U4922 = ~P3_U3170; 
assign P3_U4974 = ~P3_U3174; 
assign P3_U5026 = ~P3_U3178; 
assign P3_U5525 = ~P3_U3221; 
assign P3_U5619 = ~(P3_U5618 & P3_U5617); 
assign P3_U5622 = ~(P3_U5621 & P3_U5620); 
assign P3_U5633 = ~(P3_SUB_357_1258_U69 & P3_U2393); 
assign P3_U5636 = ~(P3_U4299 & P3_ADD_547_U5); 
assign P3_U5660 = ~(P3_ADD_547_U85 & P3_U4299); 
assign P3_U5684 = ~(P3_ADD_547_U74 & P3_U4299); 
assign P3_U5708 = ~(P3_ADD_547_U71 & P3_U4299); 
assign P3_U5732 = ~(P3_ADD_547_U70 & P3_U4299); 
assign P3_U5756 = ~(P3_ADD_547_U69 & P3_U4299); 
assign P3_U5780 = ~(P3_ADD_547_U68 & P3_U4299); 
assign P3_U5804 = ~(P3_ADD_547_U67 & P3_U4299); 
assign P3_U5827 = ~(P3_ADD_553_U66 & P3_U4298); 
assign P3_U5828 = ~(P3_ADD_547_U66 & P3_U4299); 
assign P3_U5831 = ~(P3_ADD_531_U66 & P3_U2354); 
assign P3_U5839 = ~(P3_ADD_385_U66 & P3_U2358); 
assign P3_U5840 = ~(P3_ADD_380_U66 & P3_U2359); 
assign P3_U5841 = ~(P3_ADD_349_U66 & P3_U4306); 
assign P3_U5842 = ~(P3_ADD_344_U66 & P3_U2362); 
assign P3_U5857 = ~(P3_ADD_515_U62 & P3_U4302); 
assign P3_U5858 = ~(P3_ADD_494_U62 & P3_U2356); 
assign P3_U5859 = ~(P3_ADD_476_U62 & P3_U4303); 
assign P3_U5860 = ~(P3_ADD_441_U62 & P3_U4304); 
assign P3_U5861 = ~(P3_ADD_405_U63 & P3_U4305); 
assign P3_U5862 = ~(P3_ADD_394_U63 & P3_U2357); 
assign P3_U5976 = ~(P3_ADD_526_U77 & P3_U2355); 
assign P3_U6000 = ~(P3_ADD_526_U76 & P3_U2355); 
assign P3_U6401 = ~(P3_U6400 & P3_U6399); 
assign P3_U6663 = ~(P3_U6662 & P3_U6661); 
assign P3_U6997 = ~(P3_U3242 & P3_U6996); 
assign P3_U7942 = ~(P3_U4505 & P3_U3211); 
assign P3_U7943 = ~(P3_U3104 & P3_U3214); 
assign P3_U7944 = ~(P3_U4505 & P3_U3213); 
assign P3_U7945 = ~(P3_U3104 & P3_U3210); 
assign P3_U7950 = ~(P3_U4505 & P3_U3237); 
assign P3_U7951 = ~(P3_U3104 & P3_U3238); 
assign P3_U7975 = ~(P3_U4539 & P3_U5512); 
assign P3_U7981 = ~(P3_U3221 & P3_U3094 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_U7993 = ~(P3_U3221 & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P2_U2747 = ~(P2_U7886 & P2_U7721 & P2_U4389 & P2_U4388 & P2_U7717); 
assign P2_U2748 = ~(P2_U7583 & P2_U7582); 
assign P2_U2749 = ~(P2_U4380 & P2_U7584); 
assign P2_U2750 = ~(P2_U4382 & P2_U7588); 
assign P2_U4408 = ~P2_R2219_U8; 
assign P2_U5663 = ~(P2_R2096_U68 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U8345 = ~(P2_R2219_U8 & P2_U2617); 
assign P2_U8417 = ~(P2_R2337_U90 & P2_U3284); 
assign P1_U2617 = ~(P1_U6750 & P1_U4003); 
assign P1_U2741 = ~(P1_U4078 & P1_U7096); 
assign P1_U2743 = P1_U7506 & P1_U7470; 
assign P1_U3737 = P1_U3736 & P1_U5470; 
assign P1_U4498 = ~(P1_U4477 & P1_U3388); 
assign P1_U4507 = ~(P1_U4215 & P1_U3388); 
assign P1_U5569 = ~(P1_U3758 & P1_U2519); 
assign P1_U6749 = ~(P1_R2337_U62 & P1_U2352); 
assign P1_U6880 = ~(P1_ADD_371_U18 & P1_U4208); 
assign P1_U7492 = ~(P1_U4109 & P1_U7094); 
assign P1_U7509 = ~(P1_U3746 & P1_U2519); 
assign P1_U7740 = ~(P1_U4477 & P1_U3388); 
assign P3_ADD_526_U34 = ~(P3_ADD_526_U89 & P3_ADD_526_U117); 
assign P3_ADD_526_U106 = ~(P3_ADD_526_U117 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_526_U187 = ~(P3_ADD_526_U117 & P3_ADD_526_U30); 
assign P3_ADD_526_U190 = ~(P3_ADD_526_U137 & P3_ADD_526_U28); 
assign P3_ADD_552_U34 = ~(P3_ADD_552_U89 & P3_ADD_552_U117); 
assign P3_ADD_552_U106 = ~(P3_ADD_552_U117 & P3_EBX_REG_17__SCAN_IN); 
assign P3_ADD_552_U187 = ~(P3_ADD_552_U117 & P3_ADD_552_U30); 
assign P3_ADD_552_U190 = ~(P3_ADD_552_U137 & P3_ADD_552_U28); 
assign P3_ADD_546_U34 = ~(P3_ADD_546_U89 & P3_ADD_546_U117); 
assign P3_ADD_546_U106 = ~(P3_ADD_546_U117 & P3_EAX_REG_17__SCAN_IN); 
assign P3_ADD_546_U187 = ~(P3_ADD_546_U117 & P3_ADD_546_U30); 
assign P3_ADD_546_U190 = ~(P3_ADD_546_U137 & P3_ADD_546_U28); 
assign P3_ADD_391_1180_U23 = ~(P3_ADD_391_1180_U46 & P3_ADD_391_1180_U45); 
assign P3_ADD_391_1180_U30 = ~P3_ADD_391_1180_U10; 
assign P3_ADD_391_1180_U43 = ~(P3_U2616 & P3_ADD_391_1180_U10); 
assign P3_ADD_476_U22 = ~(P3_ADD_476_U101 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_476_U182 = ~(P3_ADD_476_U101 & P3_ADD_476_U21); 
assign P3_ADD_531_U23 = ~(P3_ADD_531_U105 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_531_U129 = ~(P3_ADD_531_U105 & P3_ADD_531_U21); 
assign P3_SUB_320_U20 = P3_SUB_320_U88 & P3_SUB_320_U24; 
assign P3_SUB_320_U52 = ~P3_ADD_318_U62; 
assign P3_SUB_320_U86 = ~P3_SUB_320_U24; 
assign P3_SUB_320_U128 = ~(P3_ADD_318_U62 & P3_SUB_320_U24); 
assign P3_ADD_318_U22 = ~(P3_ADD_318_U101 & P3_PHYADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_318_U182 = ~(P3_ADD_318_U101 & P3_ADD_318_U21); 
assign P3_ADD_315_U22 = ~(P3_ADD_315_U98 & P3_PHYADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_315_U174 = ~(P3_ADD_315_U98 & P3_ADD_315_U21); 
assign P3_ADD_360_1242_U19 = ~(P3_ADD_360_1242_U248 & P3_ADD_360_1242_U247 & P3_ADD_360_1242_U192); 
assign P3_ADD_360_1242_U117 = P3_ADD_360_1242_U232 & P3_ADD_360_1242_U231; 
assign P3_ADD_360_1242_U128 = ~P3_ADD_360_1242_U118; 
assign P3_ADD_360_1242_U130 = ~(P3_ADD_360_1242_U129 & P3_ADD_360_1242_U118); 
assign P3_ADD_360_1242_U225 = ~(P3_ADD_360_1242_U22 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_360_1242_U235 = ~(P3_ADD_360_1242_U234 & P3_ADD_360_1242_U233); 
assign P3_ADD_467_U22 = ~(P3_ADD_467_U101 & P3_REIP_REG_10__SCAN_IN); 
assign P3_ADD_467_U182 = ~(P3_ADD_467_U101 & P3_ADD_467_U21); 
assign P3_ADD_430_U22 = ~(P3_ADD_430_U101 & P3_REIP_REG_10__SCAN_IN); 
assign P3_ADD_430_U182 = ~(P3_ADD_430_U101 & P3_ADD_430_U21); 
assign P3_ADD_380_U23 = ~(P3_ADD_380_U105 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_380_U129 = ~(P3_ADD_380_U105 & P3_ADD_380_U21); 
assign P3_ADD_344_U23 = ~(P3_ADD_344_U105 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_344_U129 = ~(P3_ADD_344_U105 & P3_ADD_344_U21); 
assign P3_ADD_339_U22 = ~(P3_ADD_339_U101 & P3_PHYADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_339_U182 = ~(P3_ADD_339_U101 & P3_ADD_339_U21); 
assign P3_ADD_360_U19 = ~(P3_ADD_360_U36 & P3_ADD_360_U35); 
assign P3_ADD_360_U26 = ~P3_ADD_360_U11; 
assign P3_ADD_360_U33 = ~(P3_U2626 & P3_ADD_360_U11); 
assign P3_ADD_541_U22 = ~(P3_ADD_541_U101 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_541_U182 = ~(P3_ADD_541_U101 & P3_ADD_541_U21); 
assign P3_SUB_357_1258_U26 = ~P3_ADD_357_U19; 
assign P3_SUB_357_1258_U97 = P3_SUB_357_1258_U164 & P3_SUB_357_1258_U163; 
assign P3_SUB_357_1258_U127 = ~(P3_SUB_357_1258_U270 & P3_SUB_357_1258_U66 & P3_SUB_357_1258_U271); 
assign P3_SUB_357_1258_U158 = ~P3_SUB_357_1258_U66; 
assign P3_SUB_357_1258_U160 = P3_ADD_357_U19 | P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_SUB_357_1258_U162 = ~(P3_ADD_357_U19 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_SUB_357_1258_U166 = ~(P3_SUB_357_1258_U271 & P3_SUB_357_1258_U270 & P3_SUB_357_1258_U159 & P3_SUB_357_1258_U66); 
assign P3_SUB_357_1258_U260 = ~(P3_SUB_357_1258_U185 & P3_SUB_357_1258_U163); 
assign P3_SUB_357_1258_U261 = ~(P3_SUB_357_1258_U164 & P3_SUB_357_1258_U159); 
assign P3_SUB_357_1258_U342 = ~(P3_ADD_357_U19 & P3_SUB_357_1258_U27); 
assign P3_SUB_357_1258_U346 = ~(P3_SUB_357_1258_U35 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_SUB_357_1258_U362 = ~(P3_SUB_357_1258_U32 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_SUB_357_1258_U424 = ~(P3_SUB_357_1258_U423 & P3_SUB_357_1258_U422); 
assign P3_ADD_515_U22 = ~(P3_ADD_515_U101 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_515_U182 = ~(P3_ADD_515_U101 & P3_ADD_515_U21); 
assign P3_ADD_394_U22 = ~(P3_ADD_394_U104 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_394_U186 = ~(P3_ADD_394_U104 & P3_ADD_394_U21); 
assign P3_SUB_414_U9 = P3_SUB_414_U120 & P3_SUB_414_U31; 
assign P3_SUB_414_U32 = ~(P3_SUB_414_U45 & P3_SUB_414_U75 & P3_SUB_414_U96); 
assign P3_SUB_414_U117 = ~(P3_SUB_414_U96 & P3_SUB_414_U75); 
assign P3_SUB_414_U153 = ~(P3_SUB_414_U96 & P3_SUB_414_U75); 
assign P3_ADD_441_U22 = ~(P3_ADD_441_U101 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_441_U182 = ~(P3_ADD_441_U101 & P3_ADD_441_U21); 
assign P3_ADD_349_U23 = ~(P3_ADD_349_U105 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_349_U129 = ~(P3_ADD_349_U105 & P3_ADD_349_U21); 
assign P3_ADD_405_U22 = ~(P3_ADD_405_U104 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_405_U186 = ~(P3_ADD_405_U104 & P3_ADD_405_U21); 
assign P3_ADD_553_U23 = ~(P3_ADD_553_U105 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_553_U129 = ~(P3_ADD_553_U105 & P3_ADD_553_U21); 
assign P3_ADD_558_U23 = ~(P3_ADD_558_U105 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_558_U129 = ~(P3_ADD_558_U105 & P3_ADD_558_U21); 
assign P3_ADD_385_U23 = ~(P3_ADD_385_U105 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_385_U129 = ~(P3_ADD_385_U105 & P3_ADD_385_U21); 
assign P3_ADD_357_U6 = ~(P3_ADD_357_U15 & P3_ADD_357_U23); 
assign P3_ADD_357_U8 = P3_ADD_357_U27 & P3_ADD_357_U12; 
assign P3_ADD_357_U24 = ~(P3_ADD_357_U23 & P3_ADD_357_U16); 
assign P3_ADD_357_U31 = ~(P3_ADD_357_U23 & P3_ADD_357_U16); 
assign P3_ADD_547_U23 = ~(P3_ADD_547_U105 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_547_U129 = ~(P3_ADD_547_U105 & P3_ADD_547_U21); 
assign P3_ADD_371_1212_U30 = ~P3_ADD_371_U25; 
assign P3_ADD_371_1212_U123 = ~(P3_ADD_371_1212_U122 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_371_1212_U129 = ~(P3_ADD_371_U25 & P3_ADD_371_1212_U126); 
assign P3_ADD_371_1212_U161 = ~(P3_ADD_371_U25 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_371_1212_U202 = ~(P3_ADD_371_U25 & P3_ADD_371_1212_U125); 
assign P3_ADD_371_1212_U203 = ~(P3_ADD_371_1212_U120 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_ADD_371_1212_U235 = ~(P3_ADD_371_U25 & P3_ADD_371_1212_U28); 
assign P3_ADD_371_1212_U242 = ~(P3_ADD_371_1212_U241 & P3_ADD_371_1212_U240); 
assign P3_ADD_371_1212_U255 = ~(P3_ADD_371_1212_U253 & P3_ADD_371_1212_U35); 
assign P3_ADD_371_U20 = ~(P3_ADD_371_U40 & P3_ADD_371_U39); 
assign P3_ADD_371_U29 = ~P3_ADD_371_U11; 
assign P3_ADD_371_U37 = ~(P3_U2626 & P3_ADD_371_U11); 
assign P3_ADD_494_U22 = ~(P3_ADD_494_U101 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_494_U182 = ~(P3_ADD_494_U101 & P3_ADD_494_U21); 
assign P3_ADD_536_U22 = ~(P3_ADD_536_U101 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_536_U182 = ~(P3_ADD_536_U101 & P3_ADD_536_U21); 
assign P3_ADD_402_1132_U23 = ~(P3_ADD_402_1132_U46 & P3_ADD_402_1132_U45); 
assign P3_ADD_402_1132_U30 = ~P3_ADD_402_1132_U10; 
assign P3_ADD_402_1132_U43 = ~(P3_U2616 & P3_ADD_402_1132_U10); 
assign P2_R2099_U7 = ~P2_U2751; 
assign P2_ADD_391_1196_U19 = ~P2_R2096_U68; 
assign P2_ADD_402_1132_U25 = ~(P2_ADD_402_1132_U50 & P2_ADD_402_1132_U49); 
assign P2_ADD_402_1132_U30 = ~P2_ADD_402_1132_U10; 
assign P2_ADD_402_1132_U41 = ~(P2_U2594 & P2_ADD_402_1132_U10); 
assign P2_R2182_U52 = ~P2_U2689; 
assign P2_R2182_U54 = ~P2_U2688; 
assign P2_R2182_U155 = P2_U2689 | P2_U2665; 
assign P2_R2182_U157 = ~(P2_U2665 & P2_U2689); 
assign P2_R2182_U159 = P2_U2688 | P2_U2664; 
assign P2_R2182_U161 = ~(P2_U2664 & P2_U2688); 
assign P2_R2182_U260 = ~(P2_U2688 & P2_R2182_U55); 
assign P2_R2182_U262 = ~(P2_U2688 & P2_R2182_U55); 
assign P2_R2182_U267 = ~(P2_U2689 & P2_R2182_U53); 
assign P2_R2182_U269 = ~(P2_U2689 & P2_R2182_U53); 
assign P2_R2027_U23 = ~(P2_R2027_U105 & P2_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P2_R2027_U129 = ~(P2_R2027_U105 & P2_R2027_U21); 
assign P2_R2337_U23 = ~(P2_R2337_U102 & P2_PHYADDRPOINTER_REG_11__SCAN_IN); 
assign P2_R2337_U180 = ~(P2_R2337_U102 & P2_R2337_U22); 
assign P2_R2219_U19 = ~(P2_R2219_U72 & P2_R2219_U76); 
assign P2_R2219_U31 = P2_R2219_U6 & P2_R2219_U55; 
assign P2_R2219_U44 = ~(P2_R2219_U78 & P2_R2219_U70); 
assign P2_R2219_U81 = ~(P2_R2219_U80 & P2_R2219_U70); 
assign P2_R2219_U99 = ~P2_R2219_U35; 
assign P2_R2219_U104 = ~P2_R2219_U36; 
assign P2_R2219_U109 = ~P2_R2219_U37; 
assign P2_R2219_U114 = ~P2_R2219_U38; 
assign P2_R2219_U116 = ~(P2_R2219_U38 & P2_R2219_U45); 
assign P2_R2096_U111 = ~(P2_R2096_U113 & P2_R2096_U118); 
assign P2_R2096_U114 = P2_R2096_U243 & P2_R2096_U242; 
assign P2_R2096_U241 = ~(P2_R2096_U240 & P2_R2096_U239); 
assign P2_R1957_U20 = P2_R1957_U88 & P2_R1957_U24; 
assign P2_R1957_U52 = ~P2_U3653; 
assign P2_R1957_U86 = ~P2_R1957_U24; 
assign P2_R1957_U128 = ~(P2_U3653 & P2_R1957_U24); 
assign P2_R2088_U6 = ~(P2_U3648 | P2_R2088_U7); 
assign P2_ADD_394_U22 = ~(P2_ADD_394_U104 & P2_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P2_ADD_394_U168 = ~(P2_ADD_394_U104 & P2_ADD_394_U21); 
assign P1_R2027_U34 = ~(P1_R2027_U89 & P1_R2027_U117); 
assign P1_R2027_U106 = ~(P1_R2027_U117 & P1_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P1_R2027_U187 = ~(P1_R2027_U117 & P1_R2027_U30); 
assign P1_R2027_U190 = ~(P1_R2027_U137 & P1_R2027_U28); 
assign P1_R2182_U6 = P1_R2182_U60 & P1_R2182_U16; 
assign P1_R2182_U7 = ~P1_U2744; 
assign P1_R2182_U8 = ~P1_U3246; 
assign P1_R2182_U9 = ~(P1_U3246 & P1_U2744); 
assign P1_R2182_U49 = ~P1_R2182_U16; 
assign P1_R2182_U82 = ~(P1_U2738 & P1_R2182_U16); 
assign P1_R2144_U63 = P1_R2144_U6 & P1_R2144_U64; 
assign P1_R2144_U164 = ~(P1_U2355 & P1_R2144_U68); 
assign P1_R2144_U166 = ~(P1_U2355 & P1_R2144_U69); 
assign P1_R2144_U168 = ~(P1_U2355 & P1_R2144_U70); 
assign P1_R2144_U171 = ~(P1_U2355 & P1_R2144_U68); 
assign P1_R2144_U174 = ~(P1_U2355 & P1_R2144_U70); 
assign P1_R2144_U176 = ~(P1_U2355 & P1_R2144_U71); 
assign P1_R2144_U179 = ~(P1_U2355 & P1_R2144_U69); 
assign P1_R2144_U200 = ~(P1_U2355 & P1_R2144_U71); 
assign P1_R2358_U404 = ~(P1_U2352 & P1_R2358_U144); 
assign P1_R2358_U419 = ~(P1_U2352 & P1_R2358_U144); 
assign P1_R2099_U86 = ~(P1_R2099_U349 & P1_R2099_U348); 
assign P1_R2099_U139 = P1_R2099_U319 & P1_R2099_U318; 
assign P1_R2099_U149 = ~P1_R2099_U140; 
assign P1_R2099_U151 = ~(P1_R2099_U150 & P1_R2099_U140); 
assign P1_R2099_U322 = ~(P1_R2099_U321 & P1_R2099_U320); 
assign P1_R2167_U19 = P1_R2167_U32 & P1_R2167_U33; 
assign P1_R2167_U31 = ~(P1_R2167_U18 & P1_R2167_U28); 
assign P1_R2167_U36 = ~(P1_U2717 & P1_R2167_U14); 
assign P1_R2167_U38 = ~(P1_U2711 & P1_R2167_U13); 
assign P1_R2167_U39 = ~(P1_U2356 & P1_R2167_U6); 
assign P1_R2167_U46 = ~(P1_R2167_U6 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_R2337_U22 = ~(P1_R2337_U101 & P1_PHYADDRPOINTER_REG_10__SCAN_IN); 
assign P1_R2337_U182 = ~(P1_R2337_U101 & P1_R2337_U21); 
assign P1_R2096_U22 = ~(P1_R2096_U101 & P1_REIP_REG_10__SCAN_IN); 
assign P1_R2096_U182 = ~(P1_R2096_U101 & P1_R2096_U21); 
assign P1_ADD_371_U14 = ~(P1_U3232 & P1_ADD_371_U29); 
assign P1_ADD_371_U38 = ~(P1_ADD_371_U29 & P1_ADD_371_U12); 
assign P1_ADD_405_U22 = ~(P1_ADD_405_U104 & P1_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P1_ADD_405_U168 = ~(P1_ADD_405_U104 & P1_ADD_405_U21); 
assign P1_ADD_515_U22 = ~(P1_ADD_515_U101 & P1_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P1_ADD_515_U166 = ~(P1_ADD_515_U101 & P1_ADD_515_U21); 
assign P3_U3184 = ~(P3_U3183 & P3_U3181); 
assign P3_U3188 = ~(P3_U3187 & P3_U5130); 
assign P3_U3192 = ~(P3_U3191 & P3_U5182); 
assign P3_U3220 = ~(P3_U7976 & P3_U7975 & P3_U3667); 
assign P3_U3250 = ~(P3_U2390 & P3_U6663); 
assign P3_U3253 = ~(P3_U2390 & P3_U6997); 
assign P3_U3357 = P3_U4612 & P3_U4611 & P3_U4610 & P3_U4609; 
assign P3_U3358 = P3_U4616 & P3_U4615 & P3_U4614 & P3_U4613; 
assign P3_U3672 = P3_U3245 & P3_U3244 & P3_U3671; 
assign P3_U3692 = P3_U5636 & P3_U5635; 
assign P3_U3698 = P3_U3697 & P3_U3696; 
assign P3_U3699 = P3_U5660 & P3_U5659; 
assign P3_U3707 = P3_U5684 & P3_U5683; 
assign P3_U3715 = P3_U5708 & P3_U5707; 
assign P3_U3723 = P3_U5732 & P3_U5731; 
assign P3_U3731 = P3_U5756 & P3_U5755; 
assign P3_U3739 = P3_U5780 & P3_U5779; 
assign P3_U3747 = P3_U5804 & P3_U5803; 
assign P3_U3755 = P3_U5828 & P3_U5827; 
assign P3_U3756 = P3_U5833 & P3_U5832 & P3_U5831; 
assign P3_U3759 = P3_U5842 & P3_U5841 & P3_U5840 & P3_U5839; 
assign P3_U3763 = P3_U5857 & P3_U5856; 
assign P3_U3765 = P3_U5859 & P3_U5858 & P3_U5860 & P3_U5862 & P3_U5861; 
assign P3_U4280 = P3_U7943 & P3_U7942; 
assign P3_U4282 = P3_U7951 & P3_U7950; 
assign P3_U4300 = ~P3_U3244; 
assign P3_U4301 = ~P3_U3245; 
assign P3_U4618 = ~(P3_U2463 & P3_U4522 & P3_U3360 & P3_U7945 & P3_U7944); 
assign P3_U4668 = ~P3_U3145; 
assign P3_U4669 = ~(P3_U2489 & P3_U3145); 
assign P3_U4677 = ~(P3_U2435 & P3_U4661); 
assign P3_U4682 = ~(P3_U2433 & P3_U4661); 
assign P3_U4687 = ~(P3_U2431 & P3_U4661); 
assign P3_U4692 = ~(P3_U2429 & P3_U4661); 
assign P3_U4697 = ~(P3_U2427 & P3_U4661); 
assign P3_U4702 = ~(P3_U2425 & P3_U4661); 
assign P3_U4707 = ~(P3_U2423 & P3_U4661); 
assign P3_U4712 = ~(P3_U2421 & P3_U4661); 
assign P3_U4720 = ~P3_U3151; 
assign P3_U4721 = ~(P3_U2489 & P3_U3151); 
assign P3_U4729 = ~(P3_U4715 & P3_U2435); 
assign P3_U4734 = ~(P3_U4715 & P3_U2433); 
assign P3_U4739 = ~(P3_U4715 & P3_U2431); 
assign P3_U4744 = ~(P3_U4715 & P3_U2429); 
assign P3_U4749 = ~(P3_U4715 & P3_U2427); 
assign P3_U4754 = ~(P3_U4715 & P3_U2425); 
assign P3_U4759 = ~(P3_U4715 & P3_U2423); 
assign P3_U4764 = ~(P3_U4715 & P3_U2421); 
assign P3_U4772 = ~P3_U3159; 
assign P3_U4773 = ~(P3_U2489 & P3_U3159); 
assign P3_U4781 = ~(P3_U4767 & P3_U2435); 
assign P3_U4786 = ~(P3_U4767 & P3_U2433); 
assign P3_U4791 = ~(P3_U4767 & P3_U2431); 
assign P3_U4796 = ~(P3_U4767 & P3_U2429); 
assign P3_U4801 = ~(P3_U4767 & P3_U2427); 
assign P3_U4806 = ~(P3_U4767 & P3_U2425); 
assign P3_U4811 = ~(P3_U4767 & P3_U2423); 
assign P3_U4816 = ~(P3_U4767 & P3_U2421); 
assign P3_U4823 = ~P3_U3163; 
assign P3_U4824 = ~(P3_U2489 & P3_U3163); 
assign P3_U4832 = ~(P3_U4819 & P3_U2435); 
assign P3_U4837 = ~(P3_U4819 & P3_U2433); 
assign P3_U4842 = ~(P3_U4819 & P3_U2431); 
assign P3_U4847 = ~(P3_U4819 & P3_U2429); 
assign P3_U4852 = ~(P3_U4819 & P3_U2427); 
assign P3_U4857 = ~(P3_U4819 & P3_U2425); 
assign P3_U4862 = ~(P3_U4819 & P3_U2423); 
assign P3_U4867 = ~(P3_U4819 & P3_U2421); 
assign P3_U4875 = ~P3_U3167; 
assign P3_U4876 = ~(P3_U2489 & P3_U3167); 
assign P3_U4884 = ~(P3_U4870 & P3_U2435); 
assign P3_U4889 = ~(P3_U4870 & P3_U2433); 
assign P3_U4894 = ~(P3_U4870 & P3_U2431); 
assign P3_U4899 = ~(P3_U4870 & P3_U2429); 
assign P3_U4904 = ~(P3_U4870 & P3_U2427); 
assign P3_U4909 = ~(P3_U4870 & P3_U2425); 
assign P3_U4914 = ~(P3_U4870 & P3_U2423); 
assign P3_U4919 = ~(P3_U4870 & P3_U2421); 
assign P3_U4927 = ~P3_U3171; 
assign P3_U4928 = ~(P3_U2489 & P3_U3171); 
assign P3_U4936 = ~(P3_U4922 & P3_U2435); 
assign P3_U4941 = ~(P3_U4922 & P3_U2433); 
assign P3_U4946 = ~(P3_U4922 & P3_U2431); 
assign P3_U4951 = ~(P3_U4922 & P3_U2429); 
assign P3_U4956 = ~(P3_U4922 & P3_U2427); 
assign P3_U4961 = ~(P3_U4922 & P3_U2425); 
assign P3_U4966 = ~(P3_U4922 & P3_U2423); 
assign P3_U4971 = ~(P3_U4922 & P3_U2421); 
assign P3_U4979 = ~P3_U3175; 
assign P3_U4980 = ~(P3_U2489 & P3_U3175); 
assign P3_U4988 = ~(P3_U4974 & P3_U2435); 
assign P3_U4993 = ~(P3_U4974 & P3_U2433); 
assign P3_U4998 = ~(P3_U4974 & P3_U2431); 
assign P3_U5003 = ~(P3_U4974 & P3_U2429); 
assign P3_U5008 = ~(P3_U4974 & P3_U2427); 
assign P3_U5013 = ~(P3_U4974 & P3_U2425); 
assign P3_U5018 = ~(P3_U4974 & P3_U2423); 
assign P3_U5023 = ~(P3_U4974 & P3_U2421); 
assign P3_U5030 = ~P3_U3179; 
assign P3_U5031 = ~(P3_U2489 & P3_U3179); 
assign P3_U5039 = ~(P3_U5026 & P3_U2435); 
assign P3_U5044 = ~(P3_U5026 & P3_U2433); 
assign P3_U5049 = ~(P3_U5026 & P3_U2431); 
assign P3_U5054 = ~(P3_U5026 & P3_U2429); 
assign P3_U5059 = ~(P3_U5026 & P3_U2427); 
assign P3_U5064 = ~(P3_U5026 & P3_U2425); 
assign P3_U5069 = ~(P3_U5026 & P3_U2423); 
assign P3_U5074 = ~(P3_U5026 & P3_U2421); 
assign P3_U5077 = ~P3_U3183; 
assign P3_U5126 = ~P3_U3187; 
assign P3_U5178 = ~P3_U3191; 
assign P3_U5230 = ~P3_U3195; 
assign P3_U5234 = ~(P3_U3195 & P3_U5233); 
assign P3_U5280 = ~P3_U3197; 
assign P3_U5285 = ~(P3_U3197 & P3_U5284); 
assign P3_U5331 = ~P3_U3200; 
assign P3_U5336 = ~(P3_U3200 & P3_U5335); 
assign P3_U5382 = ~P3_U3203; 
assign P3_U5387 = ~(P3_U3203 & P3_U5386); 
assign P3_U5433 = ~P3_U3206; 
assign P3_U5437 = ~(P3_U3206 & P3_U5436); 
assign P3_U5488 = ~P3_U3255; 
assign P3_U5491 = ~P3_U3254; 
assign P3_U5492 = ~(P3_U3254 & P3_U2630); 
assign P3_U5494 = ~(P3_U4294 & P3_U3255); 
assign P3_U5585 = ~(P3_U3183 & P3_U5584); 
assign P3_U5656 = ~(P3_ADD_360_1242_U19 & P3_U2395); 
assign P3_U6402 = ~(P3_U2390 & P3_U6401); 
assign P3_U6757 = ~(P3_U3986 & P3_U3255); 
assign P3_U8000 = ~(P3_U5622 & P3_U3104); 
assign P3_U8001 = ~(P3_U4505 & P3_U5619); 
assign P2_U2446 = P2_R2088_U6 & P2_U4424; 
assign P2_U2687 = P2_ADD_402_1132_U25 & P2_U2355; 
assign P2_U2714 = ~(P2_U7871 & P2_U4408 & P2_STATE2_REG_0__SCAN_IN); 
assign P2_U3520 = ~P2_R2088_U6; 
assign P2_U3646 = ~(P2_U8346 & P2_U8345); 
assign P2_U3681 = ~(P2_U8418 & P2_U8417); 
assign P2_U5579 = ~(P2_U5578 & P2_U3265 & P2_R2088_U6); 
assign P2_U5668 = ~(P2_U8122 & P2_U8121 & P2_U3265 & P2_R2088_U6); 
assign P2_U6566 = ~(P2_R2088_U6 & P2_U4603); 
assign P1_U2742 = P1_U7492 & P1_U7491; 
assign P1_U3437 = ~(P1_U2447 & P1_U4498); 
assign P1_U3738 = P1_U3737 & P1_U2518; 
assign P1_U4002 = P1_U6749 & P1_U6748; 
assign P1_U6804 = ~(P1_R2182_U6 & P1_U6746); 
assign P3_ADD_526_U74 = ~(P3_ADD_526_U188 & P3_ADD_526_U187); 
assign P3_ADD_526_U75 = ~(P3_ADD_526_U190 & P3_ADD_526_U189); 
assign P3_ADD_526_U114 = ~P3_ADD_526_U34; 
assign P3_ADD_526_U136 = ~P3_ADD_526_U106; 
assign P3_ADD_526_U184 = ~(P3_ADD_526_U34 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_526_U185 = ~(P3_ADD_526_U106 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_552_U74 = ~(P3_ADD_552_U188 & P3_ADD_552_U187); 
assign P3_ADD_552_U75 = ~(P3_ADD_552_U190 & P3_ADD_552_U189); 
assign P3_ADD_552_U114 = ~P3_ADD_552_U34; 
assign P3_ADD_552_U136 = ~P3_ADD_552_U106; 
assign P3_ADD_552_U184 = ~(P3_ADD_552_U34 & P3_EBX_REG_19__SCAN_IN); 
assign P3_ADD_552_U185 = ~(P3_ADD_552_U106 & P3_EBX_REG_18__SCAN_IN); 
assign P3_ADD_546_U74 = ~(P3_ADD_546_U188 & P3_ADD_546_U187); 
assign P3_ADD_546_U75 = ~(P3_ADD_546_U190 & P3_ADD_546_U189); 
assign P3_ADD_546_U114 = ~P3_ADD_546_U34; 
assign P3_ADD_546_U136 = ~P3_ADD_546_U106; 
assign P3_ADD_546_U184 = ~(P3_ADD_546_U34 & P3_EAX_REG_19__SCAN_IN); 
assign P3_ADD_546_U185 = ~(P3_ADD_546_U106 & P3_EAX_REG_18__SCAN_IN); 
assign P3_ADD_391_1180_U12 = ~(P3_U2616 & P3_ADD_391_1180_U30); 
assign P3_ADD_391_1180_U44 = ~(P3_ADD_391_1180_U30 & P3_ADD_391_1180_U11); 
assign P3_ADD_476_U91 = ~(P3_ADD_476_U182 & P3_ADD_476_U181); 
assign P3_ADD_476_U102 = ~P3_ADD_476_U22; 
assign P3_ADD_476_U179 = ~(P3_ADD_476_U22 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_531_U65 = ~(P3_ADD_531_U129 & P3_ADD_531_U128); 
assign P3_ADD_531_U106 = ~P3_ADD_531_U23; 
assign P3_ADD_531_U188 = ~(P3_ADD_531_U23 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_SUB_320_U125 = ~(P3_SUB_320_U86 & P3_SUB_320_U52); 
assign P3_SUB_320_U129 = ~(P3_SUB_320_U86 & P3_SUB_320_U52); 
assign P3_ADD_318_U91 = ~(P3_ADD_318_U182 & P3_ADD_318_U181); 
assign P3_ADD_318_U102 = ~P3_ADD_318_U22; 
assign P3_ADD_318_U179 = ~(P3_ADD_318_U22 & P3_PHYADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_315_U87 = ~(P3_ADD_315_U174 & P3_ADD_315_U173); 
assign P3_ADD_315_U99 = ~P3_ADD_315_U22; 
assign P3_ADD_315_U171 = ~(P3_ADD_315_U22 & P3_PHYADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_360_1242_U20 = ~P3_ADD_360_U19; 
assign P3_ADD_360_1242_U40 = ~(P3_ADD_360_1242_U131 & P3_ADD_360_1242_U130); 
assign P3_ADD_360_1242_U115 = P3_ADD_360_1242_U226 & P3_ADD_360_1242_U225; 
assign P3_ADD_360_1242_U123 = P3_ADD_360_U19 | P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_360_1242_U125 = ~(P3_ADD_360_U19 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_360_1242_U224 = ~(P3_ADD_360_U19 & P3_ADD_360_1242_U21); 
assign P3_ADD_360_1242_U236 = ~(P3_ADD_360_1242_U117 & P3_ADD_360_1242_U118); 
assign P3_ADD_360_1242_U237 = ~(P3_ADD_360_1242_U128 & P3_ADD_360_1242_U235); 
assign P3_ADD_467_U91 = ~(P3_ADD_467_U182 & P3_ADD_467_U181); 
assign P3_ADD_467_U102 = ~P3_ADD_467_U22; 
assign P3_ADD_467_U179 = ~(P3_ADD_467_U22 & P3_REIP_REG_11__SCAN_IN); 
assign P3_ADD_430_U91 = ~(P3_ADD_430_U182 & P3_ADD_430_U181); 
assign P3_ADD_430_U102 = ~P3_ADD_430_U22; 
assign P3_ADD_430_U179 = ~(P3_ADD_430_U22 & P3_REIP_REG_11__SCAN_IN); 
assign P3_ADD_380_U65 = ~(P3_ADD_380_U129 & P3_ADD_380_U128); 
assign P3_ADD_380_U106 = ~P3_ADD_380_U23; 
assign P3_ADD_380_U188 = ~(P3_ADD_380_U23 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_344_U65 = ~(P3_ADD_344_U129 & P3_ADD_344_U128); 
assign P3_ADD_344_U106 = ~P3_ADD_344_U23; 
assign P3_ADD_344_U188 = ~(P3_ADD_344_U23 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_339_U91 = ~(P3_ADD_339_U182 & P3_ADD_339_U181); 
assign P3_ADD_339_U102 = ~P3_ADD_339_U22; 
assign P3_ADD_339_U179 = ~(P3_ADD_339_U22 & P3_PHYADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_360_U13 = ~(P3_U2626 & P3_ADD_360_U26); 
assign P3_ADD_360_U34 = ~(P3_ADD_360_U26 & P3_ADD_360_U12); 
assign P3_ADD_541_U91 = ~(P3_ADD_541_U182 & P3_ADD_541_U181); 
assign P3_ADD_541_U102 = ~P3_ADD_541_U22; 
assign P3_ADD_541_U179 = ~(P3_ADD_541_U22 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_SUB_357_1258_U24 = ~P3_ADD_357_U8; 
assign P3_SUB_357_1258_U39 = ~P3_ADD_357_U6; 
assign P3_SUB_357_1258_U94 = P3_SUB_357_1258_U163 & P3_SUB_357_1258_U164 & P3_SUB_357_1258_U160; 
assign P3_SUB_357_1258_U155 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_SUB_357_1258_U156 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_SUB_357_1258_U157 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_SUB_357_1258_U165 = ~P3_SUB_357_1258_U127; 
assign P3_SUB_357_1258_U168 = ~(P3_SUB_357_1258_U95 & P3_SUB_357_1258_U160); 
assign P3_SUB_357_1258_U170 = P3_ADD_357_U8 | P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_SUB_357_1258_U178 = P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P3_SUB_357_1258_U179 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_SUB_357_1258_U180 = ~(P3_SUB_357_1258_U97 & P3_SUB_357_1258_U166); 
assign P3_SUB_357_1258_U183 = ~(P3_SUB_357_1258_U127 & P3_SUB_357_1258_U164); 
assign P3_SUB_357_1258_U186 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_SUB_357_1258_U187 = P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P3_SUB_357_1258_U188 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_SUB_357_1258_U189 = P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P3_SUB_357_1258_U190 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_SUB_357_1258_U192 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_SUB_357_1258_U193 = P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P3_SUB_357_1258_U195 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_SUB_357_1258_U197 = P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P3_SUB_357_1258_U199 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_SUB_357_1258_U204 = P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P3_SUB_357_1258_U205 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_SUB_357_1258_U206 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_SUB_357_1258_U210 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_SUB_357_1258_U211 = P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P3_SUB_357_1258_U212 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_SUB_357_1258_U213 = P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P3_SUB_357_1258_U214 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_SUB_357_1258_U215 = P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P3_SUB_357_1258_U216 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_SUB_357_1258_U219 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_SUB_357_1258_U228 = P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_SUB_357_1258_U232 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_SUB_357_1258_U234 = P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P3_SUB_357_1258_U245 = P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P3_SUB_357_1258_U250 = P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_SUB_357_1258_U254 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_SUB_357_1258_U256 = P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P3_SUB_357_1258_U257 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_SUB_357_1258_U259 = ~(P3_SUB_357_1258_U162 & P3_SUB_357_1258_U160); 
assign P3_SUB_357_1258_U266 = ~(P3_ADD_357_U8 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_SUB_357_1258_U268 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_SUB_357_1258_U269 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_SUB_357_1258_U273 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_SUB_357_1258_U275 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_SUB_357_1258_U307 = ~(P3_SUB_357_1258_U158 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_SUB_357_1258_U308 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U41); 
assign P3_SUB_357_1258_U313 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U40); 
assign P3_SUB_357_1258_U315 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U40); 
assign P3_SUB_357_1258_U335 = ~(P3_ADD_357_U8 & P3_SUB_357_1258_U25); 
assign P3_SUB_357_1258_U337 = ~(P3_ADD_357_U8 & P3_SUB_357_1258_U25); 
assign P3_SUB_357_1258_U341 = ~(P3_SUB_357_1258_U26 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_SUB_357_1258_U348 = ~(P3_SUB_357_1258_U347 & P3_SUB_357_1258_U346); 
assign P3_SUB_357_1258_U353 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_SUB_357_1258_U355 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U60); 
assign P3_SUB_357_1258_U357 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U60); 
assign P3_SUB_357_1258_U364 = ~(P3_SUB_357_1258_U363 & P3_SUB_357_1258_U362); 
assign P3_SUB_357_1258_U365 = ~(P3_SUB_357_1258_U261 & P3_SUB_357_1258_U127); 
assign P3_SUB_357_1258_U367 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U59); 
assign P3_SUB_357_1258_U369 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U59); 
assign P3_SUB_357_1258_U376 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_SUB_357_1258_U379 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U58); 
assign P3_SUB_357_1258_U381 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U58); 
assign P3_SUB_357_1258_U386 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U43); 
assign P3_SUB_357_1258_U388 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U42); 
assign P3_SUB_357_1258_U393 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U44); 
assign P3_SUB_357_1258_U395 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U44); 
assign P3_SUB_357_1258_U400 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U45); 
assign P3_SUB_357_1258_U402 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U45); 
assign P3_SUB_357_1258_U407 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U46); 
assign P3_SUB_357_1258_U409 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U46); 
assign P3_SUB_357_1258_U414 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U48); 
assign P3_SUB_357_1258_U416 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U48); 
assign P3_SUB_357_1258_U426 = ~(P3_SUB_357_1258_U424 & P3_SUB_357_1258_U31); 
assign P3_SUB_357_1258_U428 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U47); 
assign P3_SUB_357_1258_U433 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U49); 
assign P3_SUB_357_1258_U435 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U49); 
assign P3_SUB_357_1258_U441 = ~(P3_ADD_357_U6 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_SUB_357_1258_U444 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U56); 
assign P3_SUB_357_1258_U446 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U56); 
assign P3_SUB_357_1258_U451 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U55); 
assign P3_SUB_357_1258_U453 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U55); 
assign P3_SUB_357_1258_U458 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U54); 
assign P3_SUB_357_1258_U460 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U54); 
assign P3_SUB_357_1258_U465 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U51); 
assign P3_SUB_357_1258_U467 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U50); 
assign P3_SUB_357_1258_U472 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U52); 
assign P3_SUB_357_1258_U474 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U52); 
assign P3_SUB_357_1258_U479 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U53); 
assign P3_ADD_515_U91 = ~(P3_ADD_515_U182 & P3_ADD_515_U181); 
assign P3_ADD_515_U102 = ~P3_ADD_515_U22; 
assign P3_ADD_515_U179 = ~(P3_ADD_515_U22 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_394_U91 = ~(P3_ADD_394_U186 & P3_ADD_394_U185); 
assign P3_ADD_394_U105 = ~P3_ADD_394_U22; 
assign P3_ADD_394_U183 = ~(P3_ADD_394_U22 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_SUB_414_U76 = P3_SUB_414_U153 & P3_SUB_414_U152; 
assign P3_SUB_414_U97 = ~P3_SUB_414_U32; 
assign P3_SUB_414_U118 = ~(P3_SUB_414_U117 & P3_EBX_REG_18__SCAN_IN); 
assign P3_SUB_414_U150 = ~(P3_SUB_414_U32 & P3_EBX_REG_19__SCAN_IN); 
assign P3_ADD_441_U91 = ~(P3_ADD_441_U182 & P3_ADD_441_U181); 
assign P3_ADD_441_U102 = ~P3_ADD_441_U22; 
assign P3_ADD_441_U179 = ~(P3_ADD_441_U22 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_349_U65 = ~(P3_ADD_349_U129 & P3_ADD_349_U128); 
assign P3_ADD_349_U106 = ~P3_ADD_349_U23; 
assign P3_ADD_349_U188 = ~(P3_ADD_349_U23 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_405_U91 = ~(P3_ADD_405_U186 & P3_ADD_405_U185); 
assign P3_ADD_405_U105 = ~P3_ADD_405_U22; 
assign P3_ADD_405_U183 = ~(P3_ADD_405_U22 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_553_U65 = ~(P3_ADD_553_U129 & P3_ADD_553_U128); 
assign P3_ADD_553_U106 = ~P3_ADD_553_U23; 
assign P3_ADD_553_U188 = ~(P3_ADD_553_U23 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_558_U65 = ~(P3_ADD_558_U129 & P3_ADD_558_U128); 
assign P3_ADD_558_U106 = ~P3_ADD_558_U23; 
assign P3_ADD_558_U188 = ~(P3_ADD_558_U23 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_385_U65 = ~(P3_ADD_385_U129 & P3_ADD_385_U128); 
assign P3_ADD_385_U106 = ~P3_ADD_385_U23; 
assign P3_ADD_385_U188 = ~(P3_ADD_385_U23 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_357_U17 = P3_ADD_357_U31 & P3_ADD_357_U30; 
assign P3_ADD_357_U25 = ~(P3_SUB_357_U8 & P3_ADD_357_U24); 
assign P3_ADD_547_U65 = ~(P3_ADD_547_U129 & P3_ADD_547_U128); 
assign P3_ADD_547_U106 = ~P3_ADD_547_U23; 
assign P3_ADD_547_U188 = ~(P3_ADD_547_U23 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_371_1212_U20 = ~(P3_ADD_371_1212_U255 & P3_ADD_371_1212_U254 & P3_ADD_371_1212_U203); 
assign P3_ADD_371_1212_U21 = ~P3_ADD_371_U20; 
assign P3_ADD_371_1212_U24 = ~(P3_ADD_371_U20 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_371_1212_U44 = ~(P3_ADD_371_1212_U77 & P3_ADD_371_1212_U123); 
assign P3_ADD_371_1212_U119 = ~(P3_ADD_371_1212_U202 & P3_ADD_371_1212_U201); 
assign P3_ADD_371_1212_U127 = ~(P3_ADD_371_1212_U30 & P3_ADD_371_1212_U29); 
assign P3_ADD_371_1212_U133 = P3_ADD_371_U20 | P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_371_1212_U150 = P3_ADD_371_U20 | P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_371_1212_U156 = P3_ADD_371_U20 | P3_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P3_ADD_371_1212_U230 = ~(P3_ADD_371_U20 & P3_ADD_371_1212_U22); 
assign P3_ADD_371_1212_U234 = ~(P3_ADD_371_1212_U30 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_371_U13 = ~(P3_U2626 & P3_ADD_371_U29); 
assign P3_ADD_371_U38 = ~(P3_ADD_371_U29 & P3_ADD_371_U12); 
assign P3_ADD_494_U91 = ~(P3_ADD_494_U182 & P3_ADD_494_U181); 
assign P3_ADD_494_U102 = ~P3_ADD_494_U22; 
assign P3_ADD_494_U179 = ~(P3_ADD_494_U22 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_536_U91 = ~(P3_ADD_536_U182 & P3_ADD_536_U181); 
assign P3_ADD_536_U102 = ~P3_ADD_536_U22; 
assign P3_ADD_536_U179 = ~(P3_ADD_536_U22 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_402_1132_U12 = ~(P3_U2616 & P3_ADD_402_1132_U30); 
assign P3_ADD_402_1132_U44 = ~(P3_ADD_402_1132_U30 & P3_ADD_402_1132_U11); 
assign P2_R2099_U6 = ~P2_U2747; 
assign P2_R2099_U8 = ~P2_U2750; 
assign P2_R2099_U10 = ~P2_U2749; 
assign P2_R2099_U12 = ~P2_U2748; 
assign P2_R2099_U105 = ~(P2_U2751 & P2_U2747); 
assign P2_R2099_U106 = ~(P2_U2746 & P2_U2747 & P2_U2751); 
assign P2_R2099_U112 = P2_U2749 | P2_U2745; 
assign P2_R2099_U114 = ~(P2_U2745 & P2_U2749); 
assign P2_R2099_U116 = P2_U2748 | P2_U2744; 
assign P2_R2099_U118 = ~(P2_U2744 & P2_U2748); 
assign P2_R2099_U162 = ~(P2_U2748 & P2_R2099_U13); 
assign P2_R2099_U164 = ~(P2_U2748 & P2_R2099_U13); 
assign P2_R2099_U173 = ~(P2_U2749 & P2_R2099_U11); 
assign P2_R2099_U175 = ~(P2_U2749 & P2_R2099_U11); 
assign P2_R2099_U225 = ~(P2_U2747 & P2_R2099_U7); 
assign P2_ADD_402_1132_U12 = ~(P2_U2594 & P2_ADD_402_1132_U30); 
assign P2_ADD_402_1132_U42 = ~(P2_ADD_402_1132_U30 & P2_ADD_402_1132_U11); 
assign P2_R2182_U259 = ~(P2_U2664 & P2_R2182_U54); 
assign P2_R2182_U261 = ~(P2_U2664 & P2_R2182_U54); 
assign P2_R2182_U266 = ~(P2_U2665 & P2_R2182_U52); 
assign P2_R2182_U268 = ~(P2_U2665 & P2_R2182_U52); 
assign P2_R2027_U65 = ~(P2_R2027_U129 & P2_R2027_U128); 
assign P2_R2027_U106 = ~P2_R2027_U23; 
assign P2_R2027_U188 = ~(P2_R2027_U23 & P2_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P2_R2337_U89 = ~(P2_R2337_U180 & P2_R2337_U179); 
assign P2_R2337_U103 = ~P2_R2337_U23; 
assign P2_R2337_U177 = ~(P2_R2337_U23 & P2_PHYADDRPOINTER_REG_12__SCAN_IN); 
assign P2_R2219_U49 = ~(P2_R2219_U48 & P2_R2219_U81); 
assign P2_R2219_U71 = ~(P2_R2219_U6 & P2_R2219_U44); 
assign P2_R2219_U73 = ~P2_R2219_U19; 
assign P2_R2219_U74 = ~(P2_R2219_U31 & P2_R2219_U44); 
assign P2_R2219_U79 = ~P2_R2219_U44; 
assign P2_R2219_U111 = ~(P2_R2219_U37 & P2_R2219_U44); 
assign P2_R2219_U115 = ~(P2_R2219_U46 & P2_R2219_U114); 
assign P2_R2096_U119 = ~P2_R2096_U111; 
assign P2_R2096_U121 = ~(P2_R2096_U120 & P2_R2096_U111); 
assign P2_R2096_U170 = ~(P2_R2096_U241 & P2_R2096_U55); 
assign P2_R2096_U217 = ~(P2_R2096_U110 & P2_R2096_U111); 
assign P2_R1957_U125 = ~(P2_R1957_U86 & P2_R1957_U52); 
assign P2_R1957_U129 = ~(P2_R1957_U86 & P2_R1957_U52); 
assign P2_ADD_394_U83 = ~(P2_ADD_394_U168 & P2_ADD_394_U167); 
assign P2_ADD_394_U105 = ~P2_ADD_394_U22; 
assign P2_ADD_394_U147 = ~(P2_ADD_394_U22 & P2_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P1_R2027_U74 = ~(P1_R2027_U188 & P1_R2027_U187); 
assign P1_R2027_U75 = ~(P1_R2027_U190 & P1_R2027_U189); 
assign P1_R2027_U114 = ~P1_R2027_U34; 
assign P1_R2027_U136 = ~P1_R2027_U106; 
assign P1_R2027_U184 = ~(P1_R2027_U34 & P1_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P1_R2027_U185 = ~(P1_R2027_U106 & P1_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P1_R2182_U11 = ~P1_U2741; 
assign P1_R2182_U19 = ~(P1_R2182_U36 & P1_R2182_U49); 
assign P1_R2182_U44 = ~(P1_R2182_U49 & P1_U2738); 
assign P1_R2182_U50 = ~P1_R2182_U9; 
assign P1_R2182_U51 = P1_U2743 | P1_U2731; 
assign P1_R2182_U52 = ~(P1_U2731 & P1_U2743); 
assign P1_R2182_U62 = ~(P1_U2731 & P1_U2743); 
assign P1_R2182_U81 = ~(P1_R2182_U49 & P1_R2182_U15); 
assign P1_R2182_U85 = ~(P1_U3246 & P1_R2182_U7); 
assign P1_R2182_U86 = ~(P1_U2744 & P1_R2182_U8); 
assign P1_R2144_U81 = ~(P1_R2144_U165 & P1_R2144_U164 & P1_R2144_U22); 
assign P1_R2144_U104 = ~(P1_R2144_U167 & P1_R2144_U166 & P1_R2144_U17); 
assign P1_R2144_U105 = ~(P1_R2144_U175 & P1_R2144_U174 & P1_R2144_U20); 
assign P1_R2144_U106 = ~(P1_R2144_U201 & P1_R2144_U200 & P1_R2144_U18); 
assign P1_R2144_U170 = ~(P1_R2144_U169 & P1_R2144_U168); 
assign P1_R2144_U173 = ~(P1_R2144_U172 & P1_R2144_U171); 
assign P1_R2144_U178 = ~(P1_R2144_U177 & P1_R2144_U176); 
assign P1_R2144_U181 = ~(P1_R2144_U180 & P1_R2144_U179); 
assign P1_R2358_U152 = ~P1_U2617; 
assign P1_R2358_U421 = ~(P1_R2358_U420 & P1_R2358_U419); 
assign P1_R2358_U445 = ~(P1_U2617 & P1_R2358_U23); 
assign P1_R2358_U447 = ~(P1_U2617 & P1_R2358_U23); 
assign P1_R2099_U137 = ~(P1_R2099_U152 & P1_R2099_U151); 
assign P1_R2099_U323 = ~(P1_R2099_U139 & P1_R2099_U140); 
assign P1_R2099_U324 = ~(P1_R2099_U149 & P1_R2099_U322); 
assign P1_R2167_U20 = P1_R2167_U35 & P1_R2167_U36; 
assign P1_R2167_U21 = P1_R2167_U38 & P1_R2167_U39; 
assign P1_R2167_U34 = ~(P1_R2167_U19 & P1_R2167_U31); 
assign P1_R2337_U91 = ~(P1_R2337_U182 & P1_R2337_U181); 
assign P1_R2337_U102 = ~P1_R2337_U22; 
assign P1_R2337_U179 = ~(P1_R2337_U22 & P1_PHYADDRPOINTER_REG_11__SCAN_IN); 
assign P1_R2096_U91 = ~(P1_R2096_U182 & P1_R2096_U181); 
assign P1_R2096_U102 = ~P1_R2096_U22; 
assign P1_R2096_U179 = ~(P1_R2096_U22 & P1_REIP_REG_11__SCAN_IN); 
assign P1_ADD_371_U19 = ~(P1_ADD_371_U38 & P1_ADD_371_U37); 
assign P1_ADD_371_U30 = ~P1_ADD_371_U14; 
assign P1_ADD_371_U33 = ~(P1_U3233 & P1_ADD_371_U14); 
assign P1_ADD_405_U83 = ~(P1_ADD_405_U168 & P1_ADD_405_U167); 
assign P1_ADD_405_U105 = ~P1_ADD_405_U22; 
assign P1_ADD_405_U147 = ~(P1_ADD_405_U22 & P1_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P1_ADD_515_U83 = ~(P1_ADD_515_U166 & P1_ADD_515_U165); 
assign P1_ADD_515_U102 = ~P1_ADD_515_U22; 
assign P1_ADD_515_U145 = ~(P1_ADD_515_U22 & P1_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_U2516 = P3_U5493 & P3_U5492; 
assign P3_U3249 = ~(P3_U6403 & P3_U6402); 
assign P3_U3251 = ~(P3_U6758 & P3_U6757); 
assign P3_U3262 = ~(P3_U2462 & P3_U3108 & P3_U4282); 
assign P3_U3371 = P3_U3370 & P3_U4677; 
assign P3_U3373 = P3_U3372 & P3_U4682; 
assign P3_U3375 = P3_U3374 & P3_U4687; 
assign P3_U3377 = P3_U3376 & P3_U4692; 
assign P3_U3379 = P3_U3378 & P3_U4697; 
assign P3_U3381 = P3_U3380 & P3_U4702; 
assign P3_U3383 = P3_U3382 & P3_U4707; 
assign P3_U3385 = P3_U3384 & P3_U4712; 
assign P3_U3389 = P3_U3388 & P3_U4729; 
assign P3_U3391 = P3_U3390 & P3_U4734; 
assign P3_U3393 = P3_U3392 & P3_U4739; 
assign P3_U3395 = P3_U3394 & P3_U4744; 
assign P3_U3397 = P3_U3396 & P3_U4749; 
assign P3_U3399 = P3_U3398 & P3_U4754; 
assign P3_U3401 = P3_U3400 & P3_U4759; 
assign P3_U3403 = P3_U3402 & P3_U4764; 
assign P3_U3407 = P3_U3406 & P3_U4781; 
assign P3_U3409 = P3_U3408 & P3_U4786; 
assign P3_U3411 = P3_U3410 & P3_U4791; 
assign P3_U3413 = P3_U3412 & P3_U4796; 
assign P3_U3415 = P3_U3414 & P3_U4801; 
assign P3_U3417 = P3_U3416 & P3_U4806; 
assign P3_U3419 = P3_U3418 & P3_U4811; 
assign P3_U3421 = P3_U3420 & P3_U4816; 
assign P3_U3425 = P3_U3424 & P3_U4832; 
assign P3_U3427 = P3_U3426 & P3_U4837; 
assign P3_U3429 = P3_U3428 & P3_U4842; 
assign P3_U3431 = P3_U3430 & P3_U4847; 
assign P3_U3433 = P3_U3432 & P3_U4852; 
assign P3_U3435 = P3_U3434 & P3_U4857; 
assign P3_U3437 = P3_U3436 & P3_U4862; 
assign P3_U3439 = P3_U3438 & P3_U4867; 
assign P3_U3442 = P3_U3441 & P3_U4884; 
assign P3_U3444 = P3_U3443 & P3_U4889; 
assign P3_U3446 = P3_U3445 & P3_U4894; 
assign P3_U3448 = P3_U3447 & P3_U4899; 
assign P3_U3450 = P3_U3449 & P3_U4904; 
assign P3_U3452 = P3_U3451 & P3_U4909; 
assign P3_U3454 = P3_U3453 & P3_U4914; 
assign P3_U3456 = P3_U3455 & P3_U4919; 
assign P3_U3460 = P3_U3459 & P3_U4936; 
assign P3_U3462 = P3_U3461 & P3_U4941; 
assign P3_U3464 = P3_U3463 & P3_U4946; 
assign P3_U3466 = P3_U3465 & P3_U4951; 
assign P3_U3468 = P3_U3467 & P3_U4956; 
assign P3_U3470 = P3_U3469 & P3_U4961; 
assign P3_U3472 = P3_U3471 & P3_U4966; 
assign P3_U3474 = P3_U3473 & P3_U4971; 
assign P3_U3478 = P3_U3477 & P3_U4988; 
assign P3_U3480 = P3_U3479 & P3_U4993; 
assign P3_U3482 = P3_U3481 & P3_U4998; 
assign P3_U3484 = P3_U3483 & P3_U5003; 
assign P3_U3486 = P3_U3485 & P3_U5008; 
assign P3_U3488 = P3_U3487 & P3_U5013; 
assign P3_U3490 = P3_U3489 & P3_U5018; 
assign P3_U3492 = P3_U3491 & P3_U5023; 
assign P3_U3495 = P3_U3494 & P3_U5039; 
assign P3_U3497 = P3_U3496 & P3_U5044; 
assign P3_U3499 = P3_U3498 & P3_U5049; 
assign P3_U3501 = P3_U3500 & P3_U5054; 
assign P3_U3503 = P3_U3502 & P3_U5059; 
assign P3_U3505 = P3_U3504 & P3_U5064; 
assign P3_U3507 = P3_U3506 & P3_U5069; 
assign P3_U3509 = P3_U3508 & P3_U5074; 
assign P3_U3657 = P3_U3656 & P3_U5494; 
assign P3_U4309 = ~P3_U3253; 
assign P3_U4311 = ~P3_U3250; 
assign P3_U4617 = ~(P3_U3358 & P3_U3357); 
assign P3_U4620 = ~(P3_U4280 & P3_U4619); 
assign P3_U4670 = ~(P3_U4664 & P3_U4669); 
assign P3_U4673 = ~(P3_U4668 & P3_U4322); 
assign P3_U4722 = ~(P3_U4718 & P3_U4721); 
assign P3_U4725 = ~(P3_U4720 & P3_U4322); 
assign P3_U4774 = ~(P3_U4770 & P3_U4773); 
assign P3_U4777 = ~(P3_U4772 & P3_U4322); 
assign P3_U4825 = ~(P3_U4824 & P3_U3070); 
assign P3_U4828 = ~(P3_U4823 & P3_U4322); 
assign P3_U4877 = ~(P3_U4873 & P3_U4876); 
assign P3_U4880 = ~(P3_U4875 & P3_U4322); 
assign P3_U4929 = ~(P3_U4925 & P3_U4928); 
assign P3_U4932 = ~(P3_U4927 & P3_U4322); 
assign P3_U4981 = ~(P3_U4977 & P3_U4980); 
assign P3_U4984 = ~(P3_U4979 & P3_U4322); 
assign P3_U5032 = ~(P3_U5031 & P3_U3071); 
assign P3_U5035 = ~(P3_U5030 & P3_U4322); 
assign P3_U5079 = ~P3_U3184; 
assign P3_U5080 = ~(P3_U2489 & P3_U3184); 
assign P3_U5088 = ~(P3_U5077 & P3_U2435); 
assign P3_U5093 = ~(P3_U5077 & P3_U2433); 
assign P3_U5098 = ~(P3_U5077 & P3_U2431); 
assign P3_U5103 = ~(P3_U5077 & P3_U2429); 
assign P3_U5108 = ~(P3_U5077 & P3_U2427); 
assign P3_U5113 = ~(P3_U5077 & P3_U2425); 
assign P3_U5118 = ~(P3_U5077 & P3_U2423); 
assign P3_U5123 = ~(P3_U5077 & P3_U2421); 
assign P3_U5131 = ~P3_U3188; 
assign P3_U5132 = ~(P3_U2489 & P3_U3188); 
assign P3_U5140 = ~(P3_U5126 & P3_U2435); 
assign P3_U5145 = ~(P3_U5126 & P3_U2433); 
assign P3_U5150 = ~(P3_U5126 & P3_U2431); 
assign P3_U5155 = ~(P3_U5126 & P3_U2429); 
assign P3_U5160 = ~(P3_U5126 & P3_U2427); 
assign P3_U5165 = ~(P3_U5126 & P3_U2425); 
assign P3_U5170 = ~(P3_U5126 & P3_U2423); 
assign P3_U5175 = ~(P3_U5126 & P3_U2421); 
assign P3_U5183 = ~P3_U3192; 
assign P3_U5184 = ~(P3_U2489 & P3_U3192); 
assign P3_U5192 = ~(P3_U5178 & P3_U2435); 
assign P3_U5197 = ~(P3_U5178 & P3_U2433); 
assign P3_U5202 = ~(P3_U5178 & P3_U2431); 
assign P3_U5207 = ~(P3_U5178 & P3_U2429); 
assign P3_U5212 = ~(P3_U5178 & P3_U2427); 
assign P3_U5217 = ~(P3_U5178 & P3_U2425); 
assign P3_U5222 = ~(P3_U5178 & P3_U2423); 
assign P3_U5227 = ~(P3_U5178 & P3_U2421); 
assign P3_U5235 = ~(P3_U2489 & P3_U5234); 
assign P3_U5242 = ~(P3_U5230 & P3_U2435); 
assign P3_U5247 = ~(P3_U5230 & P3_U2433); 
assign P3_U5252 = ~(P3_U5230 & P3_U2431); 
assign P3_U5257 = ~(P3_U5230 & P3_U2429); 
assign P3_U5262 = ~(P3_U5230 & P3_U2427); 
assign P3_U5267 = ~(P3_U5230 & P3_U2425); 
assign P3_U5272 = ~(P3_U5230 & P3_U2423); 
assign P3_U5277 = ~(P3_U5230 & P3_U2421); 
assign P3_U5286 = ~(P3_U2489 & P3_U5285); 
assign P3_U5293 = ~(P3_U5280 & P3_U2435); 
assign P3_U5298 = ~(P3_U5280 & P3_U2433); 
assign P3_U5303 = ~(P3_U5280 & P3_U2431); 
assign P3_U5308 = ~(P3_U5280 & P3_U2429); 
assign P3_U5313 = ~(P3_U5280 & P3_U2427); 
assign P3_U5318 = ~(P3_U5280 & P3_U2425); 
assign P3_U5323 = ~(P3_U5280 & P3_U2423); 
assign P3_U5328 = ~(P3_U5280 & P3_U2421); 
assign P3_U5337 = ~(P3_U2489 & P3_U5336); 
assign P3_U5344 = ~(P3_U5331 & P3_U2435); 
assign P3_U5349 = ~(P3_U5331 & P3_U2433); 
assign P3_U5354 = ~(P3_U5331 & P3_U2431); 
assign P3_U5359 = ~(P3_U5331 & P3_U2429); 
assign P3_U5364 = ~(P3_U5331 & P3_U2427); 
assign P3_U5369 = ~(P3_U5331 & P3_U2425); 
assign P3_U5374 = ~(P3_U5331 & P3_U2423); 
assign P3_U5379 = ~(P3_U5331 & P3_U2421); 
assign P3_U5388 = ~(P3_U2489 & P3_U5387); 
assign P3_U5395 = ~(P3_U5382 & P3_U2435); 
assign P3_U5400 = ~(P3_U5382 & P3_U2433); 
assign P3_U5405 = ~(P3_U5382 & P3_U2431); 
assign P3_U5410 = ~(P3_U5382 & P3_U2429); 
assign P3_U5415 = ~(P3_U5382 & P3_U2427); 
assign P3_U5420 = ~(P3_U5382 & P3_U2425); 
assign P3_U5425 = ~(P3_U5382 & P3_U2423); 
assign P3_U5430 = ~(P3_U5382 & P3_U2421); 
assign P3_U5438 = ~(P3_U2489 & P3_U5437); 
assign P3_U5445 = ~(P3_U5433 & P3_U2435); 
assign P3_U5450 = ~(P3_U5433 & P3_U2433); 
assign P3_U5455 = ~(P3_U5433 & P3_U2431); 
assign P3_U5460 = ~(P3_U5433 & P3_U2429); 
assign P3_U5465 = ~(P3_U5433 & P3_U2427); 
assign P3_U5470 = ~(P3_U5433 & P3_U2425); 
assign P3_U5475 = ~(P3_U5433 & P3_U2423); 
assign P3_U5480 = ~(P3_U5433 & P3_U2421); 
assign P3_U5522 = ~P3_U3220; 
assign P3_U5538 = ~(P3_U3670 & P3_U3220); 
assign P3_U5586 = ~(P3_U4322 & P3_U5585); 
assign P3_U5624 = ~(P3_U8001 & P3_U8000 & P3_U5623); 
assign P3_U5634 = ~(P3_ADD_558_U5 & P3_U3220); 
assign P3_U5637 = ~(P3_U4300 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_U5638 = ~(P3_U4301 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_U5658 = ~(P3_ADD_558_U85 & P3_U3220); 
assign P3_U5661 = ~(P3_ADD_541_U4 & P3_U4300); 
assign P3_U5662 = ~(P3_ADD_536_U4 & P3_U4301); 
assign P3_U5675 = ~(P3_ADD_371_1212_U20 & P3_U2360); 
assign P3_U5682 = ~(P3_ADD_558_U74 & P3_U3220); 
assign P3_U5685 = ~(P3_ADD_541_U71 & P3_U4300); 
assign P3_U5686 = ~(P3_ADD_536_U71 & P3_U4301); 
assign P3_U5706 = ~(P3_ADD_558_U71 & P3_U3220); 
assign P3_U5709 = ~(P3_ADD_541_U68 & P3_U4300); 
assign P3_U5710 = ~(P3_ADD_536_U68 & P3_U4301); 
assign P3_U5730 = ~(P3_ADD_558_U70 & P3_U3220); 
assign P3_U5733 = ~(P3_ADD_541_U67 & P3_U4300); 
assign P3_U5734 = ~(P3_ADD_536_U67 & P3_U4301); 
assign P3_U5754 = ~(P3_ADD_558_U69 & P3_U3220); 
assign P3_U5757 = ~(P3_ADD_541_U66 & P3_U4300); 
assign P3_U5758 = ~(P3_ADD_536_U66 & P3_U4301); 
assign P3_U5778 = ~(P3_ADD_558_U68 & P3_U3220); 
assign P3_U5781 = ~(P3_ADD_541_U65 & P3_U4300); 
assign P3_U5782 = ~(P3_ADD_536_U65 & P3_U4301); 
assign P3_U5802 = ~(P3_ADD_558_U67 & P3_U3220); 
assign P3_U5805 = ~(P3_ADD_541_U64 & P3_U4300); 
assign P3_U5806 = ~(P3_ADD_536_U64 & P3_U4301); 
assign P3_U5826 = ~(P3_ADD_558_U66 & P3_U3220); 
assign P3_U5829 = ~(P3_ADD_541_U63 & P3_U4300); 
assign P3_U5830 = ~(P3_ADD_536_U63 & P3_U4301); 
assign P3_U5850 = ~(P3_ADD_558_U65 & P3_U3220); 
assign P3_U5851 = ~(P3_ADD_553_U65 & P3_U4298); 
assign P3_U5852 = ~(P3_ADD_547_U65 & P3_U4299); 
assign P3_U5853 = ~(P3_ADD_541_U62 & P3_U4300); 
assign P3_U5854 = ~(P3_ADD_536_U62 & P3_U4301); 
assign P3_U5855 = ~(P3_ADD_531_U65 & P3_U2354); 
assign P3_U5863 = ~(P3_ADD_385_U65 & P3_U2358); 
assign P3_U5864 = ~(P3_ADD_380_U65 & P3_U2359); 
assign P3_U5865 = ~(P3_ADD_349_U65 & P3_U4306); 
assign P3_U5866 = ~(P3_ADD_344_U65 & P3_U2362); 
assign P3_U5877 = ~(P3_ADD_541_U91 & P3_U4300); 
assign P3_U5878 = ~(P3_ADD_536_U91 & P3_U4301); 
assign P3_U5881 = ~(P3_ADD_515_U91 & P3_U4302); 
assign P3_U5882 = ~(P3_ADD_494_U91 & P3_U2356); 
assign P3_U5883 = ~(P3_ADD_476_U91 & P3_U4303); 
assign P3_U5884 = ~(P3_ADD_441_U91 & P3_U4304); 
assign P3_U5885 = ~(P3_ADD_405_U91 & P3_U4305); 
assign P3_U5886 = ~(P3_ADD_394_U91 & P3_U2357); 
assign P3_U6024 = ~(P3_ADD_526_U75 & P3_U2355); 
assign P3_U6048 = ~(P3_ADD_526_U74 & P3_U2355); 
assign P3_U6666 = ~(P3_U3250 & P3_LWORD_REG_15__SCAN_IN); 
assign P3_U6669 = ~(P3_U3250 & P3_LWORD_REG_14__SCAN_IN); 
assign P3_U6672 = ~(P3_U3250 & P3_LWORD_REG_13__SCAN_IN); 
assign P3_U6675 = ~(P3_U3250 & P3_LWORD_REG_12__SCAN_IN); 
assign P3_U6678 = ~(P3_U3250 & P3_LWORD_REG_11__SCAN_IN); 
assign P3_U6681 = ~(P3_U3250 & P3_LWORD_REG_10__SCAN_IN); 
assign P3_U6684 = ~(P3_U3250 & P3_LWORD_REG_9__SCAN_IN); 
assign P3_U6687 = ~(P3_U3250 & P3_LWORD_REG_8__SCAN_IN); 
assign P3_U6690 = ~(P3_U3250 & P3_LWORD_REG_7__SCAN_IN); 
assign P3_U6693 = ~(P3_U3250 & P3_LWORD_REG_6__SCAN_IN); 
assign P3_U6696 = ~(P3_U3250 & P3_LWORD_REG_5__SCAN_IN); 
assign P3_U6699 = ~(P3_U3250 & P3_LWORD_REG_4__SCAN_IN); 
assign P3_U6702 = ~(P3_U3250 & P3_LWORD_REG_3__SCAN_IN); 
assign P3_U6705 = ~(P3_U3250 & P3_LWORD_REG_2__SCAN_IN); 
assign P3_U6708 = ~(P3_U3250 & P3_LWORD_REG_1__SCAN_IN); 
assign P3_U6711 = ~(P3_U3250 & P3_LWORD_REG_0__SCAN_IN); 
assign P3_U6714 = ~(P3_U3250 & P3_UWORD_REG_14__SCAN_IN); 
assign P3_U6717 = ~(P3_U3250 & P3_UWORD_REG_13__SCAN_IN); 
assign P3_U6720 = ~(P3_U3250 & P3_UWORD_REG_12__SCAN_IN); 
assign P3_U6723 = ~(P3_U3250 & P3_UWORD_REG_11__SCAN_IN); 
assign P3_U6726 = ~(P3_U3250 & P3_UWORD_REG_10__SCAN_IN); 
assign P3_U6729 = ~(P3_U3250 & P3_UWORD_REG_9__SCAN_IN); 
assign P3_U6732 = ~(P3_U3250 & P3_UWORD_REG_8__SCAN_IN); 
assign P3_U6735 = ~(P3_U3250 & P3_UWORD_REG_7__SCAN_IN); 
assign P3_U6738 = ~(P3_U3250 & P3_UWORD_REG_6__SCAN_IN); 
assign P3_U6741 = ~(P3_U3250 & P3_UWORD_REG_5__SCAN_IN); 
assign P3_U6744 = ~(P3_U3250 & P3_UWORD_REG_4__SCAN_IN); 
assign P3_U6747 = ~(P3_U3250 & P3_UWORD_REG_3__SCAN_IN); 
assign P3_U6750 = ~(P3_U3250 & P3_UWORD_REG_2__SCAN_IN); 
assign P3_U6753 = ~(P3_U3250 & P3_UWORD_REG_1__SCAN_IN); 
assign P3_U6756 = ~(P3_U3250 & P3_UWORD_REG_0__SCAN_IN); 
assign P3_U7000 = ~(P3_U3253 & P3_EBX_REG_0__SCAN_IN); 
assign P3_U7003 = ~(P3_U3253 & P3_EBX_REG_1__SCAN_IN); 
assign P3_U7006 = ~(P3_U3253 & P3_EBX_REG_2__SCAN_IN); 
assign P3_U7009 = ~(P3_U3253 & P3_EBX_REG_3__SCAN_IN); 
assign P3_U7012 = ~(P3_U3253 & P3_EBX_REG_4__SCAN_IN); 
assign P3_U7015 = ~(P3_U3253 & P3_EBX_REG_5__SCAN_IN); 
assign P3_U7018 = ~(P3_U3253 & P3_EBX_REG_6__SCAN_IN); 
assign P3_U7021 = ~(P3_U3253 & P3_EBX_REG_7__SCAN_IN); 
assign P3_U7024 = ~(P3_U3253 & P3_EBX_REG_8__SCAN_IN); 
assign P3_U7027 = ~(P3_U3253 & P3_EBX_REG_9__SCAN_IN); 
assign P3_U7030 = ~(P3_U3253 & P3_EBX_REG_10__SCAN_IN); 
assign P3_U7033 = ~(P3_U3253 & P3_EBX_REG_11__SCAN_IN); 
assign P3_U7036 = ~(P3_U3253 & P3_EBX_REG_12__SCAN_IN); 
assign P3_U7039 = ~(P3_U3253 & P3_EBX_REG_13__SCAN_IN); 
assign P3_U7042 = ~(P3_U3253 & P3_EBX_REG_14__SCAN_IN); 
assign P3_U7045 = ~(P3_U3253 & P3_EBX_REG_15__SCAN_IN); 
assign P3_U7048 = ~(P3_U3253 & P3_EBX_REG_16__SCAN_IN); 
assign P3_U7051 = ~(P3_U3253 & P3_EBX_REG_17__SCAN_IN); 
assign P3_U7054 = ~(P3_U3253 & P3_EBX_REG_18__SCAN_IN); 
assign P3_U7057 = ~(P3_U3253 & P3_EBX_REG_19__SCAN_IN); 
assign P3_U7060 = ~(P3_U3253 & P3_EBX_REG_20__SCAN_IN); 
assign P3_U7063 = ~(P3_U3253 & P3_EBX_REG_21__SCAN_IN); 
assign P3_U7066 = ~(P3_U3253 & P3_EBX_REG_22__SCAN_IN); 
assign P3_U7069 = ~(P3_U3253 & P3_EBX_REG_23__SCAN_IN); 
assign P3_U7072 = ~(P3_U3253 & P3_EBX_REG_24__SCAN_IN); 
assign P3_U7075 = ~(P3_U3253 & P3_EBX_REG_25__SCAN_IN); 
assign P3_U7078 = ~(P3_U3253 & P3_EBX_REG_26__SCAN_IN); 
assign P3_U7081 = ~(P3_U3253 & P3_EBX_REG_27__SCAN_IN); 
assign P3_U7084 = ~(P3_U3253 & P3_EBX_REG_28__SCAN_IN); 
assign P3_U7087 = ~(P3_U3253 & P3_EBX_REG_29__SCAN_IN); 
assign P3_U7090 = ~(P3_U3253 & P3_EBX_REG_30__SCAN_IN); 
assign P3_U7092 = ~(P3_U3253 & P3_EBX_REG_31__SCAN_IN); 
assign P3_U7093 = ~(P3_U5488 & P3_U5491); 
assign P3_U7946 = ~(P3_U4539 & P3_U4618); 
assign P2_U3538 = ~(P2_U4055 & P2_U2446); 
assign P2_U4456 = ~(P2_U2446 & P2_U2359); 
assign P2_U4609 = ~(P2_U4603 & P2_U3520); 
assign P2_U6228 = ~(P2_U4058 & P2_U2446); 
assign P2_U6860 = ~(P2_U4189 & P2_U2446); 
assign P2_U8055 = ~(P2_U3289 & P2_U3520); 
assign P2_U8145 = ~(P2_U7873 & P2_U3520); 
assign P2_U8415 = ~(P2_R2337_U89 & P2_U3284); 
assign P1_U2618 = ~(P1_U6747 & P1_U4002); 
assign P1_U4499 = ~P1_U3437; 
assign P1_U6858 = ~(P1_R2337_U91 & P1_U2352); 
assign P1_U6878 = ~(P1_ADD_371_U19 & P1_U4208); 
assign P1_U7679 = ~(P1_U4494 & P1_U3437); 
assign P3_ADD_526_U36 = ~(P3_ADD_526_U90 & P3_ADD_526_U114); 
assign P3_ADD_526_U105 = ~(P3_ADD_526_U114 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_526_U183 = ~(P3_ADD_526_U114 & P3_ADD_526_U33); 
assign P3_ADD_526_U186 = ~(P3_ADD_526_U136 & P3_ADD_526_U29); 
assign P3_ADD_552_U36 = ~(P3_ADD_552_U90 & P3_ADD_552_U114); 
assign P3_ADD_552_U105 = ~(P3_ADD_552_U114 & P3_EBX_REG_19__SCAN_IN); 
assign P3_ADD_552_U183 = ~(P3_ADD_552_U114 & P3_ADD_552_U33); 
assign P3_ADD_552_U186 = ~(P3_ADD_552_U136 & P3_ADD_552_U29); 
assign P3_ADD_546_U36 = ~(P3_ADD_546_U90 & P3_ADD_546_U114); 
assign P3_ADD_546_U105 = ~(P3_ADD_546_U114 & P3_EAX_REG_19__SCAN_IN); 
assign P3_ADD_546_U183 = ~(P3_ADD_546_U114 & P3_ADD_546_U33); 
assign P3_ADD_546_U186 = ~(P3_ADD_546_U136 & P3_ADD_546_U29); 
assign P3_ADD_391_1180_U22 = ~(P3_ADD_391_1180_U44 & P3_ADD_391_1180_U43); 
assign P3_ADD_391_1180_U31 = ~P3_ADD_391_1180_U12; 
assign P3_ADD_391_1180_U41 = ~(P3_U2617 & P3_ADD_391_1180_U12); 
assign P3_ADD_476_U24 = ~(P3_ADD_476_U102 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_476_U180 = ~(P3_ADD_476_U102 & P3_ADD_476_U23); 
assign P3_ADD_531_U25 = ~(P3_ADD_531_U106 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_531_U189 = ~(P3_ADD_531_U106 & P3_ADD_531_U24); 
assign P3_SUB_320_U49 = ~P3_ADD_318_U91; 
assign P3_SUB_320_U53 = P3_SUB_320_U129 & P3_SUB_320_U128; 
assign P3_SUB_320_U126 = ~(P3_ADD_318_U91 & P3_SUB_320_U125); 
assign P3_ADD_318_U24 = ~(P3_ADD_318_U102 & P3_PHYADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_318_U180 = ~(P3_ADD_318_U102 & P3_ADD_318_U23); 
assign P3_ADD_315_U24 = ~(P3_ADD_315_U99 & P3_PHYADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_315_U172 = ~(P3_ADD_315_U99 & P3_ADD_315_U23); 
assign P3_ADD_360_1242_U41 = ~(P3_ADD_360_1242_U40 & P3_ADD_360_1242_U133); 
assign P3_ADD_360_1242_U91 = ~(P3_ADD_360_1242_U237 & P3_ADD_360_1242_U236); 
assign P3_ADD_360_1242_U93 = P3_ADD_360_1242_U133 & P3_ADD_360_1242_U123; 
assign P3_ADD_360_1242_U96 = P3_ADD_360_1242_U125 & P3_ADD_360_1242_U123; 
assign P3_ADD_360_1242_U132 = ~P3_ADD_360_1242_U40; 
assign P3_ADD_360_1242_U190 = ~(P3_ADD_360_1242_U92 & P3_ADD_360_1242_U123); 
assign P3_ADD_360_1242_U223 = ~(P3_ADD_360_1242_U20 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_467_U24 = ~(P3_ADD_467_U102 & P3_REIP_REG_11__SCAN_IN); 
assign P3_ADD_467_U180 = ~(P3_ADD_467_U102 & P3_ADD_467_U23); 
assign P3_ADD_430_U24 = ~(P3_ADD_430_U102 & P3_REIP_REG_11__SCAN_IN); 
assign P3_ADD_430_U180 = ~(P3_ADD_430_U102 & P3_ADD_430_U23); 
assign P3_ADD_380_U25 = ~(P3_ADD_380_U106 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_380_U189 = ~(P3_ADD_380_U106 & P3_ADD_380_U24); 
assign P3_ADD_344_U25 = ~(P3_ADD_344_U106 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_344_U189 = ~(P3_ADD_344_U106 & P3_ADD_344_U24); 
assign P3_ADD_339_U24 = ~(P3_ADD_339_U102 & P3_PHYADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_339_U180 = ~(P3_ADD_339_U102 & P3_ADD_339_U23); 
assign P3_ADD_360_U18 = ~(P3_ADD_360_U34 & P3_ADD_360_U33); 
assign P3_ADD_360_U27 = ~P3_ADD_360_U13; 
assign P3_ADD_360_U31 = ~(P3_U2627 & P3_ADD_360_U13); 
assign P3_ADD_541_U24 = ~(P3_ADD_541_U102 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_541_U180 = ~(P3_ADD_541_U102 & P3_ADD_541_U23); 
assign P3_SUB_357_1258_U5 = P3_SUB_357_1258_U188 & P3_SUB_357_1258_U186; 
assign P3_SUB_357_1258_U6 = P3_SUB_357_1258_U187 & P3_SUB_357_1258_U178; 
assign P3_SUB_357_1258_U10 = P3_SUB_357_1258_U210 & P3_SUB_357_1258_U205 & P3_SUB_357_1258_U206 & P3_SUB_357_1258_U156; 
assign P3_SUB_357_1258_U21 = ~(P3_SUB_357_1258_U426 & P3_SUB_357_1258_U425 & P3_SUB_357_1258_U307); 
assign P3_SUB_357_1258_U37 = ~P3_ADD_357_U17; 
assign P3_SUB_357_1258_U96 = P3_SUB_357_1258_U168 & P3_SUB_357_1258_U162; 
assign P3_SUB_357_1258_U99 = P3_SUB_357_1258_U192 & P3_SUB_357_1258_U155; 
assign P3_SUB_357_1258_U102 = P3_SUB_357_1258_U199 & P3_SUB_357_1258_U56; 
assign P3_SUB_357_1258_U105 = P3_SUB_357_1258_U157 & P3_SUB_357_1258_U58 & P3_SUB_357_1258_U219; 
assign P3_SUB_357_1258_U106 = P3_SUB_357_1258_U219 & P3_SUB_357_1258_U157; 
assign P3_SUB_357_1258_U107 = P3_SUB_357_1258_U60 & P3_SUB_357_1258_U269 & P3_INSTADDRPOINTER_REG_31__SCAN_IN; 
assign P3_SUB_357_1258_U124 = ~(P3_SUB_357_1258_U181 & P3_SUB_357_1258_U180); 
assign P3_SUB_357_1258_U125 = ~(P3_SUB_357_1258_U159 & P3_SUB_357_1258_U183); 
assign P3_SUB_357_1258_U153 = ~(P3_SUB_357_1258_U217 & P3_SUB_357_1258_U39); 
assign P3_SUB_357_1258_U154 = ~(P3_SUB_357_1258_U191 & P3_SUB_357_1258_U39); 
assign P3_SUB_357_1258_U167 = ~(P3_SUB_357_1258_U94 & P3_SUB_357_1258_U166); 
assign P3_SUB_357_1258_U171 = P3_ADD_357_U17 | P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_SUB_357_1258_U173 = ~(P3_ADD_357_U17 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_SUB_357_1258_U209 = ~(P3_SUB_357_1258_U39 & P3_SUB_357_1258_U208); 
assign P3_SUB_357_1258_U243 = ~(P3_SUB_357_1258_U57 & P3_SUB_357_1258_U39); 
assign P3_SUB_357_1258_U258 = ~(P3_SUB_357_1258_U179 & P3_SUB_357_1258_U178); 
assign P3_SUB_357_1258_U262 = ~(P3_SUB_357_1258_U234 & P3_SUB_357_1258_U157); 
assign P3_SUB_357_1258_U263 = ~(P3_SUB_357_1258_U245 & P3_SUB_357_1258_U206); 
assign P3_SUB_357_1258_U264 = ~(P3_SUB_357_1258_U256 & P3_SUB_357_1258_U155); 
assign P3_SUB_357_1258_U265 = ~(P3_SUB_357_1258_U257 & P3_SUB_357_1258_U187); 
assign P3_SUB_357_1258_U309 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_SUB_357_1258_U314 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_SUB_357_1258_U316 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_SUB_357_1258_U328 = ~(P3_ADD_357_U17 & P3_SUB_357_1258_U38); 
assign P3_SUB_357_1258_U330 = ~(P3_ADD_357_U17 & P3_SUB_357_1258_U38); 
assign P3_SUB_357_1258_U334 = ~(P3_SUB_357_1258_U24 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_SUB_357_1258_U336 = ~(P3_SUB_357_1258_U24 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_SUB_357_1258_U343 = ~(P3_SUB_357_1258_U342 & P3_SUB_357_1258_U341); 
assign P3_SUB_357_1258_U351 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_SUB_357_1258_U356 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_SUB_357_1258_U358 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_SUB_357_1258_U366 = ~(P3_SUB_357_1258_U165 & P3_SUB_357_1258_U364); 
assign P3_SUB_357_1258_U368 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_SUB_357_1258_U370 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_SUB_357_1258_U374 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_SUB_357_1258_U378 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_SUB_357_1258_U380 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_SUB_357_1258_U385 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_SUB_357_1258_U387 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_SUB_357_1258_U392 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_SUB_357_1258_U394 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_SUB_357_1258_U399 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_SUB_357_1258_U401 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_SUB_357_1258_U406 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_SUB_357_1258_U408 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_SUB_357_1258_U413 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_SUB_357_1258_U415 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_SUB_357_1258_U420 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_SUB_357_1258_U427 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_SUB_357_1258_U432 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_SUB_357_1258_U434 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_SUB_357_1258_U439 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_SUB_357_1258_U443 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_SUB_357_1258_U445 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_SUB_357_1258_U450 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_SUB_357_1258_U452 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_SUB_357_1258_U457 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_SUB_357_1258_U459 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_SUB_357_1258_U464 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_SUB_357_1258_U466 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_SUB_357_1258_U471 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_SUB_357_1258_U473 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_SUB_357_1258_U478 = ~(P3_SUB_357_1258_U39 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_515_U24 = ~(P3_ADD_515_U102 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_515_U180 = ~(P3_ADD_515_U102 & P3_ADD_515_U23); 
assign P3_ADD_394_U24 = ~(P3_ADD_394_U105 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_394_U184 = ~(P3_ADD_394_U105 & P3_ADD_394_U23); 
assign P3_SUB_414_U10 = P3_SUB_414_U118 & P3_SUB_414_U32; 
assign P3_SUB_414_U33 = ~(P3_SUB_414_U44 & P3_SUB_414_U73 & P3_SUB_414_U97); 
assign P3_SUB_414_U115 = ~(P3_SUB_414_U97 & P3_SUB_414_U73); 
assign P3_SUB_414_U151 = ~(P3_SUB_414_U97 & P3_SUB_414_U73); 
assign P3_ADD_441_U24 = ~(P3_ADD_441_U102 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_441_U180 = ~(P3_ADD_441_U102 & P3_ADD_441_U23); 
assign P3_ADD_349_U25 = ~(P3_ADD_349_U106 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_349_U189 = ~(P3_ADD_349_U106 & P3_ADD_349_U24); 
assign P3_ADD_405_U24 = ~(P3_ADD_405_U105 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_405_U184 = ~(P3_ADD_405_U105 & P3_ADD_405_U23); 
assign P3_ADD_553_U25 = ~(P3_ADD_553_U106 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_553_U189 = ~(P3_ADD_553_U106 & P3_ADD_553_U24); 
assign P3_ADD_558_U25 = ~(P3_ADD_558_U106 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_558_U189 = ~(P3_ADD_558_U106 & P3_ADD_558_U24); 
assign P3_ADD_385_U25 = ~(P3_ADD_385_U106 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_385_U189 = ~(P3_ADD_385_U106 & P3_ADD_385_U24); 
assign P3_ADD_357_U9 = P3_ADD_357_U25 & P3_ADD_357_U6; 
assign P3_ADD_547_U25 = ~(P3_ADD_547_U106 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_ADD_547_U189 = ~(P3_ADD_547_U106 & P3_ADD_547_U24); 
assign P3_ADD_371_1212_U98 = P3_ADD_371_1212_U235 & P3_ADD_371_1212_U234 & P3_ADD_371_1212_U29; 
assign P3_ADD_371_1212_U124 = ~P3_ADD_371_1212_U44; 
assign P3_ADD_371_1212_U128 = ~(P3_ADD_371_1212_U127 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_ADD_371_1212_U130 = ~(P3_ADD_371_1212_U44 & P3_ADD_371_1212_U119); 
assign P3_ADD_371_1212_U134 = ~P3_ADD_371_1212_U24; 
assign P3_ADD_371_1212_U158 = ~(P3_ADD_371_1212_U157 & P3_ADD_371_1212_U44); 
assign P3_ADD_371_1212_U197 = ~(P3_ADD_371_1212_U156 & P3_ADD_371_1212_U24); 
assign P3_ADD_371_1212_U229 = ~(P3_ADD_371_1212_U21 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_ADD_371_1212_U243 = ~(P3_ADD_371_1212_U199 & P3_ADD_371_1212_U44); 
assign P3_ADD_371_U19 = ~(P3_ADD_371_U38 & P3_ADD_371_U37); 
assign P3_ADD_371_U30 = ~P3_ADD_371_U13; 
assign P3_ADD_371_U35 = ~(P3_U2627 & P3_ADD_371_U13); 
assign P3_ADD_494_U24 = ~(P3_ADD_494_U102 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_494_U180 = ~(P3_ADD_494_U102 & P3_ADD_494_U23); 
assign P3_ADD_536_U24 = ~(P3_ADD_536_U102 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_536_U180 = ~(P3_ADD_536_U102 & P3_ADD_536_U23); 
assign P3_ADD_402_1132_U22 = ~(P3_ADD_402_1132_U44 & P3_ADD_402_1132_U43); 
assign P3_ADD_402_1132_U31 = ~P3_ADD_402_1132_U12; 
assign P3_ADD_402_1132_U41 = ~(P3_U2617 & P3_ADD_402_1132_U12); 
assign P2_R2099_U108 = ~P2_R2099_U106; 
assign P2_R2099_U109 = ~(P2_R2099_U9 & P2_R2099_U105); 
assign P2_R2099_U147 = ~P2_R2099_U105; 
assign P2_R2099_U161 = ~(P2_U2744 & P2_R2099_U12); 
assign P2_R2099_U163 = ~(P2_U2744 & P2_R2099_U12); 
assign P2_R2099_U172 = ~(P2_U2745 & P2_R2099_U10); 
assign P2_R2099_U174 = ~(P2_U2745 & P2_R2099_U10); 
assign P2_R2099_U199 = ~(P2_U2750 & P2_R2099_U105); 
assign P2_R2099_U202 = ~(P2_U2746 & P2_R2099_U105 & P2_R2099_U8); 
assign P2_R2099_U224 = ~(P2_U2751 & P2_R2099_U6); 
assign P2_ADD_402_1132_U21 = ~(P2_ADD_402_1132_U42 & P2_ADD_402_1132_U41); 
assign P2_ADD_402_1132_U31 = ~P2_ADD_402_1132_U12; 
assign P2_ADD_402_1132_U43 = ~(P2_U2595 & P2_ADD_402_1132_U12); 
assign P2_R2182_U56 = ~P2_U2687; 
assign P2_R2182_U118 = P2_R2182_U260 & P2_R2182_U259; 
assign P2_R2182_U120 = P2_R2182_U267 & P2_R2182_U266; 
assign P2_R2182_U163 = P2_U2687 | P2_U2663; 
assign P2_R2182_U165 = ~(P2_U2663 & P2_U2687); 
assign P2_R2182_U253 = ~(P2_U2687 & P2_R2182_U57); 
assign P2_R2182_U255 = ~(P2_U2687 & P2_R2182_U57); 
assign P2_R2182_U263 = ~(P2_R2182_U262 & P2_R2182_U261); 
assign P2_R2182_U270 = ~(P2_R2182_U269 & P2_R2182_U268); 
assign P2_R2167_U19 = ~(P2_U2714 & P2_U2715); 
assign P2_R2167_U21 = P2_U2714 | P2_U2715; 
assign P2_R2027_U25 = ~(P2_R2027_U106 & P2_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P2_R2027_U189 = ~(P2_R2027_U106 & P2_R2027_U24); 
assign P2_R2337_U25 = ~(P2_R2337_U103 & P2_PHYADDRPOINTER_REG_12__SCAN_IN); 
assign P2_R2337_U178 = ~(P2_R2337_U103 & P2_R2337_U24); 
assign P2_R2219_U30 = ~(P2_R2219_U116 & P2_R2219_U115); 
assign P2_R2219_U42 = ~(P2_R2219_U19 & P2_R2219_U71); 
assign P2_R2219_U43 = ~(P2_R2219_U50 & P2_R2219_U49); 
assign P2_R2219_U75 = ~(P2_R2219_U73 & P2_R2219_U55); 
assign P2_R2219_U110 = ~(P2_R2219_U79 & P2_R2219_U109); 
assign P2_R2096_U51 = ~(P2_R2096_U114 & P2_R2096_U170); 
assign P2_R2096_U109 = ~(P2_R2096_U122 & P2_R2096_U121); 
assign P2_R2096_U218 = ~(P2_R2096_U119 & P2_R2096_U216); 
assign P2_R1957_U48 = ~P2_U3681; 
assign P2_R1957_U53 = P2_R1957_U129 & P2_R1957_U128; 
assign P2_R1957_U126 = ~(P2_U3681 & P2_R1957_U125); 
assign P2_ADD_394_U24 = ~(P2_ADD_394_U105 & P2_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P2_ADD_394_U148 = ~(P2_ADD_394_U105 & P2_ADD_394_U23); 
assign P2_R2267_U22 = ~P2_U3646; 
assign P2_R2267_U77 = ~(P2_U3646 & P2_R2267_U42); 
assign P1_R2027_U36 = ~(P1_R2027_U90 & P1_R2027_U114); 
assign P1_R2027_U105 = ~(P1_R2027_U114 & P1_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P1_R2027_U183 = ~(P1_R2027_U114 & P1_R2027_U33); 
assign P1_R2027_U186 = ~(P1_R2027_U136 & P1_R2027_U29); 
assign P1_R2182_U10 = ~P1_U2742; 
assign P1_R2182_U32 = ~(P1_R2182_U82 & P1_R2182_U81); 
assign P1_R2182_U34 = ~(P1_R2182_U86 & P1_R2182_U85); 
assign P1_R2182_U35 = P1_U2742 & P1_U2741; 
assign P1_R2182_U45 = ~(P1_R2182_U51 & P1_R2182_U62); 
assign P1_R2182_U46 = ~P1_R2182_U19; 
assign P1_R2182_U53 = ~(P1_R2182_U50 & P1_R2182_U51); 
assign P1_R2182_U59 = ~P1_R2182_U44; 
assign P1_R2182_U78 = ~(P1_U2736 & P1_R2182_U19); 
assign P1_R2182_U79 = ~(P1_U2737 & P1_R2182_U44); 
assign P1_R2144_U7 = P1_R2144_U104 & P1_R2144_U81; 
assign P1_R2144_U19 = ~(P1_U2748 & P1_R2144_U178); 
assign P1_R2144_U21 = ~(P1_U2747 & P1_R2144_U170); 
assign P1_R2144_U23 = ~(P1_U2746 & P1_R2144_U173); 
assign P1_R2144_U52 = P1_R2144_U106 & P1_R2144_U105; 
assign P1_R2144_U102 = ~P1_R2144_U81; 
assign P1_R2144_U103 = ~(P1_U2745 & P1_R2144_U181); 
assign P1_R2358_U444 = ~(P1_U2352 & P1_R2358_U152); 
assign P1_R2358_U446 = ~(P1_U2352 & P1_R2358_U152); 
assign P1_R2099_U7 = ~(P1_R2099_U88 & P1_R2099_U137); 
assign P1_R2099_U87 = ~(P1_R2099_U324 & P1_R2099_U323); 
assign P1_R2099_U112 = ~(P1_R2099_U35 & P1_R2099_U137); 
assign P1_R2099_U153 = ~P1_R2099_U137; 
assign P1_R2099_U297 = ~(P1_R2099_U35 & P1_R2099_U137); 
assign P1_R2167_U37 = ~(P1_R2167_U20 & P1_R2167_U34); 
assign P1_R2337_U24 = ~(P1_R2337_U102 & P1_PHYADDRPOINTER_REG_11__SCAN_IN); 
assign P1_R2337_U180 = ~(P1_R2337_U102 & P1_R2337_U23); 
assign P1_R2096_U24 = ~(P1_R2096_U102 & P1_REIP_REG_11__SCAN_IN); 
assign P1_R2096_U180 = ~(P1_R2096_U102 & P1_R2096_U23); 
assign P1_ADD_371_U6 = P1_ADD_371_U22 & P1_ADD_371_U30; 
assign P1_ADD_371_U25 = ~(P1_ADD_371_U30 & P1_U3233); 
assign P1_ADD_371_U34 = ~(P1_ADD_371_U30 & P1_ADD_371_U13); 
assign P1_ADD_405_U24 = ~(P1_ADD_405_U105 & P1_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P1_ADD_405_U148 = ~(P1_ADD_405_U105 & P1_ADD_405_U23); 
assign P1_ADD_515_U24 = ~(P1_ADD_515_U102 & P1_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P1_ADD_515_U146 = ~(P1_ADD_515_U102 & P1_ADD_515_U23); 
assign P3_U2382 = P3_U3951 & P3_U3249; 
assign P3_U2386 = P3_U3249 & P3_STATE2_REG_1__SCAN_IN; 
assign P3_U2387 = P3_U3953 & P3_U3249; 
assign P3_U2388 = P3_U3952 & P3_U3249; 
assign P3_U2389 = P3_U4354 & P3_U3249; 
assign P3_U2399 = P3_U4309 & P3_U4573; 
assign P3_U2406 = P3_U4311 & P3_U3104; 
assign P3_U2407 = P3_U4311 & P3_U4505; 
assign P3_U2408 = P3_U4309 & P3_U3218; 
assign P3_U2409 = P3_U3251 & P3_STATE2_REG_0__SCAN_IN; 
assign P3_U2410 = P3_U3251 & P3_U3121; 
assign P3_U2518 = P3_U3668 & P3_U5522; 
assign P3_U3512 = P3_U3511 & P3_U5088; 
assign P3_U3514 = P3_U3513 & P3_U5093; 
assign P3_U3516 = P3_U3515 & P3_U5098; 
assign P3_U3518 = P3_U3517 & P3_U5103; 
assign P3_U3520 = P3_U3519 & P3_U5108; 
assign P3_U3522 = P3_U3521 & P3_U5113; 
assign P3_U3524 = P3_U3523 & P3_U5118; 
assign P3_U3526 = P3_U3525 & P3_U5123; 
assign P3_U3530 = P3_U3529 & P3_U5140; 
assign P3_U3532 = P3_U3531 & P3_U5145; 
assign P3_U3534 = P3_U3533 & P3_U5150; 
assign P3_U3536 = P3_U3535 & P3_U5155; 
assign P3_U3538 = P3_U3537 & P3_U5160; 
assign P3_U3540 = P3_U3539 & P3_U5165; 
assign P3_U3542 = P3_U3541 & P3_U5170; 
assign P3_U3544 = P3_U3543 & P3_U5175; 
assign P3_U3548 = P3_U3547 & P3_U5192; 
assign P3_U3550 = P3_U3549 & P3_U5197; 
assign P3_U3552 = P3_U3551 & P3_U5202; 
assign P3_U3554 = P3_U3553 & P3_U5207; 
assign P3_U3556 = P3_U3555 & P3_U5212; 
assign P3_U3558 = P3_U3557 & P3_U5217; 
assign P3_U3560 = P3_U3559 & P3_U5222; 
assign P3_U3562 = P3_U3561 & P3_U5227; 
assign P3_U3566 = P3_U3565 & P3_U5242; 
assign P3_U3568 = P3_U3567 & P3_U5247; 
assign P3_U3570 = P3_U3569 & P3_U5252; 
assign P3_U3572 = P3_U3571 & P3_U5257; 
assign P3_U3574 = P3_U3573 & P3_U5262; 
assign P3_U3576 = P3_U3575 & P3_U5267; 
assign P3_U3578 = P3_U3577 & P3_U5272; 
assign P3_U3580 = P3_U3579 & P3_U5277; 
assign P3_U3584 = P3_U3583 & P3_U5293; 
assign P3_U3586 = P3_U3585 & P3_U5298; 
assign P3_U3588 = P3_U3587 & P3_U5303; 
assign P3_U3590 = P3_U3589 & P3_U5308; 
assign P3_U3592 = P3_U3591 & P3_U5313; 
assign P3_U3594 = P3_U3593 & P3_U5318; 
assign P3_U3596 = P3_U3595 & P3_U5323; 
assign P3_U3598 = P3_U3597 & P3_U5328; 
assign P3_U3601 = P3_U3600 & P3_U5344; 
assign P3_U3603 = P3_U3602 & P3_U5349; 
assign P3_U3605 = P3_U3604 & P3_U5354; 
assign P3_U3607 = P3_U3606 & P3_U5359; 
assign P3_U3609 = P3_U3608 & P3_U5364; 
assign P3_U3611 = P3_U3610 & P3_U5369; 
assign P3_U3613 = P3_U3612 & P3_U5374; 
assign P3_U3615 = P3_U3614 & P3_U5379; 
assign P3_U3619 = P3_U3618 & P3_U5395; 
assign P3_U3621 = P3_U3620 & P3_U5400; 
assign P3_U3623 = P3_U3622 & P3_U5405; 
assign P3_U3625 = P3_U3624 & P3_U5410; 
assign P3_U3627 = P3_U3626 & P3_U5415; 
assign P3_U3629 = P3_U3628 & P3_U5420; 
assign P3_U3631 = P3_U3630 & P3_U5425; 
assign P3_U3633 = P3_U3632 & P3_U5430; 
assign P3_U3637 = P3_U3636 & P3_U5445; 
assign P3_U3639 = P3_U3638 & P3_U5450; 
assign P3_U3641 = P3_U3640 & P3_U5455; 
assign P3_U3643 = P3_U3642 & P3_U5460; 
assign P3_U3645 = P3_U3644 & P3_U5465; 
assign P3_U3647 = P3_U3646 & P3_U5470; 
assign P3_U3649 = P3_U3648 & P3_U5475; 
assign P3_U3651 = P3_U3650 & P3_U5480; 
assign P3_U3675 = P3_U5538 & P3_U5536; 
assign P3_U3693 = P3_U5638 & P3_U5637 & P3_U3694 & P3_U5633 & P3_U5632; 
assign P3_U3705 = P3_U3704 & P3_U3703 & P3_U5675; 
assign P3_U3710 = P3_U5686 & P3_U5685 & P3_U3708; 
assign P3_U3718 = P3_U5710 & P3_U5709 & P3_U3716; 
assign P3_U3726 = P3_U5734 & P3_U5733 & P3_U3724; 
assign P3_U3734 = P3_U5758 & P3_U5757 & P3_U3732; 
assign P3_U3742 = P3_U5782 & P3_U5781 & P3_U3740; 
assign P3_U3750 = P3_U5806 & P3_U5805 & P3_U3748; 
assign P3_U3757 = P3_U5830 & P3_U5829 & P3_U3756; 
assign P3_U3762 = P3_U5852 & P3_U5851; 
assign P3_U3764 = P3_U5854 & P3_U5853 & P3_U5855 & P3_U3763; 
assign P3_U3766 = P3_U5866 & P3_U5865 & P3_U5864 & P3_U5863; 
assign P3_U3770 = P3_U5881 & P3_U5880; 
assign P3_U3772 = P3_U5883 & P3_U5882 & P3_U5884 & P3_U5886 & P3_U5885; 
assign P3_U4290 = ~(P3_U2515 & P3_U2516 & P3_U3657); 
assign P3_U4334 = ~(P3_U2390 & P3_U7093); 
assign P3_U4623 = ~P3_U3262; 
assign P3_U4672 = ~(P3_U3369 & P3_U4670); 
assign P3_U4674 = ~(P3_U2489 & P3_U4673); 
assign P3_U4724 = ~(P3_U3387 & P3_U4722); 
assign P3_U4726 = ~(P3_U2489 & P3_U4725); 
assign P3_U4776 = ~(P3_U3405 & P3_U4774); 
assign P3_U4778 = ~(P3_U2489 & P3_U4777); 
assign P3_U4827 = ~(P3_U3423 & P3_U4825); 
assign P3_U4829 = ~(P3_U2489 & P3_U4828); 
assign P3_U4879 = ~(P3_U3440 & P3_U4877); 
assign P3_U4881 = ~(P3_U2489 & P3_U4880); 
assign P3_U4931 = ~(P3_U3458 & P3_U4929); 
assign P3_U4933 = ~(P3_U2489 & P3_U4932); 
assign P3_U4983 = ~(P3_U3476 & P3_U4981); 
assign P3_U4985 = ~(P3_U2489 & P3_U4984); 
assign P3_U5034 = ~(P3_U3493 & P3_U5032); 
assign P3_U5036 = ~(P3_U2489 & P3_U5035); 
assign P3_U5081 = ~(P3_U5078 & P3_U5080); 
assign P3_U5084 = ~(P3_U5079 & P3_U4322); 
assign P3_U5133 = ~(P3_U5129 & P3_U5132); 
assign P3_U5136 = ~(P3_U5131 & P3_U4322); 
assign P3_U5185 = ~(P3_U5181 & P3_U5184); 
assign P3_U5188 = ~(P3_U5183 & P3_U4322); 
assign P3_U5236 = ~(P3_U5235 & P3_U3072); 
assign P3_U5287 = ~(P3_U5283 & P3_U5286); 
assign P3_U5338 = ~(P3_U5334 & P3_U5337); 
assign P3_U5389 = ~(P3_U5385 & P3_U5388); 
assign P3_U5439 = ~(P3_U5438 & P3_U3073); 
assign P3_U5535 = ~(P3_U3672 & P3_U5522); 
assign P3_U5549 = ~(P3_U5534 & P3_U5522); 
assign P3_U5589 = ~(P3_U3685 & P3_U5586); 
assign P3_U5628 = ~(P3_U4539 & P3_U5624); 
assign P3_U5657 = ~(P3_SUB_357_1258_U21 & P3_U2393); 
assign P3_U5680 = ~(P3_ADD_360_1242_U91 & P3_U2395); 
assign P3_U6404 = ~P3_U3249; 
assign P3_U6759 = ~P3_U3251; 
assign P3_U6853 = ~(P3_U2516 & P3_U3243); 
assign P3_U7947 = ~(P3_U4620 & P3_U3101); 
assign P2_U2686 = P2_ADD_402_1132_U21 & P2_U2355; 
assign P2_U3680 = ~(P2_U8416 & P2_U8415); 
assign P2_U3870 = P2_U4460 & P2_U4456; 
assign P2_U3894 = P2_U4460 & P2_U5668 & P2_U4456; 
assign P2_U4190 = P2_U6860 & P2_U3534; 
assign P2_U4442 = ~P2_U3538; 
assign P2_U5659 = ~(P2_R2096_U51 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U6136 = ~(P2_U3538 & P2_LWORD_REG_15__SCAN_IN); 
assign P2_U6139 = ~(P2_U3538 & P2_LWORD_REG_14__SCAN_IN); 
assign P2_U6142 = ~(P2_U3538 & P2_LWORD_REG_13__SCAN_IN); 
assign P2_U6145 = ~(P2_U3538 & P2_LWORD_REG_12__SCAN_IN); 
assign P2_U6148 = ~(P2_U3538 & P2_LWORD_REG_11__SCAN_IN); 
assign P2_U6151 = ~(P2_U3538 & P2_LWORD_REG_10__SCAN_IN); 
assign P2_U6154 = ~(P2_U3538 & P2_LWORD_REG_9__SCAN_IN); 
assign P2_U6157 = ~(P2_U3538 & P2_LWORD_REG_8__SCAN_IN); 
assign P2_U6160 = ~(P2_U3538 & P2_LWORD_REG_7__SCAN_IN); 
assign P2_U6163 = ~(P2_U3538 & P2_LWORD_REG_6__SCAN_IN); 
assign P2_U6166 = ~(P2_U3538 & P2_LWORD_REG_5__SCAN_IN); 
assign P2_U6169 = ~(P2_U3538 & P2_LWORD_REG_4__SCAN_IN); 
assign P2_U6172 = ~(P2_U3538 & P2_LWORD_REG_3__SCAN_IN); 
assign P2_U6175 = ~(P2_U3538 & P2_LWORD_REG_2__SCAN_IN); 
assign P2_U6178 = ~(P2_U3538 & P2_LWORD_REG_1__SCAN_IN); 
assign P2_U6181 = ~(P2_U3538 & P2_LWORD_REG_0__SCAN_IN); 
assign P2_U6184 = ~(P2_U3538 & P2_UWORD_REG_14__SCAN_IN); 
assign P2_U6187 = ~(P2_U3538 & P2_UWORD_REG_13__SCAN_IN); 
assign P2_U6190 = ~(P2_U3538 & P2_UWORD_REG_12__SCAN_IN); 
assign P2_U6193 = ~(P2_U3538 & P2_UWORD_REG_11__SCAN_IN); 
assign P2_U6196 = ~(P2_U3538 & P2_UWORD_REG_10__SCAN_IN); 
assign P2_U6199 = ~(P2_U3538 & P2_UWORD_REG_9__SCAN_IN); 
assign P2_U6202 = ~(P2_U3538 & P2_UWORD_REG_8__SCAN_IN); 
assign P2_U6205 = ~(P2_U3538 & P2_UWORD_REG_7__SCAN_IN); 
assign P2_U6208 = ~(P2_U3538 & P2_UWORD_REG_6__SCAN_IN); 
assign P2_U6211 = ~(P2_U3538 & P2_UWORD_REG_5__SCAN_IN); 
assign P2_U6214 = ~(P2_U3538 & P2_UWORD_REG_4__SCAN_IN); 
assign P2_U6217 = ~(P2_U3538 & P2_UWORD_REG_3__SCAN_IN); 
assign P2_U6220 = ~(P2_U3538 & P2_UWORD_REG_2__SCAN_IN); 
assign P2_U6223 = ~(P2_U3538 & P2_UWORD_REG_1__SCAN_IN); 
assign P2_U6226 = ~(P2_U3538 & P2_UWORD_REG_0__SCAN_IN); 
assign P2_U7725 = ~(P2_R2219_U30 & P2_U7723); 
assign P2_U8343 = ~(P2_R2219_U30 & P2_U2617); 
assign P1_U3318 = ~P1_R2182_U34; 
assign P1_U4026 = P1_U6858 & P1_U6857; 
assign P1_U5530 = ~(P1_R2182_U34 & P1_U7509); 
assign P1_U5555 = ~(P1_R2182_U34 & P1_U5538); 
assign P1_U6800 = ~(P1_R2182_U32 & P1_U6746); 
assign P1_U6864 = ~(P1_R2182_U34 & P1_U6746); 
assign P1_U6872 = ~(P1_ADD_371_U6 & P1_U4208); 
assign P1_U7046 = ~(P1_R2182_U34 & P1_U3294); 
assign P3_ADD_526_U72 = ~(P3_ADD_526_U184 & P3_ADD_526_U183); 
assign P3_ADD_526_U73 = ~(P3_ADD_526_U186 & P3_ADD_526_U185); 
assign P3_ADD_526_U121 = ~P3_ADD_526_U36; 
assign P3_ADD_526_U135 = ~P3_ADD_526_U105; 
assign P3_ADD_526_U178 = ~(P3_ADD_526_U36 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_526_U179 = ~(P3_ADD_526_U105 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_552_U72 = ~(P3_ADD_552_U184 & P3_ADD_552_U183); 
assign P3_ADD_552_U73 = ~(P3_ADD_552_U186 & P3_ADD_552_U185); 
assign P3_ADD_552_U121 = ~P3_ADD_552_U36; 
assign P3_ADD_552_U135 = ~P3_ADD_552_U105; 
assign P3_ADD_552_U178 = ~(P3_ADD_552_U36 & P3_EBX_REG_21__SCAN_IN); 
assign P3_ADD_552_U179 = ~(P3_ADD_552_U105 & P3_EBX_REG_20__SCAN_IN); 
assign P3_ADD_546_U72 = ~(P3_ADD_546_U184 & P3_ADD_546_U183); 
assign P3_ADD_546_U73 = ~(P3_ADD_546_U186 & P3_ADD_546_U185); 
assign P3_ADD_546_U121 = ~P3_ADD_546_U36; 
assign P3_ADD_546_U135 = ~P3_ADD_546_U105; 
assign P3_ADD_546_U178 = ~(P3_ADD_546_U36 & P3_EAX_REG_21__SCAN_IN); 
assign P3_ADD_546_U179 = ~(P3_ADD_546_U105 & P3_EAX_REG_20__SCAN_IN); 
assign P3_ADD_391_1180_U14 = ~(P3_U2617 & P3_ADD_391_1180_U31); 
assign P3_ADD_391_1180_U42 = ~(P3_ADD_391_1180_U31 & P3_ADD_391_1180_U13); 
assign P3_ADD_476_U90 = ~(P3_ADD_476_U180 & P3_ADD_476_U179); 
assign P3_ADD_476_U103 = ~P3_ADD_476_U24; 
assign P3_ADD_476_U177 = ~(P3_ADD_476_U24 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_531_U95 = ~(P3_ADD_531_U189 & P3_ADD_531_U188); 
assign P3_ADD_531_U107 = ~P3_ADD_531_U25; 
assign P3_ADD_531_U186 = ~(P3_ADD_531_U25 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_SUB_320_U28 = ~(P3_SUB_320_U52 & P3_SUB_320_U49 & P3_SUB_320_U86); 
assign P3_ADD_318_U90 = ~(P3_ADD_318_U180 & P3_ADD_318_U179); 
assign P3_ADD_318_U103 = ~P3_ADD_318_U24; 
assign P3_ADD_318_U177 = ~(P3_ADD_318_U24 & P3_PHYADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_315_U86 = ~(P3_ADD_315_U172 & P3_ADD_315_U171); 
assign P3_ADD_315_U100 = ~P3_ADD_315_U24; 
assign P3_ADD_315_U169 = ~(P3_ADD_315_U24 & P3_PHYADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_360_1242_U32 = ~P3_ADD_360_U18; 
assign P3_ADD_360_1242_U94 = P3_ADD_360_1242_U190 & P3_ADD_360_1242_U125; 
assign P3_ADD_360_1242_U95 = P3_ADD_360_1242_U224 & P3_ADD_360_1242_U223 & P3_ADD_360_1242_U135; 
assign P3_ADD_360_1242_U134 = ~P3_ADD_360_1242_U41; 
assign P3_ADD_360_1242_U150 = ~(P3_ADD_360_1242_U135 & P3_ADD_360_1242_U41); 
assign P3_ADD_360_1242_U152 = ~(P3_ADD_360_1242_U115 & P3_ADD_360_1242_U132); 
assign P3_ADD_360_1242_U188 = ~(P3_ADD_360_U18 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_360_1242_U191 = ~(P3_ADD_360_1242_U93 & P3_ADD_360_1242_U40); 
assign P3_ADD_360_1242_U217 = ~(P3_ADD_360_U18 & P3_ADD_360_1242_U31); 
assign P3_ADD_360_1242_U219 = ~(P3_ADD_360_U18 & P3_ADD_360_1242_U31); 
assign P3_ADD_467_U90 = ~(P3_ADD_467_U180 & P3_ADD_467_U179); 
assign P3_ADD_467_U103 = ~P3_ADD_467_U24; 
assign P3_ADD_467_U177 = ~(P3_ADD_467_U24 & P3_REIP_REG_12__SCAN_IN); 
assign P3_ADD_430_U90 = ~(P3_ADD_430_U180 & P3_ADD_430_U179); 
assign P3_ADD_430_U103 = ~P3_ADD_430_U24; 
assign P3_ADD_430_U177 = ~(P3_ADD_430_U24 & P3_REIP_REG_12__SCAN_IN); 
assign P3_ADD_380_U95 = ~(P3_ADD_380_U189 & P3_ADD_380_U188); 
assign P3_ADD_380_U107 = ~P3_ADD_380_U25; 
assign P3_ADD_380_U186 = ~(P3_ADD_380_U25 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_344_U95 = ~(P3_ADD_344_U189 & P3_ADD_344_U188); 
assign P3_ADD_344_U107 = ~P3_ADD_344_U25; 
assign P3_ADD_344_U186 = ~(P3_ADD_344_U25 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_339_U90 = ~(P3_ADD_339_U180 & P3_ADD_339_U179); 
assign P3_ADD_339_U103 = ~P3_ADD_339_U24; 
assign P3_ADD_339_U177 = ~(P3_ADD_339_U24 & P3_PHYADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_360_U5 = P3_ADD_360_U22 & P3_ADD_360_U27; 
assign P3_ADD_360_U23 = ~(P3_U2627 & P3_ADD_360_U27); 
assign P3_ADD_360_U32 = ~(P3_ADD_360_U27 & P3_ADD_360_U15); 
assign P3_ADD_541_U90 = ~(P3_ADD_541_U180 & P3_ADD_541_U179); 
assign P3_ADD_541_U103 = ~P3_ADD_541_U24; 
assign P3_ADD_541_U177 = ~(P3_ADD_541_U24 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_SUB_357_1258_U7 = P3_SUB_357_1258_U6 & P3_SUB_357_1258_U189; 
assign P3_SUB_357_1258_U8 = P3_SUB_357_1258_U5 & P3_SUB_357_1258_U190; 
assign P3_SUB_357_1258_U9 = P3_SUB_357_1258_U209 & P3_SUB_357_1258_U204; 
assign P3_SUB_357_1258_U12 = P3_SUB_357_1258_U10 & P3_SUB_357_1258_U212; 
assign P3_SUB_357_1258_U22 = ~P3_ADD_357_U9; 
assign P3_SUB_357_1258_U78 = ~(P3_SUB_357_1258_U366 & P3_SUB_357_1258_U365); 
assign P3_SUB_357_1258_U109 = P3_SUB_357_1258_U386 & P3_SUB_357_1258_U385 & P3_SUB_357_1258_U157; 
assign P3_SUB_357_1258_U110 = P3_SUB_357_1258_U232 & P3_SUB_357_1258_U153; 
assign P3_SUB_357_1258_U112 = P3_SUB_357_1258_U243 & P3_SUB_357_1258_U156; 
assign P3_SUB_357_1258_U113 = P3_SUB_357_1258_U465 & P3_SUB_357_1258_U464 & P3_SUB_357_1258_U155; 
assign P3_SUB_357_1258_U114 = P3_SUB_357_1258_U254 & P3_SUB_357_1258_U154; 
assign P3_SUB_357_1258_U116 = P3_SUB_357_1258_U314 & P3_SUB_357_1258_U313; 
assign P3_SUB_357_1258_U122 = P3_SUB_357_1258_U335 & P3_SUB_357_1258_U334; 
assign P3_SUB_357_1258_U123 = ~(P3_SUB_357_1258_U96 & P3_SUB_357_1258_U167); 
assign P3_SUB_357_1258_U126 = P3_SUB_357_1258_U356 & P3_SUB_357_1258_U355; 
assign P3_SUB_357_1258_U128 = P3_SUB_357_1258_U368 & P3_SUB_357_1258_U367; 
assign P3_SUB_357_1258_U130 = P3_SUB_357_1258_U379 & P3_SUB_357_1258_U378; 
assign P3_SUB_357_1258_U132 = P3_SUB_357_1258_U393 & P3_SUB_357_1258_U392; 
assign P3_SUB_357_1258_U134 = P3_SUB_357_1258_U400 & P3_SUB_357_1258_U399; 
assign P3_SUB_357_1258_U136 = P3_SUB_357_1258_U407 & P3_SUB_357_1258_U406; 
assign P3_SUB_357_1258_U138 = P3_SUB_357_1258_U414 & P3_SUB_357_1258_U413; 
assign P3_SUB_357_1258_U140 = P3_SUB_357_1258_U433 & P3_SUB_357_1258_U432; 
assign P3_SUB_357_1258_U142 = P3_SUB_357_1258_U444 & P3_SUB_357_1258_U443; 
assign P3_SUB_357_1258_U144 = P3_SUB_357_1258_U451 & P3_SUB_357_1258_U450; 
assign P3_SUB_357_1258_U146 = P3_SUB_357_1258_U458 & P3_SUB_357_1258_U457; 
assign P3_SUB_357_1258_U148 = P3_SUB_357_1258_U472 & P3_SUB_357_1258_U471; 
assign P3_SUB_357_1258_U175 = P3_ADD_357_U9 | P3_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P3_SUB_357_1258_U182 = ~P3_SUB_357_1258_U124; 
assign P3_SUB_357_1258_U184 = ~P3_SUB_357_1258_U125; 
assign P3_SUB_357_1258_U267 = ~(P3_ADD_357_U9 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_SUB_357_1258_U310 = ~(P3_SUB_357_1258_U309 & P3_SUB_357_1258_U308); 
assign P3_SUB_357_1258_U317 = ~(P3_SUB_357_1258_U316 & P3_SUB_357_1258_U315); 
assign P3_SUB_357_1258_U321 = ~(P3_ADD_357_U9 & P3_SUB_357_1258_U23); 
assign P3_SUB_357_1258_U323 = ~(P3_ADD_357_U9 & P3_SUB_357_1258_U23); 
assign P3_SUB_357_1258_U327 = ~(P3_SUB_357_1258_U37 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_SUB_357_1258_U329 = ~(P3_SUB_357_1258_U37 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_SUB_357_1258_U338 = ~(P3_SUB_357_1258_U337 & P3_SUB_357_1258_U336); 
assign P3_SUB_357_1258_U344 = ~(P3_SUB_357_1258_U259 & P3_SUB_357_1258_U124); 
assign P3_SUB_357_1258_U349 = ~(P3_SUB_357_1258_U260 & P3_SUB_357_1258_U125); 
assign P3_SUB_357_1258_U359 = ~(P3_SUB_357_1258_U358 & P3_SUB_357_1258_U357); 
assign P3_SUB_357_1258_U371 = ~(P3_SUB_357_1258_U370 & P3_SUB_357_1258_U369); 
assign P3_SUB_357_1258_U382 = ~(P3_SUB_357_1258_U381 & P3_SUB_357_1258_U380); 
assign P3_SUB_357_1258_U389 = ~(P3_SUB_357_1258_U388 & P3_SUB_357_1258_U387); 
assign P3_SUB_357_1258_U396 = ~(P3_SUB_357_1258_U395 & P3_SUB_357_1258_U394); 
assign P3_SUB_357_1258_U403 = ~(P3_SUB_357_1258_U402 & P3_SUB_357_1258_U401); 
assign P3_SUB_357_1258_U410 = ~(P3_SUB_357_1258_U409 & P3_SUB_357_1258_U408); 
assign P3_SUB_357_1258_U417 = ~(P3_SUB_357_1258_U416 & P3_SUB_357_1258_U415); 
assign P3_SUB_357_1258_U429 = ~(P3_SUB_357_1258_U428 & P3_SUB_357_1258_U427); 
assign P3_SUB_357_1258_U436 = ~(P3_SUB_357_1258_U435 & P3_SUB_357_1258_U434); 
assign P3_SUB_357_1258_U447 = ~(P3_SUB_357_1258_U446 & P3_SUB_357_1258_U445); 
assign P3_SUB_357_1258_U454 = ~(P3_SUB_357_1258_U453 & P3_SUB_357_1258_U452); 
assign P3_SUB_357_1258_U461 = ~(P3_SUB_357_1258_U460 & P3_SUB_357_1258_U459); 
assign P3_SUB_357_1258_U468 = ~(P3_SUB_357_1258_U467 & P3_SUB_357_1258_U466); 
assign P3_SUB_357_1258_U475 = ~(P3_SUB_357_1258_U474 & P3_SUB_357_1258_U473); 
assign P3_SUB_357_1258_U480 = ~(P3_SUB_357_1258_U479 & P3_SUB_357_1258_U478); 
assign P3_ADD_515_U90 = ~(P3_ADD_515_U180 & P3_ADD_515_U179); 
assign P3_ADD_515_U103 = ~P3_ADD_515_U24; 
assign P3_ADD_515_U177 = ~(P3_ADD_515_U24 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_394_U90 = ~(P3_ADD_394_U184 & P3_ADD_394_U183); 
assign P3_ADD_394_U106 = ~P3_ADD_394_U24; 
assign P3_ADD_394_U181 = ~(P3_ADD_394_U24 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_SUB_414_U74 = P3_SUB_414_U151 & P3_SUB_414_U150; 
assign P3_SUB_414_U98 = ~P3_SUB_414_U33; 
assign P3_SUB_414_U116 = ~(P3_SUB_414_U115 & P3_EBX_REG_20__SCAN_IN); 
assign P3_SUB_414_U146 = ~(P3_SUB_414_U33 & P3_EBX_REG_21__SCAN_IN); 
assign P3_ADD_441_U90 = ~(P3_ADD_441_U180 & P3_ADD_441_U179); 
assign P3_ADD_441_U103 = ~P3_ADD_441_U24; 
assign P3_ADD_441_U177 = ~(P3_ADD_441_U24 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_349_U95 = ~(P3_ADD_349_U189 & P3_ADD_349_U188); 
assign P3_ADD_349_U107 = ~P3_ADD_349_U25; 
assign P3_ADD_349_U186 = ~(P3_ADD_349_U25 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_405_U90 = ~(P3_ADD_405_U184 & P3_ADD_405_U183); 
assign P3_ADD_405_U106 = ~P3_ADD_405_U24; 
assign P3_ADD_405_U181 = ~(P3_ADD_405_U24 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_553_U95 = ~(P3_ADD_553_U189 & P3_ADD_553_U188); 
assign P3_ADD_553_U107 = ~P3_ADD_553_U25; 
assign P3_ADD_553_U186 = ~(P3_ADD_553_U25 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_558_U95 = ~(P3_ADD_558_U189 & P3_ADD_558_U188); 
assign P3_ADD_558_U107 = ~P3_ADD_558_U25; 
assign P3_ADD_558_U186 = ~(P3_ADD_558_U25 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_385_U95 = ~(P3_ADD_385_U189 & P3_ADD_385_U188); 
assign P3_ADD_385_U107 = ~P3_ADD_385_U25; 
assign P3_ADD_385_U186 = ~(P3_ADD_385_U25 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_547_U95 = ~(P3_ADD_547_U189 & P3_ADD_547_U188); 
assign P3_ADD_547_U107 = ~P3_ADD_547_U25; 
assign P3_ADD_547_U186 = ~(P3_ADD_547_U25 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_371_1212_U25 = ~P3_ADD_371_U19; 
assign P3_ADD_371_1212_U94 = P3_ADD_371_1212_U129 & P3_ADD_371_1212_U128; 
assign P3_ADD_371_1212_U132 = P3_ADD_371_U19 | P3_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P3_ADD_371_1212_U137 = ~(P3_ADD_371_U19 & P3_ADD_371_1212_U134); 
assign P3_ADD_371_1212_U154 = ~(P3_ADD_371_U19 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_371_1212_U159 = ~(P3_ADD_371_1212_U98 & P3_ADD_371_1212_U158); 
assign P3_ADD_371_1212_U160 = ~(P3_ADD_371_1212_U124 & P3_ADD_371_1212_U29); 
assign P3_ADD_371_1212_U228 = ~(P3_ADD_371_U19 & P3_ADD_371_1212_U23); 
assign P3_ADD_371_1212_U231 = ~(P3_ADD_371_1212_U230 & P3_ADD_371_1212_U229); 
assign P3_ADD_371_1212_U244 = ~(P3_ADD_371_1212_U242 & P3_ADD_371_1212_U124); 
assign P3_ADD_371_U6 = P3_ADD_371_U22 & P3_ADD_371_U30; 
assign P3_ADD_371_U23 = ~(P3_U2627 & P3_ADD_371_U30); 
assign P3_ADD_371_U36 = ~(P3_ADD_371_U30 & P3_ADD_371_U15); 
assign P3_ADD_494_U90 = ~(P3_ADD_494_U180 & P3_ADD_494_U179); 
assign P3_ADD_494_U103 = ~P3_ADD_494_U24; 
assign P3_ADD_494_U177 = ~(P3_ADD_494_U24 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_536_U90 = ~(P3_ADD_536_U180 & P3_ADD_536_U179); 
assign P3_ADD_536_U103 = ~P3_ADD_536_U24; 
assign P3_ADD_536_U177 = ~(P3_ADD_536_U24 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_402_1132_U14 = ~(P3_U2617 & P3_ADD_402_1132_U31); 
assign P3_ADD_402_1132_U42 = ~(P3_ADD_402_1132_U31 & P3_ADD_402_1132_U13); 
assign P2_R2099_U94 = ~(P2_R2099_U225 & P2_R2099_U224); 
assign P2_R2099_U99 = P2_R2099_U162 & P2_R2099_U161; 
assign P2_R2099_U103 = P2_R2099_U173 & P2_R2099_U172; 
assign P2_R2099_U110 = ~(P2_U2750 & P2_R2099_U109); 
assign P2_R2099_U165 = ~(P2_R2099_U164 & P2_R2099_U163); 
assign P2_R2099_U176 = ~(P2_R2099_U175 & P2_R2099_U174); 
assign P2_R2099_U200 = ~(P2_R2099_U147 & P2_R2099_U8); 
assign P2_R2099_U203 = ~(P2_R2099_U108 & P2_U2750); 
assign P2_ADD_391_1196_U23 = ~P2_R2096_U51; 
assign P2_ADD_402_1132_U14 = ~(P2_U2595 & P2_ADD_402_1132_U31); 
assign P2_ADD_402_1132_U44 = ~(P2_ADD_402_1132_U31 & P2_ADD_402_1132_U13); 
assign P2_R2182_U252 = ~(P2_U2663 & P2_R2182_U56); 
assign P2_R2182_U254 = ~(P2_U2663 & P2_R2182_U56); 
assign P2_R2167_U20 = ~(P2_U2707 & P2_R2167_U19); 
assign P2_R2027_U95 = ~(P2_R2027_U189 & P2_R2027_U188); 
assign P2_R2027_U107 = ~P2_R2027_U25; 
assign P2_R2027_U186 = ~(P2_R2027_U25 & P2_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P2_R2337_U88 = ~(P2_R2337_U178 & P2_R2337_U177); 
assign P2_R2337_U104 = ~P2_R2337_U25; 
assign P2_R2337_U175 = ~(P2_R2337_U25 & P2_PHYADDRPOINTER_REG_13__SCAN_IN); 
assign P2_R2219_U29 = ~(P2_R2219_U111 & P2_R2219_U110); 
assign P2_R2219_U41 = ~(P2_R2219_U75 & P2_R2219_U56 & P2_R2219_U74); 
assign P2_R2219_U51 = ~P2_R2219_U43; 
assign P2_R2219_U54 = ~P2_R2219_U42; 
assign P2_R2219_U101 = ~(P2_R2219_U35 & P2_R2219_U42); 
assign P2_R2219_U106 = ~(P2_R2219_U36 & P2_R2219_U43); 
assign P2_R2096_U77 = ~(P2_R2096_U218 & P2_R2096_U217); 
assign P2_R2096_U123 = ~P2_R2096_U109; 
assign P2_R2096_U125 = ~(P2_R2096_U124 & P2_R2096_U109); 
assign P2_R2096_U208 = ~(P2_R2096_U108 & P2_R2096_U109); 
assign P2_GTE_370_U9 = P2_R2219_U8 | P2_R2219_U30; 
assign P2_R1957_U27 = ~(P2_R1957_U52 & P2_R1957_U86 & P2_R1957_U48); 
assign P2_ADD_394_U73 = ~(P2_ADD_394_U148 & P2_ADD_394_U147); 
assign P2_ADD_394_U106 = ~P2_ADD_394_U24; 
assign P2_ADD_394_U179 = ~(P2_ADD_394_U24 & P2_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P2_R2267_U88 = ~P2_R2267_U77; 
assign P2_R2267_U134 = ~(P2_U2617 & P2_R2267_U22); 
assign P1_R2027_U72 = ~(P1_R2027_U184 & P1_R2027_U183); 
assign P1_R2027_U73 = ~(P1_R2027_U186 & P1_R2027_U185); 
assign P1_R2027_U121 = ~P1_R2027_U36; 
assign P1_R2027_U135 = ~P1_R2027_U105; 
assign P1_R2027_U178 = ~(P1_R2027_U36 & P1_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P1_R2027_U179 = ~(P1_R2027_U105 & P1_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P1_R2182_U21 = ~(P1_R2182_U37 & P1_R2182_U46); 
assign P1_R2182_U41 = ~(P1_R2182_U52 & P1_R2182_U53); 
assign P1_R2182_U43 = ~(P1_R2182_U46 & P1_U2736); 
assign P1_R2182_U61 = ~P1_R2182_U45; 
assign P1_R2182_U77 = ~(P1_R2182_U46 & P1_R2182_U17); 
assign P1_R2182_U80 = ~(P1_R2182_U59 & P1_R2182_U14); 
assign P1_R2182_U83 = ~(P1_R2182_U50 & P1_R2182_U45); 
assign P1_R2144_U5 = P1_R2144_U104 & P1_R2144_U103; 
assign P1_R2144_U44 = P1_R2144_U21 & P1_R2144_U105; 
assign P1_R2144_U46 = P1_R2144_U19 & P1_R2144_U106; 
assign P1_R2144_U53 = P1_R2144_U7 & P1_R2144_U52; 
assign P1_R2144_U61 = P1_R2144_U23 & P1_R2144_U81; 
assign P1_R2144_U107 = ~P1_R2144_U21; 
assign P1_R2144_U108 = ~P1_R2144_U23; 
assign P1_R2144_U120 = ~P1_R2144_U19; 
assign P1_R2144_U126 = ~(P1_R2144_U23 & P1_R2144_U81); 
assign P1_R2144_U149 = ~(P1_R2144_U21 & P1_R2144_U105); 
assign P1_R2144_U150 = ~(P1_R2144_U19 & P1_R2144_U106); 
assign P1_R2144_U156 = ~(P1_R2144_U104 & P1_R2144_U103); 
assign P1_R2358_U143 = ~P1_U2618; 
assign P1_R2358_U400 = ~(P1_U2618 & P1_R2358_U23); 
assign P1_R2358_U402 = ~(P1_U2618 & P1_R2358_U23); 
assign P1_R2358_U448 = ~(P1_R2358_U447 & P1_R2358_U446); 
assign P1_R2099_U154 = ~P1_R2099_U112; 
assign P1_R2099_U155 = ~P1_R2099_U7; 
assign P1_R2099_U223 = ~(P1_R2099_U30 & P1_R2099_U7); 
assign P1_R2099_U225 = ~(P1_R2099_U34 & P1_R2099_U112); 
assign P1_R2099_U296 = ~(P1_R2099_U153 & P1_R2099_U193); 
assign P1_R2167_U40 = ~(P1_R2167_U21 & P1_R2167_U37); 
assign P1_R2337_U90 = ~(P1_R2337_U180 & P1_R2337_U179); 
assign P1_R2337_U103 = ~P1_R2337_U24; 
assign P1_R2337_U177 = ~(P1_R2337_U24 & P1_PHYADDRPOINTER_REG_12__SCAN_IN); 
assign P1_R2096_U90 = ~(P1_R2096_U180 & P1_R2096_U179); 
assign P1_R2096_U103 = ~P1_R2096_U24; 
assign P1_R2096_U177 = ~(P1_R2096_U24 & P1_REIP_REG_12__SCAN_IN); 
assign P1_ADD_371_U17 = ~(P1_ADD_371_U34 & P1_ADD_371_U33); 
assign P1_ADD_371_U32 = ~P1_ADD_371_U25; 
assign P1_ADD_371_U43 = ~(P1_U3234 & P1_ADD_371_U25); 
assign P1_ADD_405_U73 = ~(P1_ADD_405_U148 & P1_ADD_405_U147); 
assign P1_ADD_405_U106 = ~P1_ADD_405_U24; 
assign P1_ADD_405_U179 = ~(P1_ADD_405_U24 & P1_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P1_ADD_515_U73 = ~(P1_ADD_515_U146 & P1_ADD_515_U145); 
assign P1_ADD_515_U103 = ~P1_ADD_515_U24; 
assign P1_ADD_515_U175 = ~(P1_ADD_515_U24 & P1_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_U2371 = P3_U5036 & P3_U5028; 
assign P3_U2372 = P3_U4985 & P3_U3176; 
assign P3_U2373 = P3_U4933 & P3_U3172; 
assign P3_U2374 = P3_U4881 & P3_U3168; 
assign P3_U2375 = P3_U4829 & P3_U4821; 
assign P3_U2376 = P3_U4778 & P3_U3160; 
assign P3_U2377 = P3_U4726 & P3_U3152; 
assign P3_U2378 = P3_U4674 & P3_U3146; 
assign P3_U2394 = P3_U2382 & P3_U2628; 
assign P3_U2396 = P3_U2382 & P3_U3241; 
assign P3_U2397 = P3_U2386 & P3_STATEBS16_REG_SCAN_IN; 
assign P3_U2398 = P3_U2386 & P3_U2631; 
assign P3_U2447 = P3_U2409 & P3_U3108; 
assign P3_U2604 = P3_U7947 & P3_U7946; 
assign P3_U2736 = P3_U6759 & P3_DATAO_REG_31__SCAN_IN; 
assign P3_U3230 = ~(P3_U2518 & P3_U3243); 
assign P3_U3252 = ~(P3_U2390 & P3_U6853); 
assign P3_U3260 = ~(P3_U4030 & P3_U4334); 
assign P3_U3700 = P3_U5662 & P3_U5661 & P3_U3701 & P3_U5657; 
assign P3_U4287 = ~(P3_U4151 & P3_U4334); 
assign P3_U4288 = ~(P3_U4334 & P3_U3239); 
assign P3_U4679 = ~(P3_U4672 & P3_INSTQUEUE_REG_15__7__SCAN_IN); 
assign P3_U4684 = ~(P3_U4672 & P3_INSTQUEUE_REG_15__6__SCAN_IN); 
assign P3_U4689 = ~(P3_U4672 & P3_INSTQUEUE_REG_15__5__SCAN_IN); 
assign P3_U4694 = ~(P3_U4672 & P3_INSTQUEUE_REG_15__4__SCAN_IN); 
assign P3_U4699 = ~(P3_U4672 & P3_INSTQUEUE_REG_15__3__SCAN_IN); 
assign P3_U4704 = ~(P3_U4672 & P3_INSTQUEUE_REG_15__2__SCAN_IN); 
assign P3_U4709 = ~(P3_U4672 & P3_INSTQUEUE_REG_15__1__SCAN_IN); 
assign P3_U4714 = ~(P3_U4672 & P3_INSTQUEUE_REG_15__0__SCAN_IN); 
assign P3_U4731 = ~(P3_U4724 & P3_INSTQUEUE_REG_14__7__SCAN_IN); 
assign P3_U4736 = ~(P3_U4724 & P3_INSTQUEUE_REG_14__6__SCAN_IN); 
assign P3_U4741 = ~(P3_U4724 & P3_INSTQUEUE_REG_14__5__SCAN_IN); 
assign P3_U4746 = ~(P3_U4724 & P3_INSTQUEUE_REG_14__4__SCAN_IN); 
assign P3_U4751 = ~(P3_U4724 & P3_INSTQUEUE_REG_14__3__SCAN_IN); 
assign P3_U4756 = ~(P3_U4724 & P3_INSTQUEUE_REG_14__2__SCAN_IN); 
assign P3_U4761 = ~(P3_U4724 & P3_INSTQUEUE_REG_14__1__SCAN_IN); 
assign P3_U4766 = ~(P3_U4724 & P3_INSTQUEUE_REG_14__0__SCAN_IN); 
assign P3_U4783 = ~(P3_U4776 & P3_INSTQUEUE_REG_13__7__SCAN_IN); 
assign P3_U4788 = ~(P3_U4776 & P3_INSTQUEUE_REG_13__6__SCAN_IN); 
assign P3_U4793 = ~(P3_U4776 & P3_INSTQUEUE_REG_13__5__SCAN_IN); 
assign P3_U4798 = ~(P3_U4776 & P3_INSTQUEUE_REG_13__4__SCAN_IN); 
assign P3_U4803 = ~(P3_U4776 & P3_INSTQUEUE_REG_13__3__SCAN_IN); 
assign P3_U4808 = ~(P3_U4776 & P3_INSTQUEUE_REG_13__2__SCAN_IN); 
assign P3_U4813 = ~(P3_U4776 & P3_INSTQUEUE_REG_13__1__SCAN_IN); 
assign P3_U4818 = ~(P3_U4776 & P3_INSTQUEUE_REG_13__0__SCAN_IN); 
assign P3_U4834 = ~(P3_U4827 & P3_INSTQUEUE_REG_12__7__SCAN_IN); 
assign P3_U4839 = ~(P3_U4827 & P3_INSTQUEUE_REG_12__6__SCAN_IN); 
assign P3_U4844 = ~(P3_U4827 & P3_INSTQUEUE_REG_12__5__SCAN_IN); 
assign P3_U4849 = ~(P3_U4827 & P3_INSTQUEUE_REG_12__4__SCAN_IN); 
assign P3_U4854 = ~(P3_U4827 & P3_INSTQUEUE_REG_12__3__SCAN_IN); 
assign P3_U4859 = ~(P3_U4827 & P3_INSTQUEUE_REG_12__2__SCAN_IN); 
assign P3_U4864 = ~(P3_U4827 & P3_INSTQUEUE_REG_12__1__SCAN_IN); 
assign P3_U4869 = ~(P3_U4827 & P3_INSTQUEUE_REG_12__0__SCAN_IN); 
assign P3_U4886 = ~(P3_U4879 & P3_INSTQUEUE_REG_11__7__SCAN_IN); 
assign P3_U4891 = ~(P3_U4879 & P3_INSTQUEUE_REG_11__6__SCAN_IN); 
assign P3_U4896 = ~(P3_U4879 & P3_INSTQUEUE_REG_11__5__SCAN_IN); 
assign P3_U4901 = ~(P3_U4879 & P3_INSTQUEUE_REG_11__4__SCAN_IN); 
assign P3_U4906 = ~(P3_U4879 & P3_INSTQUEUE_REG_11__3__SCAN_IN); 
assign P3_U4911 = ~(P3_U4879 & P3_INSTQUEUE_REG_11__2__SCAN_IN); 
assign P3_U4916 = ~(P3_U4879 & P3_INSTQUEUE_REG_11__1__SCAN_IN); 
assign P3_U4921 = ~(P3_U4879 & P3_INSTQUEUE_REG_11__0__SCAN_IN); 
assign P3_U4938 = ~(P3_U4931 & P3_INSTQUEUE_REG_10__7__SCAN_IN); 
assign P3_U4943 = ~(P3_U4931 & P3_INSTQUEUE_REG_10__6__SCAN_IN); 
assign P3_U4948 = ~(P3_U4931 & P3_INSTQUEUE_REG_10__5__SCAN_IN); 
assign P3_U4953 = ~(P3_U4931 & P3_INSTQUEUE_REG_10__4__SCAN_IN); 
assign P3_U4958 = ~(P3_U4931 & P3_INSTQUEUE_REG_10__3__SCAN_IN); 
assign P3_U4963 = ~(P3_U4931 & P3_INSTQUEUE_REG_10__2__SCAN_IN); 
assign P3_U4968 = ~(P3_U4931 & P3_INSTQUEUE_REG_10__1__SCAN_IN); 
assign P3_U4973 = ~(P3_U4931 & P3_INSTQUEUE_REG_10__0__SCAN_IN); 
assign P3_U4990 = ~(P3_U4983 & P3_INSTQUEUE_REG_9__7__SCAN_IN); 
assign P3_U4995 = ~(P3_U4983 & P3_INSTQUEUE_REG_9__6__SCAN_IN); 
assign P3_U5000 = ~(P3_U4983 & P3_INSTQUEUE_REG_9__5__SCAN_IN); 
assign P3_U5005 = ~(P3_U4983 & P3_INSTQUEUE_REG_9__4__SCAN_IN); 
assign P3_U5010 = ~(P3_U4983 & P3_INSTQUEUE_REG_9__3__SCAN_IN); 
assign P3_U5015 = ~(P3_U4983 & P3_INSTQUEUE_REG_9__2__SCAN_IN); 
assign P3_U5020 = ~(P3_U4983 & P3_INSTQUEUE_REG_9__1__SCAN_IN); 
assign P3_U5025 = ~(P3_U4983 & P3_INSTQUEUE_REG_9__0__SCAN_IN); 
assign P3_U5041 = ~(P3_U5034 & P3_INSTQUEUE_REG_8__7__SCAN_IN); 
assign P3_U5046 = ~(P3_U5034 & P3_INSTQUEUE_REG_8__6__SCAN_IN); 
assign P3_U5051 = ~(P3_U5034 & P3_INSTQUEUE_REG_8__5__SCAN_IN); 
assign P3_U5056 = ~(P3_U5034 & P3_INSTQUEUE_REG_8__4__SCAN_IN); 
assign P3_U5061 = ~(P3_U5034 & P3_INSTQUEUE_REG_8__3__SCAN_IN); 
assign P3_U5066 = ~(P3_U5034 & P3_INSTQUEUE_REG_8__2__SCAN_IN); 
assign P3_U5071 = ~(P3_U5034 & P3_INSTQUEUE_REG_8__1__SCAN_IN); 
assign P3_U5076 = ~(P3_U5034 & P3_INSTQUEUE_REG_8__0__SCAN_IN); 
assign P3_U5083 = ~(P3_U3510 & P3_U5081); 
assign P3_U5085 = ~(P3_U2489 & P3_U5084); 
assign P3_U5135 = ~(P3_U3528 & P3_U5133); 
assign P3_U5137 = ~(P3_U2489 & P3_U5136); 
assign P3_U5187 = ~(P3_U3546 & P3_U5185); 
assign P3_U5189 = ~(P3_U2489 & P3_U5188); 
assign P3_U5238 = ~(P3_U3564 & P3_U5236); 
assign P3_U5289 = ~(P3_U3582 & P3_U5287); 
assign P3_U5340 = ~(P3_U3599 & P3_U5338); 
assign P3_U5391 = ~(P3_U3617 & P3_U5389); 
assign P3_U5441 = ~(P3_U3635 & P3_U5439); 
assign P3_U5496 = ~P3_U4290; 
assign P3_U5497 = ~(P3_U2390 & P3_U4290); 
assign P3_U5529 = ~(P3_U2518 & P3_U3217); 
assign P3_U5539 = ~(P3_U5504 & P3_U5535); 
assign P3_U5551 = ~(P3_U5547 & P3_U5549); 
assign P3_U5590 = ~(P3_U5589 & P3_U3233); 
assign P3_U5629 = ~(P3_U2515 & P3_U5627 & P3_U3687 & P3_U5628); 
assign P3_U5652 = ~(P3_U3692 & P3_U5634 & P3_U3693 & P3_U3698); 
assign P3_U5681 = ~(P3_SUB_357_1258_U78 & P3_U2393); 
assign P3_U5874 = ~(P3_ADD_558_U95 & P3_U3220); 
assign P3_U5875 = ~(P3_ADD_553_U95 & P3_U4298); 
assign P3_U5876 = ~(P3_ADD_547_U95 & P3_U4299); 
assign P3_U5879 = ~(P3_ADD_531_U95 & P3_U2354); 
assign P3_U5887 = ~(P3_ADD_385_U95 & P3_U2358); 
assign P3_U5888 = ~(P3_ADD_380_U95 & P3_U2359); 
assign P3_U5889 = ~(P3_ADD_349_U95 & P3_U4306); 
assign P3_U5890 = ~(P3_ADD_344_U95 & P3_U2362); 
assign P3_U5901 = ~(P3_ADD_541_U90 & P3_U4300); 
assign P3_U5902 = ~(P3_ADD_536_U90 & P3_U4301); 
assign P3_U5905 = ~(P3_ADD_515_U90 & P3_U4302); 
assign P3_U5906 = ~(P3_ADD_494_U90 & P3_U2356); 
assign P3_U5907 = ~(P3_ADD_476_U90 & P3_U4303); 
assign P3_U5908 = ~(P3_ADD_441_U90 & P3_U4304); 
assign P3_U5909 = ~(P3_ADD_405_U90 & P3_U4305); 
assign P3_U5910 = ~(P3_ADD_394_U90 & P3_U2357); 
assign P3_U6072 = ~(P3_ADD_526_U73 & P3_U2355); 
assign P3_U6096 = ~(P3_ADD_526_U72 & P3_U2355); 
assign P3_U6409 = ~(P3_U2389 & P3_REIP_REG_0__SCAN_IN); 
assign P3_U6410 = ~(P3_U2388 & P3_PHYADDRPOINTER_REG_0__SCAN_IN); 
assign P3_U6411 = ~(P3_U2387 & P3_ADD_371_1212_U87); 
assign P3_U6412 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_0__SCAN_IN); 
assign P3_U6417 = ~(P3_U2389 & P3_REIP_REG_1__SCAN_IN); 
assign P3_U6418 = ~(P3_ADD_339_U4 & P3_U2388); 
assign P3_U6419 = ~(P3_U2387 & P3_ADD_371_1212_U20); 
assign P3_U6420 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_1__SCAN_IN); 
assign P3_U6425 = ~(P3_U2389 & P3_REIP_REG_2__SCAN_IN); 
assign P3_U6426 = ~(P3_ADD_339_U71 & P3_U2388); 
assign P3_U6428 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_2__SCAN_IN); 
assign P3_U6433 = ~(P3_U2389 & P3_REIP_REG_3__SCAN_IN); 
assign P3_U6434 = ~(P3_ADD_339_U68 & P3_U2388); 
assign P3_U6436 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_3__SCAN_IN); 
assign P3_U6441 = ~(P3_U2389 & P3_REIP_REG_4__SCAN_IN); 
assign P3_U6442 = ~(P3_ADD_339_U67 & P3_U2388); 
assign P3_U6444 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_4__SCAN_IN); 
assign P3_U6449 = ~(P3_U2389 & P3_REIP_REG_5__SCAN_IN); 
assign P3_U6450 = ~(P3_ADD_339_U66 & P3_U2388); 
assign P3_U6452 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_5__SCAN_IN); 
assign P3_U6457 = ~(P3_U2389 & P3_REIP_REG_6__SCAN_IN); 
assign P3_U6458 = ~(P3_ADD_339_U65 & P3_U2388); 
assign P3_U6460 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_6__SCAN_IN); 
assign P3_U6465 = ~(P3_U2389 & P3_REIP_REG_7__SCAN_IN); 
assign P3_U6466 = ~(P3_ADD_339_U64 & P3_U2388); 
assign P3_U6468 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_7__SCAN_IN); 
assign P3_U6473 = ~(P3_U2389 & P3_REIP_REG_8__SCAN_IN); 
assign P3_U6474 = ~(P3_ADD_339_U63 & P3_U2388); 
assign P3_U6476 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_8__SCAN_IN); 
assign P3_U6481 = ~(P3_U2389 & P3_REIP_REG_9__SCAN_IN); 
assign P3_U6482 = ~(P3_ADD_339_U62 & P3_U2388); 
assign P3_U6484 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_9__SCAN_IN); 
assign P3_U6489 = ~(P3_U2389 & P3_REIP_REG_10__SCAN_IN); 
assign P3_U6490 = ~(P3_ADD_339_U91 & P3_U2388); 
assign P3_U6492 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_10__SCAN_IN); 
assign P3_U6497 = ~(P3_U2389 & P3_REIP_REG_11__SCAN_IN); 
assign P3_U6498 = ~(P3_ADD_339_U90 & P3_U2388); 
assign P3_U6500 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_11__SCAN_IN); 
assign P3_U6505 = ~(P3_U2389 & P3_REIP_REG_12__SCAN_IN); 
assign P3_U6508 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_12__SCAN_IN); 
assign P3_U6513 = ~(P3_U2389 & P3_REIP_REG_13__SCAN_IN); 
assign P3_U6516 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_13__SCAN_IN); 
assign P3_U6521 = ~(P3_U2389 & P3_REIP_REG_14__SCAN_IN); 
assign P3_U6524 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_14__SCAN_IN); 
assign P3_U6529 = ~(P3_U2389 & P3_REIP_REG_15__SCAN_IN); 
assign P3_U6532 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_15__SCAN_IN); 
assign P3_U6537 = ~(P3_U2389 & P3_REIP_REG_16__SCAN_IN); 
assign P3_U6540 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_16__SCAN_IN); 
assign P3_U6545 = ~(P3_U2389 & P3_REIP_REG_17__SCAN_IN); 
assign P3_U6548 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_17__SCAN_IN); 
assign P3_U6553 = ~(P3_U2389 & P3_REIP_REG_18__SCAN_IN); 
assign P3_U6556 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_18__SCAN_IN); 
assign P3_U6561 = ~(P3_U2389 & P3_REIP_REG_19__SCAN_IN); 
assign P3_U6564 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_19__SCAN_IN); 
assign P3_U6569 = ~(P3_U2389 & P3_REIP_REG_20__SCAN_IN); 
assign P3_U6572 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_20__SCAN_IN); 
assign P3_U6577 = ~(P3_U2389 & P3_REIP_REG_21__SCAN_IN); 
assign P3_U6580 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_21__SCAN_IN); 
assign P3_U6585 = ~(P3_U2389 & P3_REIP_REG_22__SCAN_IN); 
assign P3_U6588 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_22__SCAN_IN); 
assign P3_U6593 = ~(P3_U2389 & P3_REIP_REG_23__SCAN_IN); 
assign P3_U6596 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_23__SCAN_IN); 
assign P3_U6601 = ~(P3_U2389 & P3_REIP_REG_24__SCAN_IN); 
assign P3_U6604 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_24__SCAN_IN); 
assign P3_U6609 = ~(P3_U2389 & P3_REIP_REG_25__SCAN_IN); 
assign P3_U6612 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_25__SCAN_IN); 
assign P3_U6617 = ~(P3_U2389 & P3_REIP_REG_26__SCAN_IN); 
assign P3_U6620 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_26__SCAN_IN); 
assign P3_U6625 = ~(P3_U2389 & P3_REIP_REG_27__SCAN_IN); 
assign P3_U6628 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_27__SCAN_IN); 
assign P3_U6633 = ~(P3_U2389 & P3_REIP_REG_28__SCAN_IN); 
assign P3_U6636 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_28__SCAN_IN); 
assign P3_U6641 = ~(P3_U2389 & P3_REIP_REG_29__SCAN_IN); 
assign P3_U6644 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_29__SCAN_IN); 
assign P3_U6649 = ~(P3_U2389 & P3_REIP_REG_30__SCAN_IN); 
assign P3_U6652 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_30__SCAN_IN); 
assign P3_U6657 = ~(P3_U2389 & P3_REIP_REG_31__SCAN_IN); 
assign P3_U6660 = ~(P3_U6404 & P3_PHYADDRPOINTER_REG_31__SCAN_IN); 
assign P3_U6664 = ~(P3_U2407 & P3_EAX_REG_15__SCAN_IN); 
assign P3_U6665 = ~(P3_U2406 & BUF2_REG_15__SCAN_IN); 
assign P3_U6667 = ~(P3_U2407 & P3_EAX_REG_14__SCAN_IN); 
assign P3_U6668 = ~(P3_U2406 & BUF2_REG_14__SCAN_IN); 
assign P3_U6670 = ~(P3_U2407 & P3_EAX_REG_13__SCAN_IN); 
assign P3_U6671 = ~(P3_U2406 & BUF2_REG_13__SCAN_IN); 
assign P3_U6673 = ~(P3_U2407 & P3_EAX_REG_12__SCAN_IN); 
assign P3_U6674 = ~(P3_U2406 & BUF2_REG_12__SCAN_IN); 
assign P3_U6676 = ~(P3_U2407 & P3_EAX_REG_11__SCAN_IN); 
assign P3_U6677 = ~(P3_U2406 & BUF2_REG_11__SCAN_IN); 
assign P3_U6679 = ~(P3_U2407 & P3_EAX_REG_10__SCAN_IN); 
assign P3_U6680 = ~(P3_U2406 & BUF2_REG_10__SCAN_IN); 
assign P3_U6682 = ~(P3_U2407 & P3_EAX_REG_9__SCAN_IN); 
assign P3_U6683 = ~(P3_U2406 & BUF2_REG_9__SCAN_IN); 
assign P3_U6685 = ~(P3_U2407 & P3_EAX_REG_8__SCAN_IN); 
assign P3_U6686 = ~(P3_U2406 & BUF2_REG_8__SCAN_IN); 
assign P3_U6688 = ~(P3_U2407 & P3_EAX_REG_7__SCAN_IN); 
assign P3_U6689 = ~(P3_U2406 & BUF2_REG_7__SCAN_IN); 
assign P3_U6691 = ~(P3_U2407 & P3_EAX_REG_6__SCAN_IN); 
assign P3_U6692 = ~(P3_U2406 & BUF2_REG_6__SCAN_IN); 
assign P3_U6694 = ~(P3_U2407 & P3_EAX_REG_5__SCAN_IN); 
assign P3_U6695 = ~(P3_U2406 & BUF2_REG_5__SCAN_IN); 
assign P3_U6697 = ~(P3_U2407 & P3_EAX_REG_4__SCAN_IN); 
assign P3_U6698 = ~(P3_U2406 & BUF2_REG_4__SCAN_IN); 
assign P3_U6700 = ~(P3_U2407 & P3_EAX_REG_3__SCAN_IN); 
assign P3_U6701 = ~(P3_U2406 & BUF2_REG_3__SCAN_IN); 
assign P3_U6703 = ~(P3_U2407 & P3_EAX_REG_2__SCAN_IN); 
assign P3_U6704 = ~(P3_U2406 & BUF2_REG_2__SCAN_IN); 
assign P3_U6706 = ~(P3_U2407 & P3_EAX_REG_1__SCAN_IN); 
assign P3_U6707 = ~(P3_U2406 & BUF2_REG_1__SCAN_IN); 
assign P3_U6709 = ~(P3_U2407 & P3_EAX_REG_0__SCAN_IN); 
assign P3_U6710 = ~(P3_U2406 & BUF2_REG_0__SCAN_IN); 
assign P3_U6712 = ~(P3_U2407 & P3_EAX_REG_30__SCAN_IN); 
assign P3_U6713 = ~(P3_U2406 & BUF2_REG_14__SCAN_IN); 
assign P3_U6715 = ~(P3_U2407 & P3_EAX_REG_29__SCAN_IN); 
assign P3_U6716 = ~(P3_U2406 & BUF2_REG_13__SCAN_IN); 
assign P3_U6718 = ~(P3_U2407 & P3_EAX_REG_28__SCAN_IN); 
assign P3_U6719 = ~(P3_U2406 & BUF2_REG_12__SCAN_IN); 
assign P3_U6721 = ~(P3_U2407 & P3_EAX_REG_27__SCAN_IN); 
assign P3_U6722 = ~(P3_U2406 & BUF2_REG_11__SCAN_IN); 
assign P3_U6724 = ~(P3_U2407 & P3_EAX_REG_26__SCAN_IN); 
assign P3_U6725 = ~(P3_U2406 & BUF2_REG_10__SCAN_IN); 
assign P3_U6727 = ~(P3_U2407 & P3_EAX_REG_25__SCAN_IN); 
assign P3_U6728 = ~(P3_U2406 & BUF2_REG_9__SCAN_IN); 
assign P3_U6730 = ~(P3_U2407 & P3_EAX_REG_24__SCAN_IN); 
assign P3_U6731 = ~(P3_U2406 & BUF2_REG_8__SCAN_IN); 
assign P3_U6733 = ~(P3_U2407 & P3_EAX_REG_23__SCAN_IN); 
assign P3_U6734 = ~(P3_U2406 & BUF2_REG_7__SCAN_IN); 
assign P3_U6736 = ~(P3_U2407 & P3_EAX_REG_22__SCAN_IN); 
assign P3_U6737 = ~(P3_U2406 & BUF2_REG_6__SCAN_IN); 
assign P3_U6739 = ~(P3_U2407 & P3_EAX_REG_21__SCAN_IN); 
assign P3_U6740 = ~(P3_U2406 & BUF2_REG_5__SCAN_IN); 
assign P3_U6742 = ~(P3_U2407 & P3_EAX_REG_20__SCAN_IN); 
assign P3_U6743 = ~(P3_U2406 & BUF2_REG_4__SCAN_IN); 
assign P3_U6745 = ~(P3_U2407 & P3_EAX_REG_19__SCAN_IN); 
assign P3_U6746 = ~(P3_U2406 & BUF2_REG_3__SCAN_IN); 
assign P3_U6748 = ~(P3_U2407 & P3_EAX_REG_18__SCAN_IN); 
assign P3_U6749 = ~(P3_U2406 & BUF2_REG_2__SCAN_IN); 
assign P3_U6751 = ~(P3_U2407 & P3_EAX_REG_17__SCAN_IN); 
assign P3_U6752 = ~(P3_U2406 & BUF2_REG_1__SCAN_IN); 
assign P3_U6754 = ~(P3_U2407 & P3_EAX_REG_16__SCAN_IN); 
assign P3_U6755 = ~(P3_U2406 & BUF2_REG_0__SCAN_IN); 
assign P3_U6760 = ~(P3_U2410 & P3_LWORD_REG_0__SCAN_IN); 
assign P3_U6761 = ~(P3_U2409 & P3_EAX_REG_0__SCAN_IN); 
assign P3_U6762 = ~(P3_U6759 & P3_DATAO_REG_0__SCAN_IN); 
assign P3_U6763 = ~(P3_U2410 & P3_LWORD_REG_1__SCAN_IN); 
assign P3_U6764 = ~(P3_U2409 & P3_EAX_REG_1__SCAN_IN); 
assign P3_U6765 = ~(P3_U6759 & P3_DATAO_REG_1__SCAN_IN); 
assign P3_U6766 = ~(P3_U2410 & P3_LWORD_REG_2__SCAN_IN); 
assign P3_U6767 = ~(P3_U2409 & P3_EAX_REG_2__SCAN_IN); 
assign P3_U6768 = ~(P3_U6759 & P3_DATAO_REG_2__SCAN_IN); 
assign P3_U6769 = ~(P3_U2410 & P3_LWORD_REG_3__SCAN_IN); 
assign P3_U6770 = ~(P3_U2409 & P3_EAX_REG_3__SCAN_IN); 
assign P3_U6771 = ~(P3_U6759 & P3_DATAO_REG_3__SCAN_IN); 
assign P3_U6772 = ~(P3_U2410 & P3_LWORD_REG_4__SCAN_IN); 
assign P3_U6773 = ~(P3_U2409 & P3_EAX_REG_4__SCAN_IN); 
assign P3_U6774 = ~(P3_U6759 & P3_DATAO_REG_4__SCAN_IN); 
assign P3_U6775 = ~(P3_U2410 & P3_LWORD_REG_5__SCAN_IN); 
assign P3_U6776 = ~(P3_U2409 & P3_EAX_REG_5__SCAN_IN); 
assign P3_U6777 = ~(P3_U6759 & P3_DATAO_REG_5__SCAN_IN); 
assign P3_U6778 = ~(P3_U2410 & P3_LWORD_REG_6__SCAN_IN); 
assign P3_U6779 = ~(P3_U2409 & P3_EAX_REG_6__SCAN_IN); 
assign P3_U6780 = ~(P3_U6759 & P3_DATAO_REG_6__SCAN_IN); 
assign P3_U6781 = ~(P3_U2410 & P3_LWORD_REG_7__SCAN_IN); 
assign P3_U6782 = ~(P3_U2409 & P3_EAX_REG_7__SCAN_IN); 
assign P3_U6783 = ~(P3_U6759 & P3_DATAO_REG_7__SCAN_IN); 
assign P3_U6784 = ~(P3_U2410 & P3_LWORD_REG_8__SCAN_IN); 
assign P3_U6785 = ~(P3_U2409 & P3_EAX_REG_8__SCAN_IN); 
assign P3_U6786 = ~(P3_U6759 & P3_DATAO_REG_8__SCAN_IN); 
assign P3_U6787 = ~(P3_U2410 & P3_LWORD_REG_9__SCAN_IN); 
assign P3_U6788 = ~(P3_U2409 & P3_EAX_REG_9__SCAN_IN); 
assign P3_U6789 = ~(P3_U6759 & P3_DATAO_REG_9__SCAN_IN); 
assign P3_U6790 = ~(P3_U2410 & P3_LWORD_REG_10__SCAN_IN); 
assign P3_U6791 = ~(P3_U2409 & P3_EAX_REG_10__SCAN_IN); 
assign P3_U6792 = ~(P3_U6759 & P3_DATAO_REG_10__SCAN_IN); 
assign P3_U6793 = ~(P3_U2410 & P3_LWORD_REG_11__SCAN_IN); 
assign P3_U6794 = ~(P3_U2409 & P3_EAX_REG_11__SCAN_IN); 
assign P3_U6795 = ~(P3_U6759 & P3_DATAO_REG_11__SCAN_IN); 
assign P3_U6796 = ~(P3_U2410 & P3_LWORD_REG_12__SCAN_IN); 
assign P3_U6797 = ~(P3_U2409 & P3_EAX_REG_12__SCAN_IN); 
assign P3_U6798 = ~(P3_U6759 & P3_DATAO_REG_12__SCAN_IN); 
assign P3_U6799 = ~(P3_U2410 & P3_LWORD_REG_13__SCAN_IN); 
assign P3_U6800 = ~(P3_U2409 & P3_EAX_REG_13__SCAN_IN); 
assign P3_U6801 = ~(P3_U6759 & P3_DATAO_REG_13__SCAN_IN); 
assign P3_U6802 = ~(P3_U2410 & P3_LWORD_REG_14__SCAN_IN); 
assign P3_U6803 = ~(P3_U2409 & P3_EAX_REG_14__SCAN_IN); 
assign P3_U6804 = ~(P3_U6759 & P3_DATAO_REG_14__SCAN_IN); 
assign P3_U6805 = ~(P3_U2410 & P3_LWORD_REG_15__SCAN_IN); 
assign P3_U6806 = ~(P3_U2409 & P3_EAX_REG_15__SCAN_IN); 
assign P3_U6807 = ~(P3_U6759 & P3_DATAO_REG_15__SCAN_IN); 
assign P3_U6809 = ~(P3_U2410 & P3_UWORD_REG_0__SCAN_IN); 
assign P3_U6810 = ~(P3_U6759 & P3_DATAO_REG_16__SCAN_IN); 
assign P3_U6812 = ~(P3_U2410 & P3_UWORD_REG_1__SCAN_IN); 
assign P3_U6813 = ~(P3_U6759 & P3_DATAO_REG_17__SCAN_IN); 
assign P3_U6815 = ~(P3_U2410 & P3_UWORD_REG_2__SCAN_IN); 
assign P3_U6816 = ~(P3_U6759 & P3_DATAO_REG_18__SCAN_IN); 
assign P3_U6818 = ~(P3_U2410 & P3_UWORD_REG_3__SCAN_IN); 
assign P3_U6819 = ~(P3_U6759 & P3_DATAO_REG_19__SCAN_IN); 
assign P3_U6821 = ~(P3_U2410 & P3_UWORD_REG_4__SCAN_IN); 
assign P3_U6822 = ~(P3_U6759 & P3_DATAO_REG_20__SCAN_IN); 
assign P3_U6824 = ~(P3_U2410 & P3_UWORD_REG_5__SCAN_IN); 
assign P3_U6825 = ~(P3_U6759 & P3_DATAO_REG_21__SCAN_IN); 
assign P3_U6827 = ~(P3_U2410 & P3_UWORD_REG_6__SCAN_IN); 
assign P3_U6828 = ~(P3_U6759 & P3_DATAO_REG_22__SCAN_IN); 
assign P3_U6830 = ~(P3_U2410 & P3_UWORD_REG_7__SCAN_IN); 
assign P3_U6831 = ~(P3_U6759 & P3_DATAO_REG_23__SCAN_IN); 
assign P3_U6833 = ~(P3_U2410 & P3_UWORD_REG_8__SCAN_IN); 
assign P3_U6834 = ~(P3_U6759 & P3_DATAO_REG_24__SCAN_IN); 
assign P3_U6836 = ~(P3_U2410 & P3_UWORD_REG_9__SCAN_IN); 
assign P3_U6837 = ~(P3_U6759 & P3_DATAO_REG_25__SCAN_IN); 
assign P3_U6839 = ~(P3_U2410 & P3_UWORD_REG_10__SCAN_IN); 
assign P3_U6840 = ~(P3_U6759 & P3_DATAO_REG_26__SCAN_IN); 
assign P3_U6842 = ~(P3_U2410 & P3_UWORD_REG_11__SCAN_IN); 
assign P3_U6843 = ~(P3_U6759 & P3_DATAO_REG_27__SCAN_IN); 
assign P3_U6845 = ~(P3_U2410 & P3_UWORD_REG_12__SCAN_IN); 
assign P3_U6846 = ~(P3_U6759 & P3_DATAO_REG_28__SCAN_IN); 
assign P3_U6848 = ~(P3_U2410 & P3_UWORD_REG_13__SCAN_IN); 
assign P3_U6849 = ~(P3_U6759 & P3_DATAO_REG_29__SCAN_IN); 
assign P3_U6851 = ~(P3_U2410 & P3_UWORD_REG_14__SCAN_IN); 
assign P3_U6852 = ~(P3_U6759 & P3_DATAO_REG_30__SCAN_IN); 
assign P3_U6998 = ~(P3_U2408 & P3_INSTQUEUE_REG_0__0__SCAN_IN); 
assign P3_U6999 = ~(P3_ADD_552_U5 & P3_U2399); 
assign P3_U7001 = ~(P3_U2408 & P3_INSTQUEUE_REG_0__1__SCAN_IN); 
assign P3_U7002 = ~(P3_ADD_552_U71 & P3_U2399); 
assign P3_U7004 = ~(P3_U2408 & P3_INSTQUEUE_REG_0__2__SCAN_IN); 
assign P3_U7005 = ~(P3_ADD_552_U60 & P3_U2399); 
assign P3_U7007 = ~(P3_U2408 & P3_INSTQUEUE_REG_0__3__SCAN_IN); 
assign P3_U7008 = ~(P3_ADD_552_U57 & P3_U2399); 
assign P3_U7010 = ~(P3_U2408 & P3_INSTQUEUE_REG_0__4__SCAN_IN); 
assign P3_U7011 = ~(P3_ADD_552_U56 & P3_U2399); 
assign P3_U7013 = ~(P3_U2408 & P3_INSTQUEUE_REG_0__5__SCAN_IN); 
assign P3_U7014 = ~(P3_ADD_552_U55 & P3_U2399); 
assign P3_U7016 = ~(P3_U2408 & P3_INSTQUEUE_REG_0__6__SCAN_IN); 
assign P3_U7017 = ~(P3_ADD_552_U54 & P3_U2399); 
assign P3_U7019 = ~(P3_U2408 & P3_INSTQUEUE_REG_0__7__SCAN_IN); 
assign P3_U7020 = ~(P3_ADD_552_U53 & P3_U2399); 
assign P3_U7022 = ~(P3_U2605 & P3_U2408); 
assign P3_U7023 = ~(P3_ADD_552_U52 & P3_U2399); 
assign P3_U7025 = ~(P3_U2606 & P3_U2408); 
assign P3_U7026 = ~(P3_ADD_552_U51 & P3_U2399); 
assign P3_U7028 = ~(P3_U2607 & P3_U2408); 
assign P3_U7029 = ~(P3_ADD_552_U81 & P3_U2399); 
assign P3_U7031 = ~(P3_U2608 & P3_U2408); 
assign P3_U7032 = ~(P3_ADD_552_U80 & P3_U2399); 
assign P3_U7034 = ~(P3_U2609 & P3_U2408); 
assign P3_U7035 = ~(P3_ADD_552_U79 & P3_U2399); 
assign P3_U7037 = ~(P3_U2610 & P3_U2408); 
assign P3_U7038 = ~(P3_ADD_552_U78 & P3_U2399); 
assign P3_U7040 = ~(P3_U2611 & P3_U2408); 
assign P3_U7041 = ~(P3_ADD_552_U77 & P3_U2399); 
assign P3_U7043 = ~(P3_U2612 & P3_U2408); 
assign P3_U7044 = ~(P3_ADD_552_U76 & P3_U2399); 
assign P3_U7046 = ~(P3_U3062 & P3_U2408); 
assign P3_U7047 = ~(P3_ADD_552_U75 & P3_U2399); 
assign P3_U7049 = ~(P3_U3063 & P3_U2408); 
assign P3_U7050 = ~(P3_ADD_552_U74 & P3_U2399); 
assign P3_U7052 = ~(P3_U3064 & P3_U2408); 
assign P3_U7053 = ~(P3_ADD_552_U73 & P3_U2399); 
assign P3_U7055 = ~(P3_U3065 & P3_U2408); 
assign P3_U7056 = ~(P3_ADD_552_U72 & P3_U2399); 
assign P3_U7058 = ~(P3_U3066 & P3_U2408); 
assign P3_U7061 = ~(P3_U3067 & P3_U2408); 
assign P3_U7064 = ~(P3_U3068 & P3_U2408); 
assign P3_U7067 = ~(P3_ADD_402_1132_U25 & P3_U2408); 
assign P3_U7070 = ~(P3_ADD_402_1132_U24 & P3_U2408); 
assign P3_U7073 = ~(P3_ADD_402_1132_U23 & P3_U2408); 
assign P3_U7076 = ~(P3_ADD_402_1132_U22 & P3_U2408); 
assign P3_U7370 = ~(P3_U4623 & P3_U2390); 
assign P3_U8044 = ~(P3_U3303 & P3_U4290); 
assign P2_U2394 = P2_U4442 & P2_U2616; 
assign P2_U2395 = P2_U4442 & P2_U7873; 
assign P2_U2713 = ~(P2_U7725 & P2_STATE2_REG_0__SCAN_IN); 
assign P2_U3323 = ~P2_R2099_U94; 
assign P2_U3645 = ~(P2_U8344 & P2_U8343); 
assign P2_U4407 = ~P2_R2219_U29; 
assign P2_U5636 = ~(P2_R2099_U94 & P2_U5603); 
assign P2_U5654 = ~(P2_R2096_U77 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U7163 = ~(P2_U4467 & P2_R2099_U94); 
assign P2_U8341 = ~(P2_R2219_U29 & P2_U2617); 
assign P2_U8413 = ~(P2_R2337_U88 & P2_U3284); 
assign P1_U2610 = ~(P1_U6856 & P1_U4026); 
assign P1_U2672 = ~(P1_U6866 & P1_U6864 & P1_U6865 & P1_U6868 & P1_U6867); 
assign P1_U2768 = ~(P1_U7046 & P1_U7044 & P1_U7045); 
assign P1_U5531 = ~(P1_U4175 & P1_U5530); 
assign P1_U6855 = ~(P1_R2337_U90 & P1_U2352); 
assign P1_U6876 = ~(P1_ADD_371_U17 & P1_U4208); 
assign P3_ADD_526_U40 = ~(P3_ADD_526_U91 & P3_ADD_526_U121); 
assign P3_ADD_526_U104 = ~(P3_ADD_526_U121 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_526_U177 = ~(P3_ADD_526_U121 & P3_ADD_526_U35); 
assign P3_ADD_526_U180 = ~(P3_ADD_526_U135 & P3_ADD_526_U32); 
assign P3_ADD_552_U40 = ~(P3_ADD_552_U91 & P3_ADD_552_U121); 
assign P3_ADD_552_U104 = ~(P3_ADD_552_U121 & P3_EBX_REG_21__SCAN_IN); 
assign P3_ADD_552_U177 = ~(P3_ADD_552_U121 & P3_ADD_552_U35); 
assign P3_ADD_552_U180 = ~(P3_ADD_552_U135 & P3_ADD_552_U32); 
assign P3_ADD_546_U40 = ~(P3_ADD_546_U91 & P3_ADD_546_U121); 
assign P3_ADD_546_U104 = ~(P3_ADD_546_U121 & P3_EAX_REG_21__SCAN_IN); 
assign P3_ADD_546_U177 = ~(P3_ADD_546_U121 & P3_ADD_546_U35); 
assign P3_ADD_546_U180 = ~(P3_ADD_546_U135 & P3_ADD_546_U32); 
assign P3_ADD_391_1180_U21 = ~(P3_ADD_391_1180_U42 & P3_ADD_391_1180_U41); 
assign P3_ADD_391_1180_U32 = ~P3_ADD_391_1180_U14; 
assign P3_ADD_391_1180_U39 = ~(P3_U2618 & P3_ADD_391_1180_U14); 
assign P3_ADD_476_U26 = ~(P3_ADD_476_U103 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_476_U178 = ~(P3_ADD_476_U103 & P3_ADD_476_U25); 
assign P3_ADD_531_U27 = ~(P3_ADD_531_U107 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_531_U187 = ~(P3_ADD_531_U107 & P3_ADD_531_U26); 
assign P3_SUB_320_U6 = P3_SUB_320_U126 & P3_SUB_320_U28; 
assign P3_SUB_320_U81 = ~P3_ADD_318_U90; 
assign P3_SUB_320_U93 = ~P3_SUB_320_U28; 
assign P3_SUB_320_U158 = ~(P3_ADD_318_U90 & P3_SUB_320_U28); 
assign P3_ADD_318_U26 = ~(P3_ADD_318_U103 & P3_PHYADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_318_U178 = ~(P3_ADD_318_U103 & P3_ADD_318_U25); 
assign P3_ADD_315_U26 = ~(P3_ADD_315_U100 & P3_PHYADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_315_U170 = ~(P3_ADD_315_U100 & P3_ADD_315_U25); 
assign P3_ADD_360_1242_U37 = ~P3_ADD_360_U5; 
assign P3_ADD_360_1242_U114 = ~(P3_ADD_360_1242_U94 & P3_ADD_360_1242_U191); 
assign P3_ADD_360_1242_U145 = P3_ADD_360_U5 | P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_360_1242_U147 = ~(P3_ADD_360_U5 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_360_1242_U149 = ~(P3_ADD_360_1242_U95 & P3_ADD_360_1242_U41); 
assign P3_ADD_360_1242_U151 = ~(P3_ADD_360_1242_U96 & P3_ADD_360_1242_U150); 
assign P3_ADD_360_1242_U153 = ~(P3_ADD_360_1242_U134 & P3_ADD_360_1242_U135); 
assign P3_ADD_360_1242_U196 = ~(P3_ADD_360_U5 & P3_ADD_360_1242_U38); 
assign P3_ADD_360_1242_U198 = ~(P3_ADD_360_U5 & P3_ADD_360_1242_U38); 
assign P3_ADD_360_1242_U216 = ~(P3_ADD_360_1242_U32 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_360_1242_U218 = ~(P3_ADD_360_1242_U32 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_467_U26 = ~(P3_ADD_467_U103 & P3_REIP_REG_12__SCAN_IN); 
assign P3_ADD_467_U178 = ~(P3_ADD_467_U103 & P3_ADD_467_U25); 
assign P3_ADD_430_U26 = ~(P3_ADD_430_U103 & P3_REIP_REG_12__SCAN_IN); 
assign P3_ADD_430_U178 = ~(P3_ADD_430_U103 & P3_ADD_430_U25); 
assign P3_ADD_380_U27 = ~(P3_ADD_380_U107 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_380_U187 = ~(P3_ADD_380_U107 & P3_ADD_380_U26); 
assign P3_ADD_344_U27 = ~(P3_ADD_344_U107 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_344_U187 = ~(P3_ADD_344_U107 & P3_ADD_344_U26); 
assign P3_ADD_339_U26 = ~(P3_ADD_339_U103 & P3_PHYADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_339_U178 = ~(P3_ADD_339_U103 & P3_ADD_339_U25); 
assign P3_ADD_360_U17 = ~(P3_ADD_360_U32 & P3_ADD_360_U31); 
assign P3_ADD_360_U28 = ~P3_ADD_360_U23; 
assign P3_ADD_360_U29 = ~(P3_U2628 & P3_ADD_360_U23); 
assign P3_ADD_541_U26 = ~(P3_ADD_541_U103 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_541_U178 = ~(P3_ADD_541_U103 & P3_ADD_541_U25); 
assign P3_SUB_357_1258_U11 = P3_SUB_357_1258_U9 & P3_SUB_357_1258_U211; 
assign P3_SUB_357_1258_U14 = P3_SUB_357_1258_U12 & P3_SUB_357_1258_U214; 
assign P3_SUB_357_1258_U98 = P3_SUB_357_1258_U7 & P3_SUB_357_1258_U154; 
assign P3_SUB_357_1258_U100 = P3_SUB_357_1258_U99 & P3_SUB_357_1258_U8; 
assign P3_SUB_357_1258_U120 = P3_SUB_357_1258_U328 & P3_SUB_357_1258_U327; 
assign P3_SUB_357_1258_U169 = ~P3_SUB_357_1258_U123; 
assign P3_SUB_357_1258_U298 = ~(P3_SUB_357_1258_U170 & P3_SUB_357_1258_U123); 
assign P3_SUB_357_1258_U320 = ~(P3_SUB_357_1258_U22 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_SUB_357_1258_U322 = ~(P3_SUB_357_1258_U22 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_SUB_357_1258_U331 = ~(P3_SUB_357_1258_U330 & P3_SUB_357_1258_U329); 
assign P3_SUB_357_1258_U339 = ~(P3_SUB_357_1258_U122 & P3_SUB_357_1258_U123); 
assign P3_SUB_357_1258_U345 = ~(P3_SUB_357_1258_U182 & P3_SUB_357_1258_U343); 
assign P3_SUB_357_1258_U350 = ~(P3_SUB_357_1258_U184 & P3_SUB_357_1258_U348); 
assign P3_ADD_515_U26 = ~(P3_ADD_515_U103 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_515_U178 = ~(P3_ADD_515_U103 & P3_ADD_515_U25); 
assign P3_ADD_394_U26 = ~(P3_ADD_394_U106 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_394_U182 = ~(P3_ADD_394_U106 & P3_ADD_394_U25); 
assign P3_SUB_414_U11 = P3_SUB_414_U116 & P3_SUB_414_U33; 
assign P3_SUB_414_U34 = ~(P3_SUB_414_U43 & P3_SUB_414_U69 & P3_SUB_414_U98); 
assign P3_SUB_414_U113 = ~(P3_SUB_414_U98 & P3_SUB_414_U69); 
assign P3_SUB_414_U147 = ~(P3_SUB_414_U98 & P3_SUB_414_U69); 
assign P3_ADD_441_U26 = ~(P3_ADD_441_U103 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_441_U178 = ~(P3_ADD_441_U103 & P3_ADD_441_U25); 
assign P3_ADD_349_U27 = ~(P3_ADD_349_U107 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_349_U187 = ~(P3_ADD_349_U107 & P3_ADD_349_U26); 
assign P3_ADD_405_U26 = ~(P3_ADD_405_U106 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_405_U182 = ~(P3_ADD_405_U106 & P3_ADD_405_U25); 
assign P3_ADD_553_U27 = ~(P3_ADD_553_U107 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_553_U187 = ~(P3_ADD_553_U107 & P3_ADD_553_U26); 
assign P3_ADD_558_U27 = ~(P3_ADD_558_U107 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_558_U187 = ~(P3_ADD_558_U107 & P3_ADD_558_U26); 
assign P3_ADD_385_U27 = ~(P3_ADD_385_U107 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_385_U187 = ~(P3_ADD_385_U107 & P3_ADD_385_U26); 
assign P3_ADD_547_U27 = ~(P3_ADD_547_U107 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_547_U187 = ~(P3_ADD_547_U107 & P3_ADD_547_U26); 
assign P3_ADD_371_1212_U4 = P3_ADD_371_1212_U133 & P3_ADD_371_1212_U132; 
assign P3_ADD_371_1212_U40 = ~P3_ADD_371_U6; 
assign P3_ADD_371_1212_U43 = ~(P3_ADD_371_1212_U94 & P3_ADD_371_1212_U130); 
assign P3_ADD_371_1212_U93 = ~(P3_ADD_371_1212_U244 & P3_ADD_371_1212_U243); 
assign P3_ADD_371_1212_U135 = ~(P3_ADD_371_1212_U25 & P3_ADD_371_1212_U24); 
assign P3_ADD_371_1212_U146 = P3_ADD_371_U6 | P3_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P3_ADD_371_1212_U148 = ~(P3_ADD_371_U6 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_371_1212_U162 = ~(P3_ADD_371_1212_U160 & P3_ADD_371_1212_U161 & P3_ADD_371_1212_U119); 
assign P3_ADD_371_1212_U207 = ~(P3_ADD_371_U6 & P3_ADD_371_1212_U41); 
assign P3_ADD_371_1212_U209 = ~(P3_ADD_371_U6 & P3_ADD_371_1212_U41); 
assign P3_ADD_371_1212_U227 = ~(P3_ADD_371_1212_U25 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_371_U18 = ~(P3_ADD_371_U36 & P3_ADD_371_U35); 
assign P3_ADD_371_U31 = ~P3_ADD_371_U23; 
assign P3_ADD_371_U33 = ~(P3_U2628 & P3_ADD_371_U23); 
assign P3_ADD_494_U26 = ~(P3_ADD_494_U103 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_494_U178 = ~(P3_ADD_494_U103 & P3_ADD_494_U25); 
assign P3_ADD_536_U26 = ~(P3_ADD_536_U103 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_536_U178 = ~(P3_ADD_536_U103 & P3_ADD_536_U25); 
assign P3_ADD_402_1132_U21 = ~(P3_ADD_402_1132_U42 & P3_ADD_402_1132_U41); 
assign P3_ADD_402_1132_U32 = ~P3_ADD_402_1132_U14; 
assign P3_ADD_402_1132_U39 = ~(P3_U2618 & P3_ADD_402_1132_U14); 
assign P2_R2099_U104 = ~(P2_R2099_U106 & P2_R2099_U110); 
assign P2_R2099_U107 = P2_R2099_U203 & P2_R2099_U202; 
assign P2_R2099_U201 = ~(P2_R2099_U200 & P2_R2099_U199); 
assign P2_ADD_391_1196_U25 = ~P2_R2096_U77; 
assign P2_ADD_402_1132_U22 = ~(P2_ADD_402_1132_U44 & P2_ADD_402_1132_U43); 
assign P2_ADD_402_1132_U32 = ~P2_ADD_402_1132_U14; 
assign P2_ADD_402_1132_U47 = ~(P2_U2596 & P2_ADD_402_1132_U14); 
assign P2_R2182_U58 = ~P2_U2686; 
assign P2_R2182_U116 = P2_R2182_U253 & P2_R2182_U252; 
assign P2_R2182_U167 = P2_U2686 | P2_U2662; 
assign P2_R2182_U169 = ~(P2_U2662 & P2_U2686); 
assign P2_R2182_U246 = ~(P2_U2686 & P2_R2182_U59); 
assign P2_R2182_U248 = ~(P2_U2686 & P2_R2182_U59); 
assign P2_R2182_U256 = ~(P2_R2182_U255 & P2_R2182_U254); 
assign P2_R2027_U27 = ~(P2_R2027_U107 & P2_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P2_R2027_U187 = ~(P2_R2027_U107 & P2_R2027_U26); 
assign P2_R2337_U27 = ~(P2_R2337_U104 & P2_PHYADDRPOINTER_REG_13__SCAN_IN); 
assign P2_R2337_U176 = ~(P2_R2337_U104 & P2_R2337_U26); 
assign P2_R2219_U57 = ~P2_R2219_U41; 
assign P2_R2219_U59 = ~(P2_R2219_U58 & P2_R2219_U41); 
assign P2_R2219_U96 = ~(P2_R2219_U34 & P2_R2219_U41); 
assign P2_R2219_U100 = ~(P2_R2219_U54 & P2_R2219_U99); 
assign P2_R2219_U105 = ~(P2_R2219_U51 & P2_R2219_U104); 
assign P2_R2096_U107 = ~(P2_R2096_U126 & P2_R2096_U125); 
assign P2_R2096_U209 = ~(P2_R2096_U123 & P2_R2096_U207); 
assign P2_GTE_370_U7 = P2_R2219_U29 & P2_GTE_370_U9; 
assign P2_R1957_U6 = P2_R1957_U126 & P2_R1957_U27; 
assign P2_R1957_U81 = ~P2_U3680; 
assign P2_R1957_U93 = ~P2_R1957_U27; 
assign P2_R1957_U158 = ~(P2_U3680 & P2_R1957_U27); 
assign P2_ADD_394_U26 = ~(P2_ADD_394_U106 & P2_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P2_ADD_394_U180 = ~(P2_ADD_394_U106 & P2_ADD_394_U25); 
assign P2_R2267_U21 = ~(P2_R2267_U77 & P2_R2267_U134); 
assign P1_R2027_U40 = ~(P1_R2027_U91 & P1_R2027_U121); 
assign P1_R2027_U104 = ~(P1_R2027_U121 & P1_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P1_R2027_U177 = ~(P1_R2027_U121 & P1_R2027_U35); 
assign P1_R2027_U180 = ~(P1_R2027_U135 & P1_R2027_U32); 
assign P1_R2182_U13 = ~(P1_R2182_U35 & P1_R2182_U41); 
assign P1_R2182_U30 = ~(P1_R2182_U78 & P1_R2182_U77); 
assign P1_R2182_U31 = ~(P1_R2182_U80 & P1_R2182_U79); 
assign P1_R2182_U38 = ~(P1_U2742 & P1_R2182_U41); 
assign P1_R2182_U48 = ~P1_R2182_U21; 
assign P1_R2182_U54 = ~P1_R2182_U41; 
assign P1_R2182_U58 = ~P1_R2182_U43; 
assign P1_R2182_U69 = ~(P1_U2742 & P1_R2182_U41); 
assign P1_R2182_U74 = ~(P1_U2734 & P1_R2182_U21); 
assign P1_R2182_U75 = ~(P1_U2735 & P1_R2182_U43); 
assign P1_R2182_U84 = ~(P1_R2182_U61 & P1_R2182_U9); 
assign P1_R2144_U57 = P1_R2144_U156 & P1_R2144_U21; 
assign P1_R2144_U59 = P1_R2144_U5 & P1_R2144_U105; 
assign P1_R2144_U60 = P1_R2144_U126 & P1_R2144_U21; 
assign P1_R2144_U151 = ~(P1_R2144_U120 & P1_R2144_U105 & P1_R2144_U7); 
assign P1_R2144_U152 = ~(P1_R2144_U107 & P1_R2144_U7); 
assign P1_R2144_U153 = ~(P1_R2144_U108 & P1_R2144_U7); 
assign P1_R2144_U213 = ~(P1_R2144_U5 & P1_R2144_U108); 
assign P1_R2144_U214 = ~(P1_R2144_U102 & P1_R2144_U156); 
assign P1_R2358_U399 = ~(P1_U2352 & P1_R2358_U143); 
assign P1_R2358_U401 = ~(P1_U2352 & P1_R2358_U143); 
assign P1_R2099_U8 = ~(P1_R2099_U89 & P1_R2099_U155); 
assign P1_R2099_U111 = ~(P1_R2099_U155 & P1_R2099_U30); 
assign P1_R2099_U138 = P1_R2099_U297 & P1_R2099_U296; 
assign P1_R2099_U222 = ~(P1_R2099_U199 & P1_R2099_U155); 
assign P1_R2099_U224 = ~(P1_R2099_U154 & P1_R2099_U196); 
assign P1_R2167_U42 = ~(P1_R2167_U40 & P1_R2167_U41); 
assign P1_R2337_U26 = ~(P1_R2337_U103 & P1_PHYADDRPOINTER_REG_12__SCAN_IN); 
assign P1_R2337_U178 = ~(P1_R2337_U103 & P1_R2337_U25); 
assign P1_R2096_U26 = ~(P1_R2096_U103 & P1_REIP_REG_12__SCAN_IN); 
assign P1_R2096_U178 = ~(P1_R2096_U103 & P1_R2096_U25); 
assign P1_ADD_371_U44 = ~(P1_ADD_371_U32 & P1_ADD_371_U16); 
assign P1_ADD_405_U26 = ~(P1_ADD_405_U106 & P1_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P1_ADD_405_U180 = ~(P1_ADD_405_U106 & P1_ADD_405_U25); 
assign P1_ADD_515_U26 = ~(P1_ADD_515_U103 & P1_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P1_ADD_515_U176 = ~(P1_ADD_515_U103 & P1_ADD_515_U25); 
assign P3_U2368 = P3_U5189 & P3_U3193; 
assign P3_U2369 = P3_U5137 & P3_U3189; 
assign P3_U2370 = P3_U5085 & P3_U3185; 
assign P3_U2380 = P3_U3260 & P3_STATE2_REG_2__SCAN_IN; 
assign P3_U2385 = P3_U3260 & P3_STATE2_REG_1__SCAN_IN; 
assign P3_U2401 = P3_U3260 & P3_STATE2_REG_3__SCAN_IN; 
assign P3_U2684 = ~(P3_U7057 & P3_U7055 & P3_U7056); 
assign P3_U2685 = ~(P3_U7054 & P3_U7052 & P3_U7053); 
assign P3_U2686 = ~(P3_U7051 & P3_U7049 & P3_U7050); 
assign P3_U2687 = ~(P3_U7048 & P3_U7046 & P3_U7047); 
assign P3_U2688 = ~(P3_U7045 & P3_U7043 & P3_U7044); 
assign P3_U2689 = ~(P3_U7042 & P3_U7040 & P3_U7041); 
assign P3_U2690 = ~(P3_U7039 & P3_U7037 & P3_U7038); 
assign P3_U2691 = ~(P3_U7036 & P3_U7034 & P3_U7035); 
assign P3_U2692 = ~(P3_U7033 & P3_U7031 & P3_U7032); 
assign P3_U2693 = ~(P3_U7030 & P3_U7028 & P3_U7029); 
assign P3_U2694 = ~(P3_U7026 & P3_U7025 & P3_U7027); 
assign P3_U2695 = ~(P3_U7023 & P3_U7022 & P3_U7024); 
assign P3_U2696 = ~(P3_U7020 & P3_U7019 & P3_U7021); 
assign P3_U2697 = ~(P3_U7017 & P3_U7016 & P3_U7018); 
assign P3_U2698 = ~(P3_U7014 & P3_U7013 & P3_U7015); 
assign P3_U2699 = ~(P3_U7011 & P3_U7010 & P3_U7012); 
assign P3_U2700 = ~(P3_U7008 & P3_U7007 & P3_U7009); 
assign P3_U2701 = ~(P3_U7005 & P3_U7004 & P3_U7006); 
assign P3_U2702 = ~(P3_U7002 & P3_U7001 & P3_U7003); 
assign P3_U2703 = ~(P3_U6999 & P3_U6998 & P3_U7000); 
assign P3_U2752 = ~(P3_U6806 & P3_U6805 & P3_U6807); 
assign P3_U2753 = ~(P3_U6803 & P3_U6802 & P3_U6804); 
assign P3_U2754 = ~(P3_U6800 & P3_U6799 & P3_U6801); 
assign P3_U2755 = ~(P3_U6797 & P3_U6796 & P3_U6798); 
assign P3_U2756 = ~(P3_U6794 & P3_U6793 & P3_U6795); 
assign P3_U2757 = ~(P3_U6791 & P3_U6790 & P3_U6792); 
assign P3_U2758 = ~(P3_U6788 & P3_U6787 & P3_U6789); 
assign P3_U2759 = ~(P3_U6785 & P3_U6784 & P3_U6786); 
assign P3_U2760 = ~(P3_U6782 & P3_U6781 & P3_U6783); 
assign P3_U2761 = ~(P3_U6779 & P3_U6778 & P3_U6780); 
assign P3_U2762 = ~(P3_U6776 & P3_U6775 & P3_U6777); 
assign P3_U2763 = ~(P3_U6773 & P3_U6772 & P3_U6774); 
assign P3_U2764 = ~(P3_U6770 & P3_U6769 & P3_U6771); 
assign P3_U2765 = ~(P3_U6767 & P3_U6766 & P3_U6768); 
assign P3_U2766 = ~(P3_U6764 & P3_U6763 & P3_U6765); 
assign P3_U2767 = ~(P3_U6761 & P3_U6760 & P3_U6762); 
assign P3_U2768 = ~(P3_U6755 & P3_U6754 & P3_U6756); 
assign P3_U2769 = ~(P3_U6752 & P3_U6751 & P3_U6753); 
assign P3_U2770 = ~(P3_U6749 & P3_U6748 & P3_U6750); 
assign P3_U2771 = ~(P3_U6746 & P3_U6745 & P3_U6747); 
assign P3_U2772 = ~(P3_U6743 & P3_U6742 & P3_U6744); 
assign P3_U2773 = ~(P3_U6740 & P3_U6739 & P3_U6741); 
assign P3_U2774 = ~(P3_U6737 & P3_U6736 & P3_U6738); 
assign P3_U2775 = ~(P3_U6734 & P3_U6733 & P3_U6735); 
assign P3_U2776 = ~(P3_U6731 & P3_U6730 & P3_U6732); 
assign P3_U2777 = ~(P3_U6728 & P3_U6727 & P3_U6729); 
assign P3_U2778 = ~(P3_U6725 & P3_U6724 & P3_U6726); 
assign P3_U2779 = ~(P3_U6722 & P3_U6721 & P3_U6723); 
assign P3_U2780 = ~(P3_U6719 & P3_U6718 & P3_U6720); 
assign P3_U2781 = ~(P3_U6716 & P3_U6715 & P3_U6717); 
assign P3_U2782 = ~(P3_U6713 & P3_U6712 & P3_U6714); 
assign P3_U2783 = ~(P3_U6710 & P3_U6709 & P3_U6711); 
assign P3_U2784 = ~(P3_U6707 & P3_U6706 & P3_U6708); 
assign P3_U2785 = ~(P3_U6704 & P3_U6703 & P3_U6705); 
assign P3_U2786 = ~(P3_U6701 & P3_U6700 & P3_U6702); 
assign P3_U2787 = ~(P3_U6698 & P3_U6697 & P3_U6699); 
assign P3_U2788 = ~(P3_U6695 & P3_U6694 & P3_U6696); 
assign P3_U2789 = ~(P3_U6692 & P3_U6691 & P3_U6693); 
assign P3_U2790 = ~(P3_U6689 & P3_U6688 & P3_U6690); 
assign P3_U2791 = ~(P3_U6686 & P3_U6685 & P3_U6687); 
assign P3_U2792 = ~(P3_U6683 & P3_U6682 & P3_U6684); 
assign P3_U2793 = ~(P3_U6680 & P3_U6679 & P3_U6681); 
assign P3_U2794 = ~(P3_U6677 & P3_U6676 & P3_U6678); 
assign P3_U2795 = ~(P3_U6674 & P3_U6673 & P3_U6675); 
assign P3_U2796 = ~(P3_U6671 & P3_U6670 & P3_U6672); 
assign P3_U2797 = ~(P3_U6668 & P3_U6667 & P3_U6669); 
assign P3_U2798 = ~(P3_U6665 & P3_U6664 & P3_U6666); 
assign P3_U2866 = ~(P3_U5591 & P3_U5590); 
assign P3_U3676 = P3_U3677 & P3_U5539 & P3_U3675; 
assign P3_U3679 = P3_U3678 & P3_U5551; 
assign P3_U3706 = P3_U3707 & P3_U5681; 
assign P3_U3769 = P3_U5876 & P3_U5875; 
assign P3_U3771 = P3_U5878 & P3_U5877 & P3_U5879 & P3_U3770; 
assign P3_U3773 = P3_U5890 & P3_U5889 & P3_U5888 & P3_U5887; 
assign P3_U3777 = P3_U5905 & P3_U5904; 
assign P3_U3779 = P3_U5907 & P3_U5906 & P3_U5908 & P3_U5910 & P3_U5909; 
assign P3_U3954 = P3_U6412 & P3_U6411 & P3_U6410 & P3_U6409; 
assign P3_U3955 = P3_U6420 & P3_U6419 & P3_U6418 & P3_U6417; 
assign P3_U3987 = P3_U6809 & P3_U6810; 
assign P3_U3988 = P3_U6812 & P3_U6813; 
assign P3_U3989 = P3_U6815 & P3_U6816; 
assign P3_U3990 = P3_U6818 & P3_U6819; 
assign P3_U3991 = P3_U6821 & P3_U6822; 
assign P3_U3992 = P3_U6824 & P3_U6825; 
assign P3_U3993 = P3_U6827 & P3_U6828; 
assign P3_U3994 = P3_U6830 & P3_U6831; 
assign P3_U3995 = P3_U6833 & P3_U6834; 
assign P3_U3996 = P3_U6836 & P3_U6837; 
assign P3_U3997 = P3_U6839 & P3_U6840; 
assign P3_U3998 = P3_U6842 & P3_U6843; 
assign P3_U3999 = P3_U6845 & P3_U6846; 
assign P3_U4000 = P3_U6848 & P3_U6849; 
assign P3_U4001 = P3_U6851 & P3_U6852; 
assign P3_U4281 = ~(P3_U3361 & P3_U2604); 
assign P3_U4283 = ~(P3_U3658 & P3_U5497); 
assign P3_U4310 = ~P3_U3252; 
assign P3_U4316 = ~(P3_U4347 & P3_U3260); 
assign P3_U4678 = ~(P3_U2378 & P3_U2420); 
assign P3_U4683 = ~(P3_U2419 & P3_U2378); 
assign P3_U4688 = ~(P3_U2418 & P3_U2378); 
assign P3_U4693 = ~(P3_U2417 & P3_U2378); 
assign P3_U4698 = ~(P3_U2416 & P3_U2378); 
assign P3_U4703 = ~(P3_U2415 & P3_U2378); 
assign P3_U4708 = ~(P3_U2414 & P3_U2378); 
assign P3_U4713 = ~(P3_U2413 & P3_U2378); 
assign P3_U4730 = ~(P3_U2377 & P3_U2420); 
assign P3_U4735 = ~(P3_U2377 & P3_U2419); 
assign P3_U4740 = ~(P3_U2377 & P3_U2418); 
assign P3_U4745 = ~(P3_U2377 & P3_U2417); 
assign P3_U4750 = ~(P3_U2377 & P3_U2416); 
assign P3_U4755 = ~(P3_U2377 & P3_U2415); 
assign P3_U4760 = ~(P3_U2377 & P3_U2414); 
assign P3_U4765 = ~(P3_U2377 & P3_U2413); 
assign P3_U4782 = ~(P3_U2376 & P3_U2420); 
assign P3_U4787 = ~(P3_U2376 & P3_U2419); 
assign P3_U4792 = ~(P3_U2376 & P3_U2418); 
assign P3_U4797 = ~(P3_U2376 & P3_U2417); 
assign P3_U4802 = ~(P3_U2376 & P3_U2416); 
assign P3_U4807 = ~(P3_U2376 & P3_U2415); 
assign P3_U4812 = ~(P3_U2376 & P3_U2414); 
assign P3_U4817 = ~(P3_U2376 & P3_U2413); 
assign P3_U4833 = ~(P3_U2375 & P3_U2420); 
assign P3_U4838 = ~(P3_U2375 & P3_U2419); 
assign P3_U4843 = ~(P3_U2375 & P3_U2418); 
assign P3_U4848 = ~(P3_U2375 & P3_U2417); 
assign P3_U4853 = ~(P3_U2375 & P3_U2416); 
assign P3_U4858 = ~(P3_U2375 & P3_U2415); 
assign P3_U4863 = ~(P3_U2375 & P3_U2414); 
assign P3_U4868 = ~(P3_U2375 & P3_U2413); 
assign P3_U4885 = ~(P3_U2374 & P3_U2420); 
assign P3_U4890 = ~(P3_U2374 & P3_U2419); 
assign P3_U4895 = ~(P3_U2374 & P3_U2418); 
assign P3_U4900 = ~(P3_U2374 & P3_U2417); 
assign P3_U4905 = ~(P3_U2374 & P3_U2416); 
assign P3_U4910 = ~(P3_U2374 & P3_U2415); 
assign P3_U4915 = ~(P3_U2374 & P3_U2414); 
assign P3_U4920 = ~(P3_U2374 & P3_U2413); 
assign P3_U4937 = ~(P3_U2373 & P3_U2420); 
assign P3_U4942 = ~(P3_U2373 & P3_U2419); 
assign P3_U4947 = ~(P3_U2373 & P3_U2418); 
assign P3_U4952 = ~(P3_U2373 & P3_U2417); 
assign P3_U4957 = ~(P3_U2373 & P3_U2416); 
assign P3_U4962 = ~(P3_U2373 & P3_U2415); 
assign P3_U4967 = ~(P3_U2373 & P3_U2414); 
assign P3_U4972 = ~(P3_U2373 & P3_U2413); 
assign P3_U4989 = ~(P3_U2372 & P3_U2420); 
assign P3_U4994 = ~(P3_U2372 & P3_U2419); 
assign P3_U4999 = ~(P3_U2372 & P3_U2418); 
assign P3_U5004 = ~(P3_U2372 & P3_U2417); 
assign P3_U5009 = ~(P3_U2372 & P3_U2416); 
assign P3_U5014 = ~(P3_U2372 & P3_U2415); 
assign P3_U5019 = ~(P3_U2372 & P3_U2414); 
assign P3_U5024 = ~(P3_U2372 & P3_U2413); 
assign P3_U5040 = ~(P3_U2371 & P3_U2420); 
assign P3_U5045 = ~(P3_U2371 & P3_U2419); 
assign P3_U5050 = ~(P3_U2371 & P3_U2418); 
assign P3_U5055 = ~(P3_U2371 & P3_U2417); 
assign P3_U5060 = ~(P3_U2371 & P3_U2416); 
assign P3_U5065 = ~(P3_U2371 & P3_U2415); 
assign P3_U5070 = ~(P3_U2371 & P3_U2414); 
assign P3_U5075 = ~(P3_U2371 & P3_U2413); 
assign P3_U5090 = ~(P3_U5083 & P3_INSTQUEUE_REG_7__7__SCAN_IN); 
assign P3_U5095 = ~(P3_U5083 & P3_INSTQUEUE_REG_7__6__SCAN_IN); 
assign P3_U5100 = ~(P3_U5083 & P3_INSTQUEUE_REG_7__5__SCAN_IN); 
assign P3_U5105 = ~(P3_U5083 & P3_INSTQUEUE_REG_7__4__SCAN_IN); 
assign P3_U5110 = ~(P3_U5083 & P3_INSTQUEUE_REG_7__3__SCAN_IN); 
assign P3_U5115 = ~(P3_U5083 & P3_INSTQUEUE_REG_7__2__SCAN_IN); 
assign P3_U5120 = ~(P3_U5083 & P3_INSTQUEUE_REG_7__1__SCAN_IN); 
assign P3_U5125 = ~(P3_U5083 & P3_INSTQUEUE_REG_7__0__SCAN_IN); 
assign P3_U5142 = ~(P3_U5135 & P3_INSTQUEUE_REG_6__7__SCAN_IN); 
assign P3_U5147 = ~(P3_U5135 & P3_INSTQUEUE_REG_6__6__SCAN_IN); 
assign P3_U5152 = ~(P3_U5135 & P3_INSTQUEUE_REG_6__5__SCAN_IN); 
assign P3_U5157 = ~(P3_U5135 & P3_INSTQUEUE_REG_6__4__SCAN_IN); 
assign P3_U5162 = ~(P3_U5135 & P3_INSTQUEUE_REG_6__3__SCAN_IN); 
assign P3_U5167 = ~(P3_U5135 & P3_INSTQUEUE_REG_6__2__SCAN_IN); 
assign P3_U5172 = ~(P3_U5135 & P3_INSTQUEUE_REG_6__1__SCAN_IN); 
assign P3_U5177 = ~(P3_U5135 & P3_INSTQUEUE_REG_6__0__SCAN_IN); 
assign P3_U5194 = ~(P3_U5187 & P3_INSTQUEUE_REG_5__7__SCAN_IN); 
assign P3_U5199 = ~(P3_U5187 & P3_INSTQUEUE_REG_5__6__SCAN_IN); 
assign P3_U5204 = ~(P3_U5187 & P3_INSTQUEUE_REG_5__5__SCAN_IN); 
assign P3_U5209 = ~(P3_U5187 & P3_INSTQUEUE_REG_5__4__SCAN_IN); 
assign P3_U5214 = ~(P3_U5187 & P3_INSTQUEUE_REG_5__3__SCAN_IN); 
assign P3_U5219 = ~(P3_U5187 & P3_INSTQUEUE_REG_5__2__SCAN_IN); 
assign P3_U5224 = ~(P3_U5187 & P3_INSTQUEUE_REG_5__1__SCAN_IN); 
assign P3_U5229 = ~(P3_U5187 & P3_INSTQUEUE_REG_5__0__SCAN_IN); 
assign P3_U5244 = ~(P3_U5238 & P3_INSTQUEUE_REG_4__7__SCAN_IN); 
assign P3_U5249 = ~(P3_U5238 & P3_INSTQUEUE_REG_4__6__SCAN_IN); 
assign P3_U5254 = ~(P3_U5238 & P3_INSTQUEUE_REG_4__5__SCAN_IN); 
assign P3_U5259 = ~(P3_U5238 & P3_INSTQUEUE_REG_4__4__SCAN_IN); 
assign P3_U5264 = ~(P3_U5238 & P3_INSTQUEUE_REG_4__3__SCAN_IN); 
assign P3_U5269 = ~(P3_U5238 & P3_INSTQUEUE_REG_4__2__SCAN_IN); 
assign P3_U5274 = ~(P3_U5238 & P3_INSTQUEUE_REG_4__1__SCAN_IN); 
assign P3_U5279 = ~(P3_U5238 & P3_INSTQUEUE_REG_4__0__SCAN_IN); 
assign P3_U5295 = ~(P3_U5289 & P3_INSTQUEUE_REG_3__7__SCAN_IN); 
assign P3_U5300 = ~(P3_U5289 & P3_INSTQUEUE_REG_3__6__SCAN_IN); 
assign P3_U5305 = ~(P3_U5289 & P3_INSTQUEUE_REG_3__5__SCAN_IN); 
assign P3_U5310 = ~(P3_U5289 & P3_INSTQUEUE_REG_3__4__SCAN_IN); 
assign P3_U5315 = ~(P3_U5289 & P3_INSTQUEUE_REG_3__3__SCAN_IN); 
assign P3_U5320 = ~(P3_U5289 & P3_INSTQUEUE_REG_3__2__SCAN_IN); 
assign P3_U5325 = ~(P3_U5289 & P3_INSTQUEUE_REG_3__1__SCAN_IN); 
assign P3_U5330 = ~(P3_U5289 & P3_INSTQUEUE_REG_3__0__SCAN_IN); 
assign P3_U5346 = ~(P3_U5340 & P3_INSTQUEUE_REG_2__7__SCAN_IN); 
assign P3_U5351 = ~(P3_U5340 & P3_INSTQUEUE_REG_2__6__SCAN_IN); 
assign P3_U5356 = ~(P3_U5340 & P3_INSTQUEUE_REG_2__5__SCAN_IN); 
assign P3_U5361 = ~(P3_U5340 & P3_INSTQUEUE_REG_2__4__SCAN_IN); 
assign P3_U5366 = ~(P3_U5340 & P3_INSTQUEUE_REG_2__3__SCAN_IN); 
assign P3_U5371 = ~(P3_U5340 & P3_INSTQUEUE_REG_2__2__SCAN_IN); 
assign P3_U5376 = ~(P3_U5340 & P3_INSTQUEUE_REG_2__1__SCAN_IN); 
assign P3_U5381 = ~(P3_U5340 & P3_INSTQUEUE_REG_2__0__SCAN_IN); 
assign P3_U5397 = ~(P3_U5391 & P3_INSTQUEUE_REG_1__7__SCAN_IN); 
assign P3_U5402 = ~(P3_U5391 & P3_INSTQUEUE_REG_1__6__SCAN_IN); 
assign P3_U5407 = ~(P3_U5391 & P3_INSTQUEUE_REG_1__5__SCAN_IN); 
assign P3_U5412 = ~(P3_U5391 & P3_INSTQUEUE_REG_1__4__SCAN_IN); 
assign P3_U5417 = ~(P3_U5391 & P3_INSTQUEUE_REG_1__3__SCAN_IN); 
assign P3_U5422 = ~(P3_U5391 & P3_INSTQUEUE_REG_1__2__SCAN_IN); 
assign P3_U5427 = ~(P3_U5391 & P3_INSTQUEUE_REG_1__1__SCAN_IN); 
assign P3_U5432 = ~(P3_U5391 & P3_INSTQUEUE_REG_1__0__SCAN_IN); 
assign P3_U5447 = ~(P3_U5441 & P3_INSTQUEUE_REG_0__7__SCAN_IN); 
assign P3_U5452 = ~(P3_U5441 & P3_INSTQUEUE_REG_0__6__SCAN_IN); 
assign P3_U5457 = ~(P3_U5441 & P3_INSTQUEUE_REG_0__5__SCAN_IN); 
assign P3_U5462 = ~(P3_U5441 & P3_INSTQUEUE_REG_0__4__SCAN_IN); 
assign P3_U5467 = ~(P3_U5441 & P3_INSTQUEUE_REG_0__3__SCAN_IN); 
assign P3_U5472 = ~(P3_U5441 & P3_INSTQUEUE_REG_0__2__SCAN_IN); 
assign P3_U5477 = ~(P3_U5441 & P3_INSTQUEUE_REG_0__1__SCAN_IN); 
assign P3_U5482 = ~(P3_U5441 & P3_INSTQUEUE_REG_0__0__SCAN_IN); 
assign P3_U5530 = ~(P3_U5529 & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P3_U5561 = ~P3_U3230; 
assign P3_U5562 = ~(P3_U2466 & P3_U3230); 
assign P3_U5630 = ~(P3_U2390 & P3_U5629); 
assign P3_U5676 = ~(P3_U5658 & P3_U3699 & P3_U5656 & P3_U3705 & P3_U3700); 
assign P3_U5699 = ~(P3_ADD_371_1212_U93 & P3_U2360); 
assign P3_U6405 = ~(P3_U2398 & P3_PHYADDRPOINTER_REG_0__SCAN_IN); 
assign P3_U6406 = ~(P3_U2397 & P3_PHYADDRPOINTER_REG_0__SCAN_IN); 
assign P3_U6407 = ~(P3_U2396 & P3_ADD_360_1242_U85); 
assign P3_U6408 = ~(P3_U2394 & P3_SUB_357_1258_U69); 
assign P3_U6413 = ~(P3_ADD_318_U4 & P3_U2398); 
assign P3_U6414 = ~(P3_U2397 & P3_PHYADDRPOINTER_REG_1__SCAN_IN); 
assign P3_U6415 = ~(P3_U2396 & P3_ADD_360_1242_U19); 
assign P3_U6416 = ~(P3_U2394 & P3_SUB_357_1258_U21); 
assign P3_U6421 = ~(P3_ADD_318_U71 & P3_U2398); 
assign P3_U6422 = ~(P3_ADD_315_U4 & P3_U2397); 
assign P3_U6423 = ~(P3_U2396 & P3_ADD_360_1242_U91); 
assign P3_U6424 = ~(P3_U2394 & P3_SUB_357_1258_U78); 
assign P3_U6427 = ~(P3_U2387 & P3_ADD_371_1212_U93); 
assign P3_U6429 = ~(P3_ADD_318_U68 & P3_U2398); 
assign P3_U6430 = ~(P3_ADD_315_U66 & P3_U2397); 
assign P3_U6437 = ~(P3_ADD_318_U67 & P3_U2398); 
assign P3_U6438 = ~(P3_ADD_315_U65 & P3_U2397); 
assign P3_U6445 = ~(P3_ADD_318_U66 & P3_U2398); 
assign P3_U6446 = ~(P3_ADD_315_U64 & P3_U2397); 
assign P3_U6453 = ~(P3_ADD_318_U65 & P3_U2398); 
assign P3_U6454 = ~(P3_ADD_315_U63 & P3_U2397); 
assign P3_U6461 = ~(P3_ADD_318_U64 & P3_U2398); 
assign P3_U6462 = ~(P3_ADD_315_U62 & P3_U2397); 
assign P3_U6469 = ~(P3_ADD_318_U63 & P3_U2398); 
assign P3_U6470 = ~(P3_ADD_315_U61 & P3_U2397); 
assign P3_U6477 = ~(P3_ADD_318_U62 & P3_U2398); 
assign P3_U6478 = ~(P3_ADD_315_U60 & P3_U2397); 
assign P3_U6485 = ~(P3_ADD_318_U91 & P3_U2398); 
assign P3_U6486 = ~(P3_ADD_315_U88 & P3_U2397); 
assign P3_U6493 = ~(P3_ADD_318_U90 & P3_U2398); 
assign P3_U6494 = ~(P3_ADD_315_U87 & P3_U2397); 
assign P3_U6502 = ~(P3_ADD_315_U86 & P3_U2397); 
assign P3_U6808 = ~(P3_U2447 & P3_EAX_REG_16__SCAN_IN); 
assign P3_U6811 = ~(P3_U2447 & P3_EAX_REG_17__SCAN_IN); 
assign P3_U6814 = ~(P3_U2447 & P3_EAX_REG_18__SCAN_IN); 
assign P3_U6817 = ~(P3_U2447 & P3_EAX_REG_19__SCAN_IN); 
assign P3_U6820 = ~(P3_U2447 & P3_EAX_REG_20__SCAN_IN); 
assign P3_U6823 = ~(P3_U2447 & P3_EAX_REG_21__SCAN_IN); 
assign P3_U6826 = ~(P3_U2447 & P3_EAX_REG_22__SCAN_IN); 
assign P3_U6829 = ~(P3_U2447 & P3_EAX_REG_23__SCAN_IN); 
assign P3_U6832 = ~(P3_U2447 & P3_EAX_REG_24__SCAN_IN); 
assign P3_U6835 = ~(P3_U2447 & P3_EAX_REG_25__SCAN_IN); 
assign P3_U6838 = ~(P3_U2447 & P3_EAX_REG_26__SCAN_IN); 
assign P3_U6841 = ~(P3_U2447 & P3_EAX_REG_27__SCAN_IN); 
assign P3_U6844 = ~(P3_U2447 & P3_EAX_REG_28__SCAN_IN); 
assign P3_U6847 = ~(P3_U2447 & P3_EAX_REG_29__SCAN_IN); 
assign P3_U6850 = ~(P3_U2447 & P3_EAX_REG_30__SCAN_IN); 
assign P3_U6857 = ~(P3_U3252 & P3_EAX_REG_0__SCAN_IN); 
assign P3_U6861 = ~(P3_U3252 & P3_EAX_REG_1__SCAN_IN); 
assign P3_U6865 = ~(P3_U3252 & P3_EAX_REG_2__SCAN_IN); 
assign P3_U6869 = ~(P3_U3252 & P3_EAX_REG_3__SCAN_IN); 
assign P3_U6873 = ~(P3_U3252 & P3_EAX_REG_4__SCAN_IN); 
assign P3_U6877 = ~(P3_U3252 & P3_EAX_REG_5__SCAN_IN); 
assign P3_U6881 = ~(P3_U3252 & P3_EAX_REG_6__SCAN_IN); 
assign P3_U6885 = ~(P3_U3252 & P3_EAX_REG_7__SCAN_IN); 
assign P3_U6889 = ~(P3_U3252 & P3_EAX_REG_8__SCAN_IN); 
assign P3_U6893 = ~(P3_U3252 & P3_EAX_REG_9__SCAN_IN); 
assign P3_U6897 = ~(P3_U3252 & P3_EAX_REG_10__SCAN_IN); 
assign P3_U6901 = ~(P3_U3252 & P3_EAX_REG_11__SCAN_IN); 
assign P3_U6905 = ~(P3_U3252 & P3_EAX_REG_12__SCAN_IN); 
assign P3_U6909 = ~(P3_U3252 & P3_EAX_REG_13__SCAN_IN); 
assign P3_U6913 = ~(P3_U3252 & P3_EAX_REG_14__SCAN_IN); 
assign P3_U6917 = ~(P3_U3252 & P3_EAX_REG_15__SCAN_IN); 
assign P3_U6922 = ~(P3_U3252 & P3_EAX_REG_16__SCAN_IN); 
assign P3_U6927 = ~(P3_U3252 & P3_EAX_REG_17__SCAN_IN); 
assign P3_U6932 = ~(P3_U3252 & P3_EAX_REG_18__SCAN_IN); 
assign P3_U6937 = ~(P3_U3252 & P3_EAX_REG_19__SCAN_IN); 
assign P3_U6942 = ~(P3_U3252 & P3_EAX_REG_20__SCAN_IN); 
assign P3_U6947 = ~(P3_U3252 & P3_EAX_REG_21__SCAN_IN); 
assign P3_U6952 = ~(P3_U3252 & P3_EAX_REG_22__SCAN_IN); 
assign P3_U6957 = ~(P3_U3252 & P3_EAX_REG_23__SCAN_IN); 
assign P3_U6962 = ~(P3_U3252 & P3_EAX_REG_24__SCAN_IN); 
assign P3_U6967 = ~(P3_U3252 & P3_EAX_REG_25__SCAN_IN); 
assign P3_U6972 = ~(P3_U3252 & P3_EAX_REG_26__SCAN_IN); 
assign P3_U6977 = ~(P3_U3252 & P3_EAX_REG_27__SCAN_IN); 
assign P3_U6982 = ~(P3_U3252 & P3_EAX_REG_28__SCAN_IN); 
assign P3_U6987 = ~(P3_U3252 & P3_EAX_REG_29__SCAN_IN); 
assign P3_U6992 = ~(P3_U3252 & P3_EAX_REG_30__SCAN_IN); 
assign P3_U6995 = ~(P3_U3252 & P3_EAX_REG_31__SCAN_IN); 
assign P3_U7079 = ~(P3_ADD_402_1132_U21 & P3_U2408); 
assign P3_U7094 = ~P3_U3260; 
assign P3_U7374 = ~P3_U4287; 
assign P3_U7380 = ~(P3_U2390 & P3_U2604); 
assign P3_U7384 = ~P3_U4288; 
assign P3_U8023 = ~(P3_U7379 & P3_U4287); 
assign P3_U8029 = ~(P3_U7385 & P3_U4288); 
assign P3_U8031 = ~(P3_U7386 & P3_U4288); 
assign P3_U8045 = ~(P3_U5496 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_U8046 = ~(P3_U5496 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_U8048 = ~(P3_U5496 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_U8050 = ~(P3_U5496 & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P3_U8052 = ~(P3_U5496 & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P2_U2685 = P2_ADD_402_1132_U22 & P2_U2355; 
assign P2_U2702 = ~(P2_U7164 & P2_U7165 & P2_U7163); 
assign P2_U2712 = ~(P2_U7871 & P2_U4407 & P2_STATE2_REG_0__SCAN_IN); 
assign P2_U3644 = ~(P2_U8342 & P2_U8341); 
assign P2_U3679 = ~(P2_U8414 & P2_U8413); 
assign P2_U5637 = ~(P2_U3890 & P2_U5636); 
assign P2_U6134 = ~(P2_U2395 & P2_EAX_REG_15__SCAN_IN); 
assign P2_U6135 = ~(U308 & P2_U2394); 
assign P2_U6137 = ~(P2_U2395 & P2_EAX_REG_14__SCAN_IN); 
assign P2_U6138 = ~(U309 & P2_U2394); 
assign P2_U6140 = ~(P2_U2395 & P2_EAX_REG_13__SCAN_IN); 
assign P2_U6141 = ~(U310 & P2_U2394); 
assign P2_U6143 = ~(P2_U2395 & P2_EAX_REG_12__SCAN_IN); 
assign P2_U6144 = ~(U311 & P2_U2394); 
assign P2_U6146 = ~(P2_U2395 & P2_EAX_REG_11__SCAN_IN); 
assign P2_U6147 = ~(U312 & P2_U2394); 
assign P2_U6149 = ~(P2_U2395 & P2_EAX_REG_10__SCAN_IN); 
assign P2_U6150 = ~(U313 & P2_U2394); 
assign P2_U6152 = ~(P2_U2395 & P2_EAX_REG_9__SCAN_IN); 
assign P2_U6153 = ~(U283 & P2_U2394); 
assign P2_U6155 = ~(P2_U2395 & P2_EAX_REG_8__SCAN_IN); 
assign P2_U6156 = ~(U284 & P2_U2394); 
assign P2_U6158 = ~(P2_U2395 & P2_EAX_REG_7__SCAN_IN); 
assign P2_U6159 = ~(P2_U2394 & U285); 
assign P2_U6161 = ~(P2_U2395 & P2_EAX_REG_6__SCAN_IN); 
assign P2_U6162 = ~(P2_U2394 & U286); 
assign P2_U6164 = ~(P2_U2395 & P2_EAX_REG_5__SCAN_IN); 
assign P2_U6165 = ~(P2_U2394 & U287); 
assign P2_U6167 = ~(P2_U2395 & P2_EAX_REG_4__SCAN_IN); 
assign P2_U6168 = ~(P2_U2394 & U288); 
assign P2_U6170 = ~(P2_U2395 & P2_EAX_REG_3__SCAN_IN); 
assign P2_U6171 = ~(P2_U2394 & U289); 
assign P2_U6173 = ~(P2_U2395 & P2_EAX_REG_2__SCAN_IN); 
assign P2_U6174 = ~(P2_U2394 & U292); 
assign P2_U6176 = ~(P2_U2395 & P2_EAX_REG_1__SCAN_IN); 
assign P2_U6177 = ~(P2_U2394 & U303); 
assign P2_U6179 = ~(P2_U2395 & P2_EAX_REG_0__SCAN_IN); 
assign P2_U6180 = ~(P2_U2394 & U314); 
assign P2_U6182 = ~(P2_U2395 & P2_EAX_REG_30__SCAN_IN); 
assign P2_U6183 = ~(U309 & P2_U2394); 
assign P2_U6185 = ~(P2_U2395 & P2_EAX_REG_29__SCAN_IN); 
assign P2_U6186 = ~(U310 & P2_U2394); 
assign P2_U6188 = ~(P2_U2395 & P2_EAX_REG_28__SCAN_IN); 
assign P2_U6189 = ~(U311 & P2_U2394); 
assign P2_U6191 = ~(P2_U2395 & P2_EAX_REG_27__SCAN_IN); 
assign P2_U6192 = ~(U312 & P2_U2394); 
assign P2_U6194 = ~(P2_U2395 & P2_EAX_REG_26__SCAN_IN); 
assign P2_U6195 = ~(U313 & P2_U2394); 
assign P2_U6197 = ~(P2_U2395 & P2_EAX_REG_25__SCAN_IN); 
assign P2_U6198 = ~(U283 & P2_U2394); 
assign P2_U6200 = ~(P2_U2395 & P2_EAX_REG_24__SCAN_IN); 
assign P2_U6201 = ~(U284 & P2_U2394); 
assign P2_U6203 = ~(P2_U2395 & P2_EAX_REG_23__SCAN_IN); 
assign P2_U6204 = ~(P2_U2394 & U285); 
assign P2_U6206 = ~(P2_U2395 & P2_EAX_REG_22__SCAN_IN); 
assign P2_U6207 = ~(P2_U2394 & U286); 
assign P2_U6209 = ~(P2_U2395 & P2_EAX_REG_21__SCAN_IN); 
assign P2_U6210 = ~(P2_U2394 & U287); 
assign P2_U6212 = ~(P2_U2395 & P2_EAX_REG_20__SCAN_IN); 
assign P2_U6213 = ~(P2_U2394 & U288); 
assign P2_U6215 = ~(P2_U2395 & P2_EAX_REG_19__SCAN_IN); 
assign P2_U6216 = ~(P2_U2394 & U289); 
assign P2_U6218 = ~(P2_U2395 & P2_EAX_REG_18__SCAN_IN); 
assign P2_U6219 = ~(P2_U2394 & U292); 
assign P2_U6221 = ~(P2_U2395 & P2_EAX_REG_17__SCAN_IN); 
assign P2_U6222 = ~(P2_U2394 & U303); 
assign P2_U6224 = ~(P2_U2395 & P2_EAX_REG_16__SCAN_IN); 
assign P2_U6225 = ~(P2_U2394 & U314); 
assign P2_U8330 = ~(P2_U3242 & P2_R2267_U21); 
assign P1_U2609 = ~(P1_U6853 & P1_U6854 & P1_U6855); 
assign P1_U5533 = ~(P1_U2427 & P1_U5531); 
assign P1_U6792 = ~(P1_R2182_U30 & P1_U6746); 
assign P1_U6796 = ~(P1_R2182_U31 & P1_U6746); 
assign P3_ADD_526_U69 = ~(P3_ADD_526_U178 & P3_ADD_526_U177); 
assign P3_ADD_526_U70 = ~(P3_ADD_526_U180 & P3_ADD_526_U179); 
assign P3_ADD_526_U115 = ~P3_ADD_526_U40; 
assign P3_ADD_526_U134 = ~P3_ADD_526_U104; 
assign P3_ADD_526_U174 = ~(P3_ADD_526_U40 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_526_U175 = ~(P3_ADD_526_U104 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_552_U69 = ~(P3_ADD_552_U178 & P3_ADD_552_U177); 
assign P3_ADD_552_U70 = ~(P3_ADD_552_U180 & P3_ADD_552_U179); 
assign P3_ADD_552_U115 = ~P3_ADD_552_U40; 
assign P3_ADD_552_U134 = ~P3_ADD_552_U104; 
assign P3_ADD_552_U174 = ~(P3_ADD_552_U40 & P3_EBX_REG_23__SCAN_IN); 
assign P3_ADD_552_U175 = ~(P3_ADD_552_U104 & P3_EBX_REG_22__SCAN_IN); 
assign P3_ADD_546_U69 = ~(P3_ADD_546_U178 & P3_ADD_546_U177); 
assign P3_ADD_546_U70 = ~(P3_ADD_546_U180 & P3_ADD_546_U179); 
assign P3_ADD_546_U115 = ~P3_ADD_546_U40; 
assign P3_ADD_546_U134 = ~P3_ADD_546_U104; 
assign P3_ADD_546_U174 = ~(P3_ADD_546_U40 & P3_EAX_REG_23__SCAN_IN); 
assign P3_ADD_546_U175 = ~(P3_ADD_546_U104 & P3_EAX_REG_22__SCAN_IN); 
assign P3_ADD_391_1180_U16 = ~(P3_U2618 & P3_ADD_391_1180_U32); 
assign P3_ADD_391_1180_U40 = ~(P3_ADD_391_1180_U32 & P3_ADD_391_1180_U15); 
assign P3_ADD_476_U89 = ~(P3_ADD_476_U178 & P3_ADD_476_U177); 
assign P3_ADD_476_U104 = ~P3_ADD_476_U26; 
assign P3_ADD_476_U175 = ~(P3_ADD_476_U26 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_531_U94 = ~(P3_ADD_531_U187 & P3_ADD_531_U186); 
assign P3_ADD_531_U108 = ~P3_ADD_531_U27; 
assign P3_ADD_531_U184 = ~(P3_ADD_531_U27 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_SUB_320_U123 = ~(P3_SUB_320_U93 & P3_SUB_320_U81); 
assign P3_SUB_320_U159 = ~(P3_SUB_320_U93 & P3_SUB_320_U81); 
assign P3_ADD_318_U89 = ~(P3_ADD_318_U178 & P3_ADD_318_U177); 
assign P3_ADD_318_U104 = ~P3_ADD_318_U26; 
assign P3_ADD_318_U175 = ~(P3_ADD_318_U26 & P3_PHYADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_315_U85 = ~(P3_ADD_315_U170 & P3_ADD_315_U169); 
assign P3_ADD_315_U101 = ~P3_ADD_315_U26; 
assign P3_ADD_315_U167 = ~(P3_ADD_315_U26 & P3_PHYADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_360_1242_U17 = P3_ADD_360_1242_U153 & P3_ADD_360_1242_U152; 
assign P3_ADD_360_1242_U18 = P3_ADD_360_1242_U151 & P3_ADD_360_1242_U149; 
assign P3_ADD_360_1242_U33 = ~P3_ADD_360_U17; 
assign P3_ADD_360_1242_U113 = P3_ADD_360_1242_U217 & P3_ADD_360_1242_U216; 
assign P3_ADD_360_1242_U121 = ~(P3_ADD_360_1242_U114 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_360_1242_U136 = ~P3_ADD_360_1242_U114; 
assign P3_ADD_360_1242_U137 = ~(P3_ADD_360_U18 & P3_ADD_360_1242_U114); 
assign P3_ADD_360_1242_U139 = P3_ADD_360_U17 | P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_360_1242_U141 = ~(P3_ADD_360_U17 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_360_1242_U195 = ~(P3_ADD_360_1242_U37 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_360_1242_U197 = ~(P3_ADD_360_1242_U37 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_360_1242_U210 = ~(P3_ADD_360_U17 & P3_ADD_360_1242_U34); 
assign P3_ADD_360_1242_U212 = ~(P3_ADD_360_U17 & P3_ADD_360_1242_U34); 
assign P3_ADD_360_1242_U220 = ~(P3_ADD_360_1242_U219 & P3_ADD_360_1242_U218); 
assign P3_ADD_467_U89 = ~(P3_ADD_467_U178 & P3_ADD_467_U177); 
assign P3_ADD_467_U104 = ~P3_ADD_467_U26; 
assign P3_ADD_467_U175 = ~(P3_ADD_467_U26 & P3_REIP_REG_13__SCAN_IN); 
assign P3_ADD_430_U89 = ~(P3_ADD_430_U178 & P3_ADD_430_U177); 
assign P3_ADD_430_U104 = ~P3_ADD_430_U26; 
assign P3_ADD_430_U175 = ~(P3_ADD_430_U26 & P3_REIP_REG_13__SCAN_IN); 
assign P3_ADD_380_U94 = ~(P3_ADD_380_U187 & P3_ADD_380_U186); 
assign P3_ADD_380_U108 = ~P3_ADD_380_U27; 
assign P3_ADD_380_U184 = ~(P3_ADD_380_U27 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_344_U94 = ~(P3_ADD_344_U187 & P3_ADD_344_U186); 
assign P3_ADD_344_U108 = ~P3_ADD_344_U27; 
assign P3_ADD_344_U184 = ~(P3_ADD_344_U27 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_339_U89 = ~(P3_ADD_339_U178 & P3_ADD_339_U177); 
assign P3_ADD_339_U104 = ~P3_ADD_339_U26; 
assign P3_ADD_339_U175 = ~(P3_ADD_339_U26 & P3_PHYADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_360_U30 = ~(P3_ADD_360_U28 & P3_ADD_360_U14); 
assign P3_ADD_541_U89 = ~(P3_ADD_541_U178 & P3_ADD_541_U177); 
assign P3_ADD_541_U104 = ~P3_ADD_541_U26; 
assign P3_ADD_541_U175 = ~(P3_ADD_541_U26 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_SUB_357_1258_U13 = P3_SUB_357_1258_U11 & P3_SUB_357_1258_U213; 
assign P3_SUB_357_1258_U75 = ~(P3_SUB_357_1258_U345 & P3_SUB_357_1258_U344); 
assign P3_SUB_357_1258_U76 = ~(P3_SUB_357_1258_U350 & P3_SUB_357_1258_U349); 
assign P3_SUB_357_1258_U104 = P3_SUB_357_1258_U14 & P3_SUB_357_1258_U216; 
assign P3_SUB_357_1258_U118 = P3_SUB_357_1258_U321 & P3_SUB_357_1258_U320; 
assign P3_SUB_357_1258_U121 = ~(P3_SUB_357_1258_U298 & P3_SUB_357_1258_U266); 
assign P3_SUB_357_1258_U324 = ~(P3_SUB_357_1258_U323 & P3_SUB_357_1258_U322); 
assign P3_SUB_357_1258_U340 = ~(P3_SUB_357_1258_U169 & P3_SUB_357_1258_U338); 
assign P3_ADD_515_U89 = ~(P3_ADD_515_U178 & P3_ADD_515_U177); 
assign P3_ADD_515_U104 = ~P3_ADD_515_U26; 
assign P3_ADD_515_U175 = ~(P3_ADD_515_U26 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_394_U89 = ~(P3_ADD_394_U182 & P3_ADD_394_U181); 
assign P3_ADD_394_U107 = ~P3_ADD_394_U26; 
assign P3_ADD_394_U179 = ~(P3_ADD_394_U26 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_SUB_414_U70 = P3_SUB_414_U147 & P3_SUB_414_U146; 
assign P3_SUB_414_U99 = ~P3_SUB_414_U34; 
assign P3_SUB_414_U114 = ~(P3_SUB_414_U113 & P3_EBX_REG_22__SCAN_IN); 
assign P3_SUB_414_U144 = ~(P3_SUB_414_U34 & P3_EBX_REG_23__SCAN_IN); 
assign P3_ADD_441_U89 = ~(P3_ADD_441_U178 & P3_ADD_441_U177); 
assign P3_ADD_441_U104 = ~P3_ADD_441_U26; 
assign P3_ADD_441_U175 = ~(P3_ADD_441_U26 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_349_U94 = ~(P3_ADD_349_U187 & P3_ADD_349_U186); 
assign P3_ADD_349_U108 = ~P3_ADD_349_U27; 
assign P3_ADD_349_U184 = ~(P3_ADD_349_U27 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_405_U89 = ~(P3_ADD_405_U182 & P3_ADD_405_U181); 
assign P3_ADD_405_U107 = ~P3_ADD_405_U26; 
assign P3_ADD_405_U179 = ~(P3_ADD_405_U26 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_553_U94 = ~(P3_ADD_553_U187 & P3_ADD_553_U186); 
assign P3_ADD_553_U108 = ~P3_ADD_553_U27; 
assign P3_ADD_553_U184 = ~(P3_ADD_553_U27 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_558_U94 = ~(P3_ADD_558_U187 & P3_ADD_558_U186); 
assign P3_ADD_558_U108 = ~P3_ADD_558_U27; 
assign P3_ADD_558_U184 = ~(P3_ADD_558_U27 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_385_U94 = ~(P3_ADD_385_U187 & P3_ADD_385_U186); 
assign P3_ADD_385_U108 = ~P3_ADD_385_U27; 
assign P3_ADD_385_U184 = ~(P3_ADD_385_U27 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_547_U94 = ~(P3_ADD_547_U187 & P3_ADD_547_U186); 
assign P3_ADD_547_U108 = ~P3_ADD_547_U27; 
assign P3_ADD_547_U184 = ~(P3_ADD_547_U27 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_371_1212_U18 = P3_ADD_371_1212_U162 & P3_ADD_371_1212_U159; 
assign P3_ADD_371_1212_U36 = ~P3_ADD_371_U18; 
assign P3_ADD_371_1212_U96 = P3_ADD_371_1212_U228 & P3_ADD_371_1212_U227 & P3_ADD_371_1212_U24; 
assign P3_ADD_371_1212_U97 = P3_ADD_371_1212_U154 & P3_ADD_371_1212_U4; 
assign P3_ADD_371_1212_U131 = ~P3_ADD_371_1212_U43; 
assign P3_ADD_371_1212_U136 = ~(P3_ADD_371_1212_U135 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_ADD_371_1212_U138 = ~(P3_ADD_371_1212_U4 & P3_ADD_371_1212_U43); 
assign P3_ADD_371_1212_U140 = P3_ADD_371_U18 | P3_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P3_ADD_371_1212_U142 = ~(P3_ADD_371_U18 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_371_1212_U151 = ~(P3_ADD_371_1212_U150 & P3_ADD_371_1212_U43); 
assign P3_ADD_371_1212_U206 = ~(P3_ADD_371_1212_U40 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_371_1212_U208 = ~(P3_ADD_371_1212_U40 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_ADD_371_1212_U221 = ~(P3_ADD_371_U18 & P3_ADD_371_1212_U37); 
assign P3_ADD_371_1212_U223 = ~(P3_ADD_371_U18 & P3_ADD_371_1212_U37); 
assign P3_ADD_371_1212_U232 = ~(P3_ADD_371_1212_U197 & P3_ADD_371_1212_U43); 
assign P3_ADD_371_U34 = ~(P3_ADD_371_U31 & P3_ADD_371_U14); 
assign P3_ADD_494_U89 = ~(P3_ADD_494_U178 & P3_ADD_494_U177); 
assign P3_ADD_494_U104 = ~P3_ADD_494_U26; 
assign P3_ADD_494_U175 = ~(P3_ADD_494_U26 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_536_U89 = ~(P3_ADD_536_U178 & P3_ADD_536_U177); 
assign P3_ADD_536_U104 = ~P3_ADD_536_U26; 
assign P3_ADD_536_U175 = ~(P3_ADD_536_U26 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_402_1132_U16 = ~(P3_U2618 & P3_ADD_402_1132_U32); 
assign P3_ADD_402_1132_U40 = ~(P3_ADD_402_1132_U32 & P3_ADD_402_1132_U15); 
assign P2_R2099_U111 = ~P2_R2099_U104; 
assign P2_R2099_U113 = ~(P2_R2099_U112 & P2_R2099_U104); 
assign P2_R2099_U148 = ~(P2_R2099_U201 & P2_R2099_U9); 
assign P2_R2099_U177 = ~(P2_R2099_U103 & P2_R2099_U104); 
assign P2_ADD_402_1132_U16 = ~(P2_U2596 & P2_ADD_402_1132_U32); 
assign P2_ADD_402_1132_U48 = ~(P2_ADD_402_1132_U32 & P2_ADD_402_1132_U15); 
assign P2_R2182_U245 = ~(P2_U2662 & P2_R2182_U58); 
assign P2_R2182_U247 = ~(P2_U2662 & P2_R2182_U58); 
assign P2_R2167_U8 = ~P2_U2713; 
assign P2_R2167_U24 = ~(P2_U2713 & P2_R2167_U7); 
assign P2_R2027_U94 = ~(P2_R2027_U187 & P2_R2027_U186); 
assign P2_R2027_U108 = ~P2_R2027_U27; 
assign P2_R2027_U184 = ~(P2_R2027_U27 & P2_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P2_R2337_U87 = ~(P2_R2337_U176 & P2_R2337_U175); 
assign P2_R2337_U105 = ~P2_R2337_U27; 
assign P2_R2337_U173 = ~(P2_R2337_U27 & P2_PHYADDRPOINTER_REG_14__SCAN_IN); 
assign P2_R2219_U27 = ~(P2_R2219_U101 & P2_R2219_U100); 
assign P2_R2219_U28 = ~(P2_R2219_U106 & P2_R2219_U105); 
assign P2_R2219_U40 = ~(P2_R2219_U60 & P2_R2219_U59); 
assign P2_R2219_U95 = ~(P2_R2219_U57 & P2_R2219_U94); 
assign P2_R2096_U75 = ~(P2_R2096_U209 & P2_R2096_U208); 
assign P2_R2096_U127 = ~P2_R2096_U107; 
assign P2_R2096_U129 = ~(P2_R2096_U128 & P2_R2096_U107); 
assign P2_R2096_U201 = ~(P2_R2096_U106 & P2_R2096_U107); 
assign P2_R1957_U123 = ~(P2_R1957_U93 & P2_R1957_U81); 
assign P2_R1957_U159 = ~(P2_R1957_U93 & P2_R1957_U81); 
assign P2_ADD_394_U88 = ~(P2_ADD_394_U180 & P2_ADD_394_U179); 
assign P2_ADD_394_U107 = ~P2_ADD_394_U26; 
assign P2_ADD_394_U139 = ~(P2_ADD_394_U26 & P2_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P2_R2267_U76 = ~P2_U3645; 
assign P2_R2267_U155 = ~(P2_U3645 & P2_R2267_U77); 
assign P1_R2027_U69 = ~(P1_R2027_U178 & P1_R2027_U177); 
assign P1_R2027_U70 = ~(P1_R2027_U180 & P1_R2027_U179); 
assign P1_R2027_U115 = ~P1_R2027_U40; 
assign P1_R2027_U134 = ~P1_R2027_U104; 
assign P1_R2027_U174 = ~(P1_R2027_U40 & P1_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P1_R2027_U175 = ~(P1_R2027_U104 & P1_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P1_R2182_U22 = ~(P1_R2182_U48 & P1_U2734); 
assign P1_R2182_U33 = ~(P1_R2182_U84 & P1_R2182_U83); 
assign P1_R2182_U47 = ~P1_R2182_U13; 
assign P1_R2182_U55 = ~P1_R2182_U38; 
assign P1_R2182_U64 = ~(P1_U2740 & P1_R2182_U13); 
assign P1_R2182_U65 = ~(P1_U2741 & P1_R2182_U38); 
assign P1_R2182_U70 = ~(P1_R2182_U54 & P1_R2182_U10); 
assign P1_R2182_U73 = ~(P1_R2182_U48 & P1_R2182_U20); 
assign P1_R2182_U76 = ~(P1_R2182_U58 & P1_R2182_U18); 
assign P1_R2144_U54 = P1_R2144_U103 & P1_R2144_U151 & P1_R2144_U153 & P1_R2144_U152; 
assign P1_R2144_U74 = ~P1_U2768; 
assign P1_R2144_U189 = ~(P1_U2768 & P1_R2144_U12); 
assign P1_R2144_U191 = ~(P1_U2768 & P1_R2144_U12); 
assign P1_R2358_U150 = ~P1_U2672; 
assign P1_R2358_U161 = ~P1_U2610; 
assign P1_R2358_U403 = ~(P1_R2358_U402 & P1_R2358_U401); 
assign P1_R2358_U429 = ~(P1_U2672 & P1_R2358_U23); 
assign P1_R2358_U434 = ~(P1_U2672 & P1_R2358_U23); 
assign P1_R2358_U476 = ~(P1_U2610 & P1_R2358_U23); 
assign P1_R2358_U478 = ~(P1_U2610 & P1_R2358_U23); 
assign P1_R2099_U41 = ~(P1_R2099_U223 & P1_R2099_U222); 
assign P1_R2099_U42 = ~(P1_R2099_U225 & P1_R2099_U224); 
assign P1_R2099_U156 = ~P1_R2099_U111; 
assign P1_R2099_U157 = ~P1_R2099_U8; 
assign P1_R2099_U219 = ~(P1_R2099_U28 & P1_R2099_U8); 
assign P1_R2099_U221 = ~(P1_R2099_U31 & P1_R2099_U111); 
assign P1_R2167_U44 = ~(P1_R2167_U42 & P1_R2167_U6); 
assign P1_R2167_U47 = ~(P1_U2716 & P1_R2167_U42); 
assign P1_R2337_U89 = ~(P1_R2337_U178 & P1_R2337_U177); 
assign P1_R2337_U104 = ~P1_R2337_U26; 
assign P1_R2337_U175 = ~(P1_R2337_U26 & P1_PHYADDRPOINTER_REG_13__SCAN_IN); 
assign P1_R2096_U89 = ~(P1_R2096_U178 & P1_R2096_U177); 
assign P1_R2096_U104 = ~P1_R2096_U26; 
assign P1_R2096_U175 = ~(P1_R2096_U26 & P1_REIP_REG_13__SCAN_IN); 
assign P1_ADD_371_U21 = ~(P1_ADD_371_U44 & P1_ADD_371_U43); 
assign P1_ADD_405_U88 = ~(P1_ADD_405_U180 & P1_ADD_405_U179); 
assign P1_ADD_405_U107 = ~P1_ADD_405_U26; 
assign P1_ADD_405_U139 = ~(P1_ADD_405_U26 & P1_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P1_ADD_515_U88 = ~(P1_ADD_515_U176 & P1_ADD_515_U175); 
assign P1_ADD_515_U104 = ~P1_ADD_515_U26; 
assign P1_ADD_515_U137 = ~(P1_ADD_515_U26 & P1_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_U2383 = P3_U2380 & P3_U4296; 
assign P3_U2384 = P3_U2380 & P3_U4297; 
assign P3_U2391 = P3_U4310 & P3_U3218; 
assign P3_U2400 = P3_U4310 & P3_U4573; 
assign P3_U2411 = P3_U4310 & P3_U4608; 
assign P3_U2454 = P3_U2380 & P3_U4323; 
assign P3_U2455 = P3_U2380 & P3_U4324; 
assign P3_U2737 = ~(P3_U4001 & P3_U6850); 
assign P3_U2738 = ~(P3_U4000 & P3_U6847); 
assign P3_U2739 = ~(P3_U3999 & P3_U6844); 
assign P3_U2740 = ~(P3_U3998 & P3_U6841); 
assign P3_U2741 = ~(P3_U3997 & P3_U6838); 
assign P3_U2742 = ~(P3_U3996 & P3_U6835); 
assign P3_U2743 = ~(P3_U3995 & P3_U6832); 
assign P3_U2744 = ~(P3_U3994 & P3_U6829); 
assign P3_U2745 = ~(P3_U3993 & P3_U6826); 
assign P3_U2746 = ~(P3_U3992 & P3_U6823); 
assign P3_U2747 = ~(P3_U3991 & P3_U6820); 
assign P3_U2748 = ~(P3_U3990 & P3_U6817); 
assign P3_U2749 = ~(P3_U3989 & P3_U6814); 
assign P3_U2750 = ~(P3_U3988 & P3_U6811); 
assign P3_U2751 = ~(P3_U3987 & P3_U6808); 
assign P3_U2829 = ~(P3_U6416 & P3_U6415 & P3_U6414 & P3_U6413 & P3_U3955); 
assign P3_U2830 = ~(P3_U6408 & P3_U6407 & P3_U6406 & P3_U6405 & P3_U3954); 
assign P3_U2868 = ~(P3_U3651 & P3_U5482); 
assign P3_U2869 = ~(P3_U3649 & P3_U5477); 
assign P3_U2870 = ~(P3_U3647 & P3_U5472); 
assign P3_U2871 = ~(P3_U3645 & P3_U5467); 
assign P3_U2872 = ~(P3_U3643 & P3_U5462); 
assign P3_U2873 = ~(P3_U3641 & P3_U5457); 
assign P3_U2874 = ~(P3_U3639 & P3_U5452); 
assign P3_U2875 = ~(P3_U3637 & P3_U5447); 
assign P3_U2876 = ~(P3_U3633 & P3_U5432); 
assign P3_U2877 = ~(P3_U3631 & P3_U5427); 
assign P3_U2878 = ~(P3_U3629 & P3_U5422); 
assign P3_U2879 = ~(P3_U3627 & P3_U5417); 
assign P3_U2880 = ~(P3_U3625 & P3_U5412); 
assign P3_U2881 = ~(P3_U3623 & P3_U5407); 
assign P3_U2882 = ~(P3_U3621 & P3_U5402); 
assign P3_U2883 = ~(P3_U3619 & P3_U5397); 
assign P3_U2884 = ~(P3_U3615 & P3_U5381); 
assign P3_U2885 = ~(P3_U3613 & P3_U5376); 
assign P3_U2886 = ~(P3_U3611 & P3_U5371); 
assign P3_U2887 = ~(P3_U3609 & P3_U5366); 
assign P3_U2888 = ~(P3_U3607 & P3_U5361); 
assign P3_U2889 = ~(P3_U3605 & P3_U5356); 
assign P3_U2890 = ~(P3_U3603 & P3_U5351); 
assign P3_U2891 = ~(P3_U3601 & P3_U5346); 
assign P3_U2892 = ~(P3_U3598 & P3_U5330); 
assign P3_U2893 = ~(P3_U3596 & P3_U5325); 
assign P3_U2894 = ~(P3_U3594 & P3_U5320); 
assign P3_U2895 = ~(P3_U3592 & P3_U5315); 
assign P3_U2896 = ~(P3_U3590 & P3_U5310); 
assign P3_U2897 = ~(P3_U3588 & P3_U5305); 
assign P3_U2898 = ~(P3_U3586 & P3_U5300); 
assign P3_U2899 = ~(P3_U3584 & P3_U5295); 
assign P3_U2900 = ~(P3_U3580 & P3_U5279); 
assign P3_U2901 = ~(P3_U3578 & P3_U5274); 
assign P3_U2902 = ~(P3_U3576 & P3_U5269); 
assign P3_U2903 = ~(P3_U3574 & P3_U5264); 
assign P3_U2904 = ~(P3_U3572 & P3_U5259); 
assign P3_U2905 = ~(P3_U3570 & P3_U5254); 
assign P3_U2906 = ~(P3_U3568 & P3_U5249); 
assign P3_U2907 = ~(P3_U3566 & P3_U5244); 
assign P3_U2932 = ~(P3_U5076 & P3_U3509 & P3_U5075); 
assign P3_U2933 = ~(P3_U5071 & P3_U3507 & P3_U5070); 
assign P3_U2934 = ~(P3_U5066 & P3_U3505 & P3_U5065); 
assign P3_U2935 = ~(P3_U5061 & P3_U3503 & P3_U5060); 
assign P3_U2936 = ~(P3_U5056 & P3_U3501 & P3_U5055); 
assign P3_U2937 = ~(P3_U5051 & P3_U3499 & P3_U5050); 
assign P3_U2938 = ~(P3_U5046 & P3_U3497 & P3_U5045); 
assign P3_U2939 = ~(P3_U5041 & P3_U3495 & P3_U5040); 
assign P3_U2940 = ~(P3_U5025 & P3_U3492 & P3_U5024); 
assign P3_U2941 = ~(P3_U5020 & P3_U3490 & P3_U5019); 
assign P3_U2942 = ~(P3_U5015 & P3_U3488 & P3_U5014); 
assign P3_U2943 = ~(P3_U5010 & P3_U3486 & P3_U5009); 
assign P3_U2944 = ~(P3_U5005 & P3_U3484 & P3_U5004); 
assign P3_U2945 = ~(P3_U5000 & P3_U3482 & P3_U4999); 
assign P3_U2946 = ~(P3_U4995 & P3_U3480 & P3_U4994); 
assign P3_U2947 = ~(P3_U4990 & P3_U3478 & P3_U4989); 
assign P3_U2948 = ~(P3_U4973 & P3_U3474 & P3_U4972); 
assign P3_U2949 = ~(P3_U4968 & P3_U3472 & P3_U4967); 
assign P3_U2950 = ~(P3_U4963 & P3_U3470 & P3_U4962); 
assign P3_U2951 = ~(P3_U4958 & P3_U3468 & P3_U4957); 
assign P3_U2952 = ~(P3_U4953 & P3_U3466 & P3_U4952); 
assign P3_U2953 = ~(P3_U4948 & P3_U3464 & P3_U4947); 
assign P3_U2954 = ~(P3_U4943 & P3_U3462 & P3_U4942); 
assign P3_U2955 = ~(P3_U4938 & P3_U3460 & P3_U4937); 
assign P3_U2956 = ~(P3_U4921 & P3_U3456 & P3_U4920); 
assign P3_U2957 = ~(P3_U4916 & P3_U3454 & P3_U4915); 
assign P3_U2958 = ~(P3_U4911 & P3_U3452 & P3_U4910); 
assign P3_U2959 = ~(P3_U4906 & P3_U3450 & P3_U4905); 
assign P3_U2960 = ~(P3_U4901 & P3_U3448 & P3_U4900); 
assign P3_U2961 = ~(P3_U4896 & P3_U3446 & P3_U4895); 
assign P3_U2962 = ~(P3_U4891 & P3_U3444 & P3_U4890); 
assign P3_U2963 = ~(P3_U4886 & P3_U3442 & P3_U4885); 
assign P3_U2964 = ~(P3_U4869 & P3_U3439 & P3_U4868); 
assign P3_U2965 = ~(P3_U4864 & P3_U3437 & P3_U4863); 
assign P3_U2966 = ~(P3_U4859 & P3_U3435 & P3_U4858); 
assign P3_U2967 = ~(P3_U4854 & P3_U3433 & P3_U4853); 
assign P3_U2968 = ~(P3_U4849 & P3_U3431 & P3_U4848); 
assign P3_U2969 = ~(P3_U4844 & P3_U3429 & P3_U4843); 
assign P3_U2970 = ~(P3_U4839 & P3_U3427 & P3_U4838); 
assign P3_U2971 = ~(P3_U4834 & P3_U3425 & P3_U4833); 
assign P3_U2972 = ~(P3_U4818 & P3_U3421 & P3_U4817); 
assign P3_U2973 = ~(P3_U4813 & P3_U3419 & P3_U4812); 
assign P3_U2974 = ~(P3_U4808 & P3_U3417 & P3_U4807); 
assign P3_U2975 = ~(P3_U4803 & P3_U3415 & P3_U4802); 
assign P3_U2976 = ~(P3_U4798 & P3_U3413 & P3_U4797); 
assign P3_U2977 = ~(P3_U4793 & P3_U3411 & P3_U4792); 
assign P3_U2978 = ~(P3_U4788 & P3_U3409 & P3_U4787); 
assign P3_U2979 = ~(P3_U4783 & P3_U3407 & P3_U4782); 
assign P3_U2980 = ~(P3_U4766 & P3_U3403 & P3_U4765); 
assign P3_U2981 = ~(P3_U4761 & P3_U3401 & P3_U4760); 
assign P3_U2982 = ~(P3_U4756 & P3_U3399 & P3_U4755); 
assign P3_U2983 = ~(P3_U4751 & P3_U3397 & P3_U4750); 
assign P3_U2984 = ~(P3_U4746 & P3_U3395 & P3_U4745); 
assign P3_U2985 = ~(P3_U4741 & P3_U3393 & P3_U4740); 
assign P3_U2986 = ~(P3_U4736 & P3_U3391 & P3_U4735); 
assign P3_U2987 = ~(P3_U4731 & P3_U3389 & P3_U4730); 
assign P3_U2988 = ~(P3_U4714 & P3_U3385 & P3_U4713); 
assign P3_U2989 = ~(P3_U4709 & P3_U3383 & P3_U4708); 
assign P3_U2990 = ~(P3_U4704 & P3_U3381 & P3_U4703); 
assign P3_U2991 = ~(P3_U4699 & P3_U3379 & P3_U4698); 
assign P3_U2992 = ~(P3_U4694 & P3_U3377 & P3_U4693); 
assign P3_U2993 = ~(P3_U4689 & P3_U3375 & P3_U4688); 
assign P3_U2994 = ~(P3_U4684 & P3_U3373 & P3_U4683); 
assign P3_U2995 = ~(P3_U4679 & P3_U3371 & P3_U4678); 
assign P3_U3248 = ~(P3_U4336 & P3_U5630); 
assign P3_U3304 = ~(P3_U8045 & P3_U8044); 
assign P3_U3681 = P3_U3682 & P3_U5562; 
assign P3_U3713 = P3_U3712 & P3_U3711 & P3_U5699; 
assign P3_U3956 = P3_U6426 & P3_U6425 & P3_U6428 & P3_U6427; 
assign P3_U4285 = ~(P3_U2390 & P3_U4281); 
assign P3_U4622 = ~P3_U4281; 
assign P3_U5089 = ~(P3_U2370 & P3_U2420); 
assign P3_U5094 = ~(P3_U2370 & P3_U2419); 
assign P3_U5099 = ~(P3_U2370 & P3_U2418); 
assign P3_U5104 = ~(P3_U2370 & P3_U2417); 
assign P3_U5109 = ~(P3_U2370 & P3_U2416); 
assign P3_U5114 = ~(P3_U2370 & P3_U2415); 
assign P3_U5119 = ~(P3_U2370 & P3_U2414); 
assign P3_U5124 = ~(P3_U2370 & P3_U2413); 
assign P3_U5141 = ~(P3_U2369 & P3_U2420); 
assign P3_U5146 = ~(P3_U2369 & P3_U2419); 
assign P3_U5151 = ~(P3_U2369 & P3_U2418); 
assign P3_U5156 = ~(P3_U2369 & P3_U2417); 
assign P3_U5161 = ~(P3_U2369 & P3_U2416); 
assign P3_U5166 = ~(P3_U2369 & P3_U2415); 
assign P3_U5171 = ~(P3_U2369 & P3_U2414); 
assign P3_U5176 = ~(P3_U2369 & P3_U2413); 
assign P3_U5193 = ~(P3_U2368 & P3_U2420); 
assign P3_U5198 = ~(P3_U2368 & P3_U2419); 
assign P3_U5203 = ~(P3_U2368 & P3_U2418); 
assign P3_U5208 = ~(P3_U2368 & P3_U2417); 
assign P3_U5213 = ~(P3_U2368 & P3_U2416); 
assign P3_U5218 = ~(P3_U2368 & P3_U2415); 
assign P3_U5223 = ~(P3_U2368 & P3_U2414); 
assign P3_U5228 = ~(P3_U2368 & P3_U2413); 
assign P3_U5499 = ~P3_U4283; 
assign P3_U5531 = ~(P3_U5525 & P3_U5530); 
assign P3_U5571 = ~(P3_U5560 & P3_U5561); 
assign P3_U5704 = ~(P3_ADD_360_1242_U17 & P3_U2395); 
assign P3_U5705 = ~(P3_SUB_357_1258_U76 & P3_U2393); 
assign P3_U5723 = ~(P3_ADD_371_1212_U18 & P3_U2360); 
assign P3_U5728 = ~(P3_ADD_360_1242_U18 & P3_U2395); 
assign P3_U5729 = ~(P3_SUB_357_1258_U75 & P3_U2393); 
assign P3_U5898 = ~(P3_ADD_558_U94 & P3_U3220); 
assign P3_U5899 = ~(P3_ADD_553_U94 & P3_U4298); 
assign P3_U5900 = ~(P3_ADD_547_U94 & P3_U4299); 
assign P3_U5903 = ~(P3_ADD_531_U94 & P3_U2354); 
assign P3_U5911 = ~(P3_ADD_385_U94 & P3_U2358); 
assign P3_U5912 = ~(P3_ADD_380_U94 & P3_U2359); 
assign P3_U5913 = ~(P3_ADD_349_U94 & P3_U4306); 
assign P3_U5914 = ~(P3_ADD_344_U94 & P3_U2362); 
assign P3_U5925 = ~(P3_ADD_541_U89 & P3_U4300); 
assign P3_U5926 = ~(P3_ADD_536_U89 & P3_U4301); 
assign P3_U5929 = ~(P3_ADD_515_U89 & P3_U4302); 
assign P3_U5930 = ~(P3_ADD_494_U89 & P3_U2356); 
assign P3_U5931 = ~(P3_ADD_476_U89 & P3_U4303); 
assign P3_U5932 = ~(P3_ADD_441_U89 & P3_U4304); 
assign P3_U5933 = ~(P3_ADD_405_U89 & P3_U4305); 
assign P3_U5934 = ~(P3_ADD_394_U89 & P3_U2357); 
assign P3_U6120 = ~(P3_ADD_526_U70 & P3_U2355); 
assign P3_U6144 = ~(P3_ADD_526_U69 & P3_U2355); 
assign P3_U6431 = ~(P3_U2396 & P3_ADD_360_1242_U17); 
assign P3_U6432 = ~(P3_U2394 & P3_SUB_357_1258_U76); 
assign P3_U6435 = ~(P3_U2387 & P3_ADD_371_1212_U18); 
assign P3_U6439 = ~(P3_U2396 & P3_ADD_360_1242_U18); 
assign P3_U6440 = ~(P3_U2394 & P3_SUB_357_1258_U75); 
assign P3_U6501 = ~(P3_ADD_318_U89 & P3_U2398); 
assign P3_U6506 = ~(P3_ADD_339_U89 & P3_U2388); 
assign P3_U6510 = ~(P3_ADD_315_U85 & P3_U2397); 
assign P3_U7059 = ~(P3_ADD_552_U70 & P3_U2399); 
assign P3_U7062 = ~(P3_ADD_552_U69 & P3_U2399); 
assign P3_U7105 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_0__SCAN_IN); 
assign P3_U7106 = ~(P3_U7094 & P3_REIP_REG_0__SCAN_IN); 
assign P3_U7115 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_1__SCAN_IN); 
assign P3_U7116 = ~(P3_U7094 & P3_REIP_REG_1__SCAN_IN); 
assign P3_U7125 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_2__SCAN_IN); 
assign P3_U7126 = ~(P3_U7094 & P3_REIP_REG_2__SCAN_IN); 
assign P3_U7135 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_3__SCAN_IN); 
assign P3_U7136 = ~(P3_U7094 & P3_REIP_REG_3__SCAN_IN); 
assign P3_U7145 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_4__SCAN_IN); 
assign P3_U7146 = ~(P3_U7094 & P3_REIP_REG_4__SCAN_IN); 
assign P3_U7155 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_5__SCAN_IN); 
assign P3_U7156 = ~(P3_U7094 & P3_REIP_REG_5__SCAN_IN); 
assign P3_U7163 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_6__SCAN_IN); 
assign P3_U7164 = ~(P3_U7094 & P3_REIP_REG_6__SCAN_IN); 
assign P3_U7171 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_7__SCAN_IN); 
assign P3_U7172 = ~(P3_U7094 & P3_REIP_REG_7__SCAN_IN); 
assign P3_U7179 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_8__SCAN_IN); 
assign P3_U7180 = ~(P3_U7094 & P3_REIP_REG_8__SCAN_IN); 
assign P3_U7187 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_9__SCAN_IN); 
assign P3_U7188 = ~(P3_U7094 & P3_REIP_REG_9__SCAN_IN); 
assign P3_U7195 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_10__SCAN_IN); 
assign P3_U7196 = ~(P3_U7094 & P3_REIP_REG_10__SCAN_IN); 
assign P3_U7203 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_11__SCAN_IN); 
assign P3_U7204 = ~(P3_U7094 & P3_REIP_REG_11__SCAN_IN); 
assign P3_U7211 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_12__SCAN_IN); 
assign P3_U7212 = ~(P3_U7094 & P3_REIP_REG_12__SCAN_IN); 
assign P3_U7219 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_13__SCAN_IN); 
assign P3_U7220 = ~(P3_U7094 & P3_REIP_REG_13__SCAN_IN); 
assign P3_U7227 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_14__SCAN_IN); 
assign P3_U7228 = ~(P3_U7094 & P3_REIP_REG_14__SCAN_IN); 
assign P3_U7235 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_15__SCAN_IN); 
assign P3_U7236 = ~(P3_U7094 & P3_REIP_REG_15__SCAN_IN); 
assign P3_U7243 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_16__SCAN_IN); 
assign P3_U7244 = ~(P3_U7094 & P3_REIP_REG_16__SCAN_IN); 
assign P3_U7251 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_17__SCAN_IN); 
assign P3_U7252 = ~(P3_U7094 & P3_REIP_REG_17__SCAN_IN); 
assign P3_U7259 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_18__SCAN_IN); 
assign P3_U7260 = ~(P3_U7094 & P3_REIP_REG_18__SCAN_IN); 
assign P3_U7267 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_19__SCAN_IN); 
assign P3_U7268 = ~(P3_U7094 & P3_REIP_REG_19__SCAN_IN); 
assign P3_U7275 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_20__SCAN_IN); 
assign P3_U7276 = ~(P3_U7094 & P3_REIP_REG_20__SCAN_IN); 
assign P3_U7283 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_21__SCAN_IN); 
assign P3_U7284 = ~(P3_U7094 & P3_REIP_REG_21__SCAN_IN); 
assign P3_U7291 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_22__SCAN_IN); 
assign P3_U7292 = ~(P3_U7094 & P3_REIP_REG_22__SCAN_IN); 
assign P3_U7299 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_23__SCAN_IN); 
assign P3_U7300 = ~(P3_U7094 & P3_REIP_REG_23__SCAN_IN); 
assign P3_U7307 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_24__SCAN_IN); 
assign P3_U7308 = ~(P3_U7094 & P3_REIP_REG_24__SCAN_IN); 
assign P3_U7315 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_25__SCAN_IN); 
assign P3_U7316 = ~(P3_U7094 & P3_REIP_REG_25__SCAN_IN); 
assign P3_U7323 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_26__SCAN_IN); 
assign P3_U7324 = ~(P3_U7094 & P3_REIP_REG_26__SCAN_IN); 
assign P3_U7331 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_27__SCAN_IN); 
assign P3_U7332 = ~(P3_U7094 & P3_REIP_REG_27__SCAN_IN); 
assign P3_U7339 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_28__SCAN_IN); 
assign P3_U7340 = ~(P3_U7094 & P3_REIP_REG_28__SCAN_IN); 
assign P3_U7347 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_29__SCAN_IN); 
assign P3_U7348 = ~(P3_U7094 & P3_REIP_REG_29__SCAN_IN); 
assign P3_U7355 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_30__SCAN_IN); 
assign P3_U7356 = ~(P3_U7094 & P3_REIP_REG_30__SCAN_IN); 
assign P3_U7364 = ~(P3_U2401 & P3_PHYADDRPOINTER_REG_31__SCAN_IN); 
assign P3_U7365 = ~(P3_U7094 & P3_REIP_REG_31__SCAN_IN); 
assign P3_U7381 = ~(P3_U7380 & P3_CODEFETCH_REG_SCAN_IN); 
assign P3_U7948 = ~(P3_U4281 & P3_U4617); 
assign P3_U7971 = ~(P3_U3283 & P3_U4283); 
assign P3_U8022 = ~(P3_U7374 & P3_REQUESTPENDING_REG_SCAN_IN); 
assign P3_U8028 = ~(P3_U7384 & P3_READREQUEST_REG_SCAN_IN); 
assign P3_U8030 = ~(P3_U7384 & P3_MEMORYFETCH_REG_SCAN_IN); 
assign P2_U2710 = P2_R2219_U27 & P2_U7723; 
assign P2_U2952 = ~(P2_U6225 & P2_U6224 & P2_U6226); 
assign P2_U2953 = ~(P2_U6222 & P2_U6221 & P2_U6223); 
assign P2_U2954 = ~(P2_U6219 & P2_U6218 & P2_U6220); 
assign P2_U2955 = ~(P2_U6216 & P2_U6215 & P2_U6217); 
assign P2_U2956 = ~(P2_U6213 & P2_U6212 & P2_U6214); 
assign P2_U2957 = ~(P2_U6210 & P2_U6209 & P2_U6211); 
assign P2_U2958 = ~(P2_U6207 & P2_U6206 & P2_U6208); 
assign P2_U2959 = ~(P2_U6204 & P2_U6203 & P2_U6205); 
assign P2_U2960 = ~(P2_U6201 & P2_U6200 & P2_U6202); 
assign P2_U2961 = ~(P2_U6198 & P2_U6197 & P2_U6199); 
assign P2_U2962 = ~(P2_U6195 & P2_U6194 & P2_U6196); 
assign P2_U2963 = ~(P2_U6192 & P2_U6191 & P2_U6193); 
assign P2_U2964 = ~(P2_U6189 & P2_U6188 & P2_U6190); 
assign P2_U2965 = ~(P2_U6186 & P2_U6185 & P2_U6187); 
assign P2_U2966 = ~(P2_U6183 & P2_U6182 & P2_U6184); 
assign P2_U2967 = ~(P2_U6180 & P2_U6179 & P2_U6181); 
assign P2_U2968 = ~(P2_U6177 & P2_U6176 & P2_U6178); 
assign P2_U2969 = ~(P2_U6174 & P2_U6173 & P2_U6175); 
assign P2_U2970 = ~(P2_U6171 & P2_U6170 & P2_U6172); 
assign P2_U2971 = ~(P2_U6168 & P2_U6167 & P2_U6169); 
assign P2_U2972 = ~(P2_U6165 & P2_U6164 & P2_U6166); 
assign P2_U2973 = ~(P2_U6162 & P2_U6161 & P2_U6163); 
assign P2_U2974 = ~(P2_U6159 & P2_U6158 & P2_U6160); 
assign P2_U2975 = ~(P2_U6156 & P2_U6155 & P2_U6157); 
assign P2_U2976 = ~(P2_U6153 & P2_U6152 & P2_U6154); 
assign P2_U2977 = ~(P2_U6150 & P2_U6149 & P2_U6151); 
assign P2_U2978 = ~(P2_U6147 & P2_U6146 & P2_U6148); 
assign P2_U2979 = ~(P2_U6144 & P2_U6143 & P2_U6145); 
assign P2_U2980 = ~(P2_U6141 & P2_U6140 & P2_U6142); 
assign P2_U2981 = ~(P2_U6138 & P2_U6137 & P2_U6139); 
assign P2_U2982 = ~(P2_U6135 & P2_U6134 & P2_U6136); 
assign P2_U5639 = ~(P2_U4466 & P2_U5637); 
assign P2_U5650 = ~(P2_R2096_U75 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U7724 = ~(P2_R2219_U28 & P2_U7723); 
assign P2_U8337 = ~(P2_R2219_U27 & P2_U2617); 
assign P2_U8339 = ~(P2_R2219_U28 & P2_U2617); 
assign P2_U8411 = ~(P2_R2337_U87 & P2_U3284); 
assign P1_U2442 = P1_R2182_U33 & P1_R2182_U34; 
assign P1_U2443 = P1_R2182_U33 & P1_U3318; 
assign P1_U2445 = ~(P1_R2182_U33 | P1_R2182_U34); 
assign P1_U3319 = ~P1_R2182_U33; 
assign P1_U5523 = ~(P1_R2182_U33 & P1_U7509); 
assign P1_U5552 = ~(P1_R2182_U33 & P1_U5538); 
assign P1_U6852 = ~(P1_R2337_U89 & P1_U2352); 
assign P1_U6859 = ~(P1_R2182_U33 & P1_U6746); 
assign P1_U6874 = ~(P1_ADD_371_U21 & P1_U4208); 
assign P1_U7043 = ~(P1_R2182_U33 & P1_U3294); 
assign P3_ADD_526_U43 = ~(P3_ADD_526_U92 & P3_ADD_526_U115); 
assign P3_ADD_526_U103 = ~(P3_ADD_526_U115 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_526_U173 = ~(P3_ADD_526_U115 & P3_ADD_526_U39); 
assign P3_ADD_526_U176 = ~(P3_ADD_526_U134 & P3_ADD_526_U37); 
assign P3_ADD_552_U43 = ~(P3_ADD_552_U92 & P3_ADD_552_U115); 
assign P3_ADD_552_U103 = ~(P3_ADD_552_U115 & P3_EBX_REG_23__SCAN_IN); 
assign P3_ADD_552_U173 = ~(P3_ADD_552_U115 & P3_ADD_552_U39); 
assign P3_ADD_552_U176 = ~(P3_ADD_552_U134 & P3_ADD_552_U37); 
assign P3_ADD_546_U43 = ~(P3_ADD_546_U92 & P3_ADD_546_U115); 
assign P3_ADD_546_U103 = ~(P3_ADD_546_U115 & P3_EAX_REG_23__SCAN_IN); 
assign P3_ADD_546_U173 = ~(P3_ADD_546_U115 & P3_ADD_546_U39); 
assign P3_ADD_546_U176 = ~(P3_ADD_546_U134 & P3_ADD_546_U37); 
assign P3_ADD_391_1180_U20 = ~(P3_ADD_391_1180_U40 & P3_ADD_391_1180_U39); 
assign P3_ADD_391_1180_U33 = ~P3_ADD_391_1180_U16; 
assign P3_ADD_391_1180_U37 = ~(P3_U2619 & P3_ADD_391_1180_U16); 
assign P3_ADD_476_U28 = ~(P3_ADD_476_U104 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_476_U176 = ~(P3_ADD_476_U104 & P3_ADD_476_U27); 
assign P3_ADD_531_U29 = ~(P3_ADD_531_U108 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_531_U185 = ~(P3_ADD_531_U108 & P3_ADD_531_U28); 
assign P3_SUB_320_U48 = ~P3_ADD_318_U89; 
assign P3_SUB_320_U82 = P3_SUB_320_U159 & P3_SUB_320_U158; 
assign P3_SUB_320_U124 = ~(P3_ADD_318_U89 & P3_SUB_320_U123); 
assign P3_ADD_318_U28 = ~(P3_ADD_318_U104 & P3_PHYADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_318_U176 = ~(P3_ADD_318_U104 & P3_ADD_318_U27); 
assign P3_ADD_315_U28 = ~(P3_ADD_315_U101 & P3_PHYADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_315_U168 = ~(P3_ADD_315_U101 & P3_ADD_315_U27); 
assign P3_ADD_360_1242_U107 = P3_ADD_360_1242_U196 & P3_ADD_360_1242_U195; 
assign P3_ADD_360_1242_U112 = ~(P3_ADD_360_1242_U137 & P3_ADD_360_1242_U121 & P3_ADD_360_1242_U188); 
assign P3_ADD_360_1242_U199 = ~(P3_ADD_360_1242_U198 & P3_ADD_360_1242_U197); 
assign P3_ADD_360_1242_U209 = ~(P3_ADD_360_1242_U33 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_360_1242_U211 = ~(P3_ADD_360_1242_U33 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_360_1242_U221 = ~(P3_ADD_360_1242_U113 & P3_ADD_360_1242_U114); 
assign P3_ADD_360_1242_U222 = ~(P3_ADD_360_1242_U136 & P3_ADD_360_1242_U220); 
assign P3_ADD_467_U28 = ~(P3_ADD_467_U104 & P3_REIP_REG_13__SCAN_IN); 
assign P3_ADD_467_U176 = ~(P3_ADD_467_U104 & P3_ADD_467_U27); 
assign P3_ADD_430_U28 = ~(P3_ADD_430_U104 & P3_REIP_REG_13__SCAN_IN); 
assign P3_ADD_430_U176 = ~(P3_ADD_430_U104 & P3_ADD_430_U27); 
assign P3_ADD_380_U29 = ~(P3_ADD_380_U108 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_380_U185 = ~(P3_ADD_380_U108 & P3_ADD_380_U28); 
assign P3_ADD_344_U29 = ~(P3_ADD_344_U108 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_344_U185 = ~(P3_ADD_344_U108 & P3_ADD_344_U28); 
assign P3_ADD_339_U28 = ~(P3_ADD_339_U104 & P3_PHYADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_339_U176 = ~(P3_ADD_339_U104 & P3_ADD_339_U27); 
assign P3_ADD_360_U16 = ~(P3_ADD_360_U30 & P3_ADD_360_U29); 
assign P3_ADD_541_U28 = ~(P3_ADD_541_U104 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_541_U176 = ~(P3_ADD_541_U104 & P3_ADD_541_U27); 
assign P3_SUB_357_1258_U74 = ~(P3_SUB_357_1258_U340 & P3_SUB_357_1258_U339); 
assign P3_SUB_357_1258_U103 = P3_SUB_357_1258_U215 & P3_SUB_357_1258_U13; 
assign P3_SUB_357_1258_U172 = ~(P3_SUB_357_1258_U171 & P3_SUB_357_1258_U121); 
assign P3_SUB_357_1258_U299 = ~P3_SUB_357_1258_U121; 
assign P3_SUB_357_1258_U332 = ~(P3_SUB_357_1258_U120 & P3_SUB_357_1258_U121); 
assign P3_ADD_515_U28 = ~(P3_ADD_515_U104 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_515_U176 = ~(P3_ADD_515_U104 & P3_ADD_515_U27); 
assign P3_ADD_394_U28 = ~(P3_ADD_394_U107 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_394_U180 = ~(P3_ADD_394_U107 & P3_ADD_394_U27); 
assign P3_SUB_414_U12 = P3_SUB_414_U114 & P3_SUB_414_U34; 
assign P3_SUB_414_U35 = ~(P3_SUB_414_U42 & P3_SUB_414_U67 & P3_SUB_414_U99); 
assign P3_SUB_414_U111 = ~(P3_SUB_414_U99 & P3_SUB_414_U67); 
assign P3_SUB_414_U145 = ~(P3_SUB_414_U99 & P3_SUB_414_U67); 
assign P3_ADD_441_U28 = ~(P3_ADD_441_U104 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_441_U176 = ~(P3_ADD_441_U104 & P3_ADD_441_U27); 
assign P3_ADD_349_U29 = ~(P3_ADD_349_U108 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_349_U185 = ~(P3_ADD_349_U108 & P3_ADD_349_U28); 
assign P3_ADD_405_U28 = ~(P3_ADD_405_U107 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_405_U180 = ~(P3_ADD_405_U107 & P3_ADD_405_U27); 
assign P3_ADD_553_U29 = ~(P3_ADD_553_U108 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_553_U185 = ~(P3_ADD_553_U108 & P3_ADD_553_U28); 
assign P3_ADD_558_U29 = ~(P3_ADD_558_U108 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_558_U185 = ~(P3_ADD_558_U108 & P3_ADD_558_U28); 
assign P3_ADD_385_U29 = ~(P3_ADD_385_U108 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_385_U185 = ~(P3_ADD_385_U108 & P3_ADD_385_U28); 
assign P3_ADD_547_U29 = ~(P3_ADD_547_U108 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_ADD_547_U185 = ~(P3_ADD_547_U108 & P3_ADD_547_U28); 
assign P3_ADD_371_1212_U95 = P3_ADD_371_1212_U137 & P3_ADD_371_1212_U136; 
assign P3_ADD_371_1212_U110 = P3_ADD_371_1212_U207 & P3_ADD_371_1212_U206; 
assign P3_ADD_371_1212_U152 = ~(P3_ADD_371_1212_U96 & P3_ADD_371_1212_U151); 
assign P3_ADD_371_1212_U153 = ~(P3_ADD_371_1212_U131 & P3_ADD_371_1212_U24); 
assign P3_ADD_371_1212_U210 = ~(P3_ADD_371_1212_U209 & P3_ADD_371_1212_U208); 
assign P3_ADD_371_1212_U220 = ~(P3_ADD_371_1212_U36 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_371_1212_U222 = ~(P3_ADD_371_1212_U36 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_ADD_371_1212_U233 = ~(P3_ADD_371_1212_U231 & P3_ADD_371_1212_U131); 
assign P3_ADD_371_U17 = ~(P3_ADD_371_U34 & P3_ADD_371_U33); 
assign P3_ADD_494_U28 = ~(P3_ADD_494_U104 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_494_U176 = ~(P3_ADD_494_U104 & P3_ADD_494_U27); 
assign P3_ADD_536_U28 = ~(P3_ADD_536_U104 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_536_U176 = ~(P3_ADD_536_U104 & P3_ADD_536_U27); 
assign P3_ADD_402_1132_U20 = ~(P3_ADD_402_1132_U40 & P3_ADD_402_1132_U39); 
assign P3_ADD_402_1132_U33 = ~P3_ADD_402_1132_U16; 
assign P3_ADD_402_1132_U37 = ~(P3_U2619 & P3_ADD_402_1132_U16); 
assign P2_R2099_U5 = ~(P2_R2099_U107 & P2_R2099_U148); 
assign P2_R2099_U100 = ~(P2_R2099_U114 & P2_R2099_U113); 
assign P2_R2099_U178 = ~(P2_R2099_U111 & P2_R2099_U176); 
assign P2_ADD_391_1196_U27 = ~P2_R2096_U75; 
assign P2_ADD_402_1132_U24 = ~(P2_ADD_402_1132_U48 & P2_ADD_402_1132_U47); 
assign P2_ADD_402_1132_U33 = ~P2_ADD_402_1132_U16; 
assign P2_ADD_402_1132_U37 = ~(P2_U2597 & P2_ADD_402_1132_U16); 
assign P2_R2182_U44 = ~P2_U2702; 
assign P2_R2182_U46 = ~(P2_U2681 & P2_U2702); 
assign P2_R2182_U60 = ~P2_U2685; 
assign P2_R2182_U114 = P2_R2182_U246 & P2_R2182_U245; 
assign P2_R2182_U171 = P2_U2685 | P2_U2661; 
assign P2_R2182_U173 = ~(P2_U2661 & P2_U2685); 
assign P2_R2182_U239 = ~(P2_U2685 & P2_R2182_U61); 
assign P2_R2182_U241 = ~(P2_U2685 & P2_R2182_U61); 
assign P2_R2182_U249 = ~(P2_R2182_U248 & P2_R2182_U247); 
assign P2_R2182_U305 = ~(P2_U2702 & P2_R2182_U45); 
assign P2_R2167_U9 = ~P2_U2712; 
assign P2_R2167_U22 = ~(P2_U2706 & P2_R2167_U8); 
assign P2_R2167_U25 = ~(P2_U2712 & P2_R2167_U10); 
assign P2_R2027_U29 = ~(P2_R2027_U108 & P2_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P2_R2027_U185 = ~(P2_R2027_U108 & P2_R2027_U28); 
assign P2_R2337_U29 = ~(P2_R2337_U105 & P2_PHYADDRPOINTER_REG_14__SCAN_IN); 
assign P2_R2337_U174 = ~(P2_R2337_U105 & P2_R2337_U28); 
assign P2_R2219_U26 = ~(P2_R2219_U96 & P2_R2219_U95); 
assign P2_R2219_U61 = ~P2_R2219_U40; 
assign P2_R2219_U63 = ~(P2_R2219_U62 & P2_R2219_U40); 
assign P2_R2219_U91 = ~(P2_R2219_U33 & P2_R2219_U40); 
assign P2_R2096_U105 = ~(P2_R2096_U130 & P2_R2096_U129); 
assign P2_R2096_U202 = ~(P2_R2096_U127 & P2_R2096_U200); 
assign P2_R1957_U47 = ~P2_U3679; 
assign P2_R1957_U82 = P2_R1957_U159 & P2_R1957_U158; 
assign P2_R1957_U124 = ~(P2_U3679 & P2_R1957_U123); 
assign P2_ADD_394_U28 = ~(P2_ADD_394_U107 & P2_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P2_ADD_394_U140 = ~(P2_ADD_394_U107 & P2_ADD_394_U27); 
assign P2_R2267_U23 = ~(P2_R2267_U76 & P2_R2267_U77); 
assign P2_R2267_U64 = ~P2_U3644; 
assign P2_R2267_U156 = ~(P2_R2267_U88 & P2_R2267_U76); 
assign P1_R2027_U43 = ~(P1_R2027_U92 & P1_R2027_U115); 
assign P1_R2027_U103 = ~(P1_R2027_U115 & P1_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P1_R2027_U173 = ~(P1_R2027_U115 & P1_R2027_U39); 
assign P1_R2027_U176 = ~(P1_R2027_U134 & P1_R2027_U37); 
assign P1_R2182_U5 = P1_R2182_U47 & P1_U2740; 
assign P1_R2182_U28 = ~(P1_R2182_U74 & P1_R2182_U73); 
assign P1_R2182_U29 = ~(P1_R2182_U76 & P1_R2182_U75); 
assign P1_R2182_U42 = P1_R2182_U70 & P1_R2182_U69; 
assign P1_R2182_U56 = ~P1_R2182_U22; 
assign P1_R2182_U63 = ~(P1_R2182_U47 & P1_R2182_U12); 
assign P1_R2182_U66 = ~(P1_R2182_U55 & P1_R2182_U11); 
assign P1_R2182_U71 = ~(P1_U2733 & P1_R2182_U22); 
assign P1_R2144_U188 = ~(P1_U2355 & P1_R2144_U74); 
assign P1_R2144_U190 = ~(P1_U2355 & P1_R2144_U74); 
assign P1_R2358_U162 = ~P1_U2609; 
assign P1_R2358_U428 = ~(P1_U2352 & P1_R2358_U150); 
assign P1_R2358_U433 = ~(P1_U2352 & P1_R2358_U150); 
assign P1_R2358_U475 = ~(P1_U2352 & P1_R2358_U161); 
assign P1_R2358_U477 = ~(P1_U2352 & P1_R2358_U161); 
assign P1_R2358_U481 = ~(P1_U2609 & P1_R2358_U23); 
assign P1_R2358_U483 = ~(P1_U2609 & P1_R2358_U23); 
assign P1_R2099_U9 = ~(P1_R2099_U90 & P1_R2099_U157); 
assign P1_R2099_U110 = ~(P1_R2099_U157 & P1_R2099_U28); 
assign P1_R2099_U218 = ~(P1_R2099_U205 & P1_R2099_U157); 
assign P1_R2099_U220 = ~(P1_R2099_U156 & P1_R2099_U202); 
assign P1_R2167_U45 = ~(P1_R2167_U44 & P1_R2167_U43); 
assign P1_R2167_U48 = ~(P1_R2167_U47 & P1_R2167_U46); 
assign P1_R2337_U28 = ~(P1_R2337_U104 & P1_PHYADDRPOINTER_REG_13__SCAN_IN); 
assign P1_R2337_U176 = ~(P1_R2337_U104 & P1_R2337_U27); 
assign P1_R2096_U28 = ~(P1_R2096_U104 & P1_REIP_REG_13__SCAN_IN); 
assign P1_R2096_U176 = ~(P1_R2096_U104 & P1_R2096_U27); 
assign P1_ADD_405_U28 = ~(P1_ADD_405_U107 & P1_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P1_ADD_405_U140 = ~(P1_ADD_405_U107 & P1_ADD_405_U27); 
assign P1_ADD_515_U28 = ~(P1_ADD_515_U104 & P1_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P1_ADD_515_U138 = ~(P1_ADD_515_U104 & P1_ADD_515_U27); 
assign P3_U2392 = P3_U2383 & P3_U4293; 
assign P3_U2402 = P3_U3248 & P3_U3090; 
assign P3_U2404 = P3_U2384 & P3_U3257; 
assign P3_U2405 = P3_U7095 & P3_U2384; 
assign P3_U2444 = P3_U2391 & P3_U3074; 
assign P3_U2446 = P3_U2391 & P3_U3113; 
assign P3_U2448 = P3_U2391 & P3_U4590; 
assign P3_U2634 = ~(P3_U7382 & P3_U7381); 
assign P3_U2682 = ~(P3_U7063 & P3_U7061 & P3_U7062); 
assign P3_U2683 = ~(P3_U7060 & P3_U7058 & P3_U7059); 
assign P3_U2828 = ~(P3_U6424 & P3_U6423 & P3_U6422 & P3_U6421 & P3_U3956); 
assign P3_U2908 = ~(P3_U5229 & P3_U3562 & P3_U5228); 
assign P3_U2909 = ~(P3_U5224 & P3_U3560 & P3_U5223); 
assign P3_U2910 = ~(P3_U5219 & P3_U3558 & P3_U5218); 
assign P3_U2911 = ~(P3_U5214 & P3_U3556 & P3_U5213); 
assign P3_U2912 = ~(P3_U5209 & P3_U3554 & P3_U5208); 
assign P3_U2913 = ~(P3_U5204 & P3_U3552 & P3_U5203); 
assign P3_U2914 = ~(P3_U5199 & P3_U3550 & P3_U5198); 
assign P3_U2915 = ~(P3_U5194 & P3_U3548 & P3_U5193); 
assign P3_U2916 = ~(P3_U5177 & P3_U3544 & P3_U5176); 
assign P3_U2917 = ~(P3_U5172 & P3_U3542 & P3_U5171); 
assign P3_U2918 = ~(P3_U5167 & P3_U3540 & P3_U5166); 
assign P3_U2919 = ~(P3_U5162 & P3_U3538 & P3_U5161); 
assign P3_U2920 = ~(P3_U5157 & P3_U3536 & P3_U5156); 
assign P3_U2921 = ~(P3_U5152 & P3_U3534 & P3_U5151); 
assign P3_U2922 = ~(P3_U5147 & P3_U3532 & P3_U5146); 
assign P3_U2923 = ~(P3_U5142 & P3_U3530 & P3_U5141); 
assign P3_U2924 = ~(P3_U5125 & P3_U3526 & P3_U5124); 
assign P3_U2925 = ~(P3_U5120 & P3_U3524 & P3_U5119); 
assign P3_U2926 = ~(P3_U5115 & P3_U3522 & P3_U5114); 
assign P3_U2927 = ~(P3_U5110 & P3_U3520 & P3_U5109); 
assign P3_U2928 = ~(P3_U5105 & P3_U3518 & P3_U5104); 
assign P3_U2929 = ~(P3_U5100 & P3_U3516 & P3_U5099); 
assign P3_U2930 = ~(P3_U5095 & P3_U3514 & P3_U5094); 
assign P3_U2931 = ~(P3_U5090 & P3_U3512 & P3_U5089); 
assign P3_U3247 = ~(P3_U3248 & P3_STATE2_REG_2__SCAN_IN); 
assign P3_U3296 = ~(P3_U8023 & P3_U8022); 
assign P3_U3298 = ~(P3_U8029 & P3_U8028); 
assign P3_U3299 = ~(P3_U8031 & P3_U8030); 
assign P3_U3714 = P3_U5705 & P3_U5704; 
assign P3_U3721 = P3_U3720 & P3_U3719 & P3_U5723; 
assign P3_U3722 = P3_U3723 & P3_U5729; 
assign P3_U3776 = P3_U5900 & P3_U5899; 
assign P3_U3778 = P3_U5902 & P3_U5901 & P3_U5903 & P3_U3777; 
assign P3_U3780 = P3_U5914 & P3_U5913 & P3_U5912 & P3_U5911; 
assign P3_U3784 = P3_U5929 & P3_U5928; 
assign P3_U3786 = P3_U5931 & P3_U5930 & P3_U5932 & P3_U5934 & P3_U5933; 
assign P3_U3957 = P3_U6434 & P3_U6433 & P3_U6436 & P3_U6435; 
assign P3_U4034 = P3_U7106 & P3_U7105; 
assign P3_U4038 = P3_U7116 & P3_U7115; 
assign P3_U4042 = P3_U7126 & P3_U7125; 
assign P3_U4046 = P3_U7136 & P3_U7135; 
assign P3_U4050 = P3_U7146 & P3_U7145; 
assign P3_U4055 = P3_U7156 & P3_U7155; 
assign P3_U4059 = P3_U7164 & P3_U7163; 
assign P3_U4062 = P3_U7172 & P3_U7171; 
assign P3_U4065 = P3_U7180 & P3_U7179; 
assign P3_U4068 = P3_U7188 & P3_U7187; 
assign P3_U4071 = P3_U7196 & P3_U7195; 
assign P3_U4074 = P3_U7204 & P3_U7203; 
assign P3_U4077 = P3_U7212 & P3_U7211; 
assign P3_U4080 = P3_U7220 & P3_U7219; 
assign P3_U4083 = P3_U7228 & P3_U7227; 
assign P3_U4086 = P3_U7236 & P3_U7235; 
assign P3_U4089 = P3_U7244 & P3_U7243; 
assign P3_U4092 = P3_U7252 & P3_U7251; 
assign P3_U4095 = P3_U7260 & P3_U7259; 
assign P3_U4098 = P3_U7268 & P3_U7267; 
assign P3_U4101 = P3_U7276 & P3_U7275; 
assign P3_U4104 = P3_U7284 & P3_U7283; 
assign P3_U4107 = P3_U7292 & P3_U7291; 
assign P3_U4110 = P3_U7300 & P3_U7299; 
assign P3_U4113 = P3_U7308 & P3_U7307; 
assign P3_U4116 = P3_U7316 & P3_U7315; 
assign P3_U4119 = P3_U7324 & P3_U7323; 
assign P3_U4122 = P3_U7332 & P3_U7331; 
assign P3_U4125 = P3_U7340 & P3_U7339; 
assign P3_U4128 = P3_U7348 & P3_U7347; 
assign P3_U4131 = P3_U7356 & P3_U7355; 
assign P3_U4132 = P3_U7364 & P3_U7365; 
assign P3_U4317 = ~(P3_U2383 & P3_U3105); 
assign P3_U5537 = ~(P3_U3669 & P3_U5531); 
assign P3_U5563 = ~(P3_U5531 & P3_U3094); 
assign P3_U5631 = ~P3_U3248; 
assign P3_U5700 = ~(P3_U5682 & P3_U3710 & P3_U5680 & P3_U3706 & P3_U3713); 
assign P3_U5753 = ~(P3_SUB_357_1258_U74 & P3_U2393); 
assign P3_U6448 = ~(P3_U2394 & P3_SUB_357_1258_U74); 
assign P3_U6855 = ~(P3_U2621 & P3_U2411); 
assign P3_U6856 = ~(P3_ADD_546_U5 & P3_U2400); 
assign P3_U6859 = ~(P3_U2622 & P3_U2411); 
assign P3_U6860 = ~(P3_ADD_546_U71 & P3_U2400); 
assign P3_U6863 = ~(P3_U2623 & P3_U2411); 
assign P3_U6864 = ~(P3_ADD_546_U60 & P3_U2400); 
assign P3_U6867 = ~(P3_U2624 & P3_U2411); 
assign P3_U6868 = ~(P3_ADD_546_U57 & P3_U2400); 
assign P3_U6871 = ~(P3_U2625 & P3_U2411); 
assign P3_U6872 = ~(P3_ADD_546_U56 & P3_U2400); 
assign P3_U6875 = ~(P3_U2626 & P3_U2411); 
assign P3_U6876 = ~(P3_ADD_546_U55 & P3_U2400); 
assign P3_U6879 = ~(P3_U2627 & P3_U2411); 
assign P3_U6880 = ~(P3_ADD_546_U54 & P3_U2400); 
assign P3_U6883 = ~(P3_U2628 & P3_U2411); 
assign P3_U6884 = ~(P3_ADD_546_U53 & P3_U2400); 
assign P3_U6887 = ~(P3_U2605 & P3_U2411); 
assign P3_U6888 = ~(P3_ADD_546_U52 & P3_U2400); 
assign P3_U6891 = ~(P3_U2606 & P3_U2411); 
assign P3_U6892 = ~(P3_ADD_546_U51 & P3_U2400); 
assign P3_U6895 = ~(P3_U2607 & P3_U2411); 
assign P3_U6896 = ~(P3_ADD_546_U81 & P3_U2400); 
assign P3_U6899 = ~(P3_U2608 & P3_U2411); 
assign P3_U6900 = ~(P3_ADD_546_U80 & P3_U2400); 
assign P3_U6903 = ~(P3_U2609 & P3_U2411); 
assign P3_U6904 = ~(P3_ADD_546_U79 & P3_U2400); 
assign P3_U6907 = ~(P3_U2610 & P3_U2411); 
assign P3_U6908 = ~(P3_ADD_546_U78 & P3_U2400); 
assign P3_U6911 = ~(P3_U2611 & P3_U2411); 
assign P3_U6912 = ~(P3_ADD_546_U77 & P3_U2400); 
assign P3_U6915 = ~(P3_U2612 & P3_U2411); 
assign P3_U6916 = ~(P3_ADD_546_U76 & P3_U2400); 
assign P3_U6920 = ~(P3_U3062 & P3_U2411); 
assign P3_U6921 = ~(P3_ADD_546_U75 & P3_U2400); 
assign P3_U6925 = ~(P3_U3063 & P3_U2411); 
assign P3_U6926 = ~(P3_ADD_546_U74 & P3_U2400); 
assign P3_U6930 = ~(P3_U3064 & P3_U2411); 
assign P3_U6931 = ~(P3_ADD_546_U73 & P3_U2400); 
assign P3_U6935 = ~(P3_U3065 & P3_U2411); 
assign P3_U6936 = ~(P3_ADD_546_U72 & P3_U2400); 
assign P3_U6940 = ~(P3_U3066 & P3_U2411); 
assign P3_U6941 = ~(P3_ADD_546_U70 & P3_U2400); 
assign P3_U6945 = ~(P3_U3067 & P3_U2411); 
assign P3_U6946 = ~(P3_ADD_546_U69 & P3_U2400); 
assign P3_U6950 = ~(P3_U3068 & P3_U2411); 
assign P3_U6955 = ~(P3_ADD_391_1180_U25 & P3_U2411); 
assign P3_U6960 = ~(P3_ADD_391_1180_U24 & P3_U2411); 
assign P3_U6965 = ~(P3_ADD_391_1180_U23 & P3_U2411); 
assign P3_U6970 = ~(P3_ADD_391_1180_U22 & P3_U2411); 
assign P3_U6975 = ~(P3_ADD_391_1180_U21 & P3_U2411); 
assign P3_U6980 = ~(P3_ADD_391_1180_U20 & P3_U2411); 
assign P3_U7082 = ~(P3_ADD_402_1132_U20 & P3_U2408); 
assign P3_U7100 = ~(P3_ADD_505_U5 & P3_U2455); 
assign P3_U7101 = ~(P3_ADD_486_U5 & P3_U2454); 
assign P3_U7110 = ~(P3_ADD_505_U17 & P3_U2455); 
assign P3_U7111 = ~(P3_ADD_486_U17 & P3_U2454); 
assign P3_U7120 = ~(P3_ADD_505_U16 & P3_U2455); 
assign P3_U7121 = ~(P3_ADD_486_U16 & P3_U2454); 
assign P3_U7130 = ~(P3_ADD_505_U15 & P3_U2455); 
assign P3_U7131 = ~(P3_ADD_486_U15 & P3_U2454); 
assign P3_U7140 = ~(P3_ADD_505_U14 & P3_U2455); 
assign P3_U7141 = ~(P3_ADD_486_U14 & P3_U2454); 
assign P3_U7150 = ~(P3_ADD_505_U6 & P3_U2455); 
assign P3_U7151 = ~(P3_ADD_486_U6 & P3_U2454); 
assign P3_U7368 = ~P3_U4285; 
assign P3_U7369 = ~(P3_U4285 & P3_FLUSH_REG_SCAN_IN); 
assign P3_U7949 = ~(P3_U4622 & P3_U4624); 
assign P3_U7972 = ~(P3_U5499 & P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P3_U7979 = ~(P3_U5499 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P3_U7982 = ~(P3_U5531 & P3_U3097 & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P3_U7989 = ~(P3_U5499 & P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P3_U7991 = ~(P3_U5499 & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P3_U7994 = ~(P3_U5571 & P3_U3093); 
assign P3_U7995 = ~(P3_U5499 & P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P3_U8019 = ~(P3_U4285 & P3_MORE_REG_SCAN_IN); 
assign P2_U2467 = P2_R2099_U5 & P2_R2099_U94; 
assign P2_U2470 = P2_R2099_U5 & P2_U3323; 
assign P2_U2479 = ~(P2_R2099_U94 | P2_R2099_U5); 
assign P2_U2684 = P2_ADD_402_1132_U24 & P2_U2355; 
assign P2_U2709 = P2_R2219_U26 & P2_U7723; 
assign P2_U2711 = ~(P2_U7724 & P2_STATE2_REG_0__SCAN_IN); 
assign P2_U3324 = ~P2_R2099_U5; 
assign P2_U3642 = ~(P2_U8338 & P2_U8337); 
assign P2_U3643 = ~(P2_U8340 & P2_U8339); 
assign P2_U3678 = ~(P2_U8412 & P2_U8411); 
assign P2_U5628 = ~(P2_R2099_U5 & P2_U5603); 
assign P2_U7160 = ~(P2_U4467 & P2_R2099_U5); 
assign P2_U8335 = ~(P2_R2219_U26 & P2_U2617); 
assign P1_U2444 = P1_R2182_U34 & P1_U3319; 
assign P1_U2616 = ~(P1_U6850 & P1_U6851 & P1_U6852); 
assign P1_U2671 = ~(P1_U6863 & P1_U6862 & P1_U4027 & P1_U6859); 
assign P1_U2767 = ~(P1_U7043 & P1_U7041 & P1_U7042); 
assign P1_U3317 = ~P1_R2182_U42; 
assign P1_U5512 = ~(P1_R2182_U42 & P1_U7509); 
assign P1_U5525 = ~(P1_U3750 & P1_U5523); 
assign P1_U5547 = ~(P1_R2182_U42 & P1_U5538); 
assign P1_U6759 = ~(P1_R2182_U5 & P1_U6746); 
assign P1_U6784 = ~(P1_R2182_U28 & P1_U6746); 
assign P1_U6788 = ~(P1_R2182_U29 & P1_U6746); 
assign P1_U6820 = ~(P1_R2182_U42 & P1_U6746); 
assign P1_U6940 = ~(P1_R2182_U42 & P1_U3294); 
assign P3_ADD_526_U67 = ~(P3_ADD_526_U174 & P3_ADD_526_U173); 
assign P3_ADD_526_U68 = ~(P3_ADD_526_U176 & P3_ADD_526_U175); 
assign P3_ADD_526_U116 = ~P3_ADD_526_U43; 
assign P3_ADD_526_U133 = ~P3_ADD_526_U103; 
assign P3_ADD_526_U170 = ~(P3_ADD_526_U43 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_526_U171 = ~(P3_ADD_526_U103 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_552_U67 = ~(P3_ADD_552_U174 & P3_ADD_552_U173); 
assign P3_ADD_552_U68 = ~(P3_ADD_552_U176 & P3_ADD_552_U175); 
assign P3_ADD_552_U116 = ~P3_ADD_552_U43; 
assign P3_ADD_552_U133 = ~P3_ADD_552_U103; 
assign P3_ADD_552_U170 = ~(P3_ADD_552_U43 & P3_EBX_REG_25__SCAN_IN); 
assign P3_ADD_552_U171 = ~(P3_ADD_552_U103 & P3_EBX_REG_24__SCAN_IN); 
assign P3_ADD_546_U67 = ~(P3_ADD_546_U174 & P3_ADD_546_U173); 
assign P3_ADD_546_U68 = ~(P3_ADD_546_U176 & P3_ADD_546_U175); 
assign P3_ADD_546_U116 = ~P3_ADD_546_U43; 
assign P3_ADD_546_U133 = ~P3_ADD_546_U103; 
assign P3_ADD_546_U170 = ~(P3_ADD_546_U43 & P3_EAX_REG_25__SCAN_IN); 
assign P3_ADD_546_U171 = ~(P3_ADD_546_U103 & P3_EAX_REG_24__SCAN_IN); 
assign P3_ADD_391_1180_U27 = ~(P3_U2619 & P3_ADD_391_1180_U33); 
assign P3_ADD_391_1180_U38 = ~(P3_ADD_391_1180_U33 & P3_ADD_391_1180_U17); 
assign P3_ADD_476_U88 = ~(P3_ADD_476_U176 & P3_ADD_476_U175); 
assign P3_ADD_476_U105 = ~P3_ADD_476_U28; 
assign P3_ADD_476_U173 = ~(P3_ADD_476_U28 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_531_U93 = ~(P3_ADD_531_U185 & P3_ADD_531_U184); 
assign P3_ADD_531_U109 = ~P3_ADD_531_U29; 
assign P3_ADD_531_U182 = ~(P3_ADD_531_U29 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_SUB_320_U29 = ~(P3_SUB_320_U48 & P3_SUB_320_U81 & P3_SUB_320_U93); 
assign P3_ADD_318_U88 = ~(P3_ADD_318_U176 & P3_ADD_318_U175); 
assign P3_ADD_318_U105 = ~P3_ADD_318_U28; 
assign P3_ADD_318_U173 = ~(P3_ADD_318_U28 & P3_PHYADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_315_U84 = ~(P3_ADD_315_U168 & P3_ADD_315_U167); 
assign P3_ADD_315_U102 = ~P3_ADD_315_U28; 
assign P3_ADD_315_U165 = ~(P3_ADD_315_U28 & P3_PHYADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_360_1242_U36 = ~P3_ADD_360_U16; 
assign P3_ADD_360_1242_U89 = ~(P3_ADD_360_1242_U222 & P3_ADD_360_1242_U221); 
assign P3_ADD_360_1242_U111 = P3_ADD_360_1242_U210 & P3_ADD_360_1242_U209; 
assign P3_ADD_360_1242_U138 = ~P3_ADD_360_1242_U112; 
assign P3_ADD_360_1242_U140 = ~(P3_ADD_360_1242_U139 & P3_ADD_360_1242_U112); 
assign P3_ADD_360_1242_U189 = ~(P3_ADD_360_U16 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_360_1242_U203 = ~(P3_ADD_360_U16 & P3_ADD_360_1242_U35); 
assign P3_ADD_360_1242_U205 = ~(P3_ADD_360_U16 & P3_ADD_360_1242_U35); 
assign P3_ADD_360_1242_U213 = ~(P3_ADD_360_1242_U212 & P3_ADD_360_1242_U211); 
assign P3_ADD_467_U88 = ~(P3_ADD_467_U176 & P3_ADD_467_U175); 
assign P3_ADD_467_U105 = ~P3_ADD_467_U28; 
assign P3_ADD_467_U173 = ~(P3_ADD_467_U28 & P3_REIP_REG_14__SCAN_IN); 
assign P3_ADD_430_U88 = ~(P3_ADD_430_U176 & P3_ADD_430_U175); 
assign P3_ADD_430_U105 = ~P3_ADD_430_U28; 
assign P3_ADD_430_U173 = ~(P3_ADD_430_U28 & P3_REIP_REG_14__SCAN_IN); 
assign P3_ADD_380_U93 = ~(P3_ADD_380_U185 & P3_ADD_380_U184); 
assign P3_ADD_380_U109 = ~P3_ADD_380_U29; 
assign P3_ADD_380_U182 = ~(P3_ADD_380_U29 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_344_U93 = ~(P3_ADD_344_U185 & P3_ADD_344_U184); 
assign P3_ADD_344_U109 = ~P3_ADD_344_U29; 
assign P3_ADD_344_U182 = ~(P3_ADD_344_U29 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_LT_563_U14 = ~P3_U3304; 
assign P3_LT_563_U26 = ~(P3_U3304 & P3_LT_563_U7); 
assign P3_ADD_339_U88 = ~(P3_ADD_339_U176 & P3_ADD_339_U175); 
assign P3_ADD_339_U105 = ~P3_ADD_339_U28; 
assign P3_ADD_339_U173 = ~(P3_ADD_339_U28 & P3_PHYADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_541_U88 = ~(P3_ADD_541_U176 & P3_ADD_541_U175); 
assign P3_ADD_541_U105 = ~P3_ADD_541_U28; 
assign P3_ADD_541_U173 = ~(P3_ADD_541_U28 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_SUB_357_1258_U119 = ~(P3_SUB_357_1258_U173 & P3_SUB_357_1258_U172); 
assign P3_SUB_357_1258_U333 = ~(P3_SUB_357_1258_U299 & P3_SUB_357_1258_U331); 
assign P3_ADD_515_U88 = ~(P3_ADD_515_U176 & P3_ADD_515_U175); 
assign P3_ADD_515_U105 = ~P3_ADD_515_U28; 
assign P3_ADD_515_U173 = ~(P3_ADD_515_U28 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_394_U88 = ~(P3_ADD_394_U180 & P3_ADD_394_U179); 
assign P3_ADD_394_U108 = ~P3_ADD_394_U28; 
assign P3_ADD_394_U177 = ~(P3_ADD_394_U28 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_SUB_414_U68 = P3_SUB_414_U145 & P3_SUB_414_U144; 
assign P3_SUB_414_U100 = ~P3_SUB_414_U35; 
assign P3_SUB_414_U112 = ~(P3_SUB_414_U111 & P3_EBX_REG_24__SCAN_IN); 
assign P3_SUB_414_U142 = ~(P3_SUB_414_U35 & P3_EBX_REG_25__SCAN_IN); 
assign P3_ADD_441_U88 = ~(P3_ADD_441_U176 & P3_ADD_441_U175); 
assign P3_ADD_441_U105 = ~P3_ADD_441_U28; 
assign P3_ADD_441_U173 = ~(P3_ADD_441_U28 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_349_U93 = ~(P3_ADD_349_U185 & P3_ADD_349_U184); 
assign P3_ADD_349_U109 = ~P3_ADD_349_U29; 
assign P3_ADD_349_U182 = ~(P3_ADD_349_U29 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_405_U88 = ~(P3_ADD_405_U180 & P3_ADD_405_U179); 
assign P3_ADD_405_U108 = ~P3_ADD_405_U28; 
assign P3_ADD_405_U177 = ~(P3_ADD_405_U28 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_553_U93 = ~(P3_ADD_553_U185 & P3_ADD_553_U184); 
assign P3_ADD_553_U109 = ~P3_ADD_553_U29; 
assign P3_ADD_553_U182 = ~(P3_ADD_553_U29 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_558_U93 = ~(P3_ADD_558_U185 & P3_ADD_558_U184); 
assign P3_ADD_558_U109 = ~P3_ADD_558_U29; 
assign P3_ADD_558_U182 = ~(P3_ADD_558_U29 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_385_U93 = ~(P3_ADD_385_U185 & P3_ADD_385_U184); 
assign P3_ADD_385_U109 = ~P3_ADD_385_U29; 
assign P3_ADD_385_U182 = ~(P3_ADD_385_U29 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_547_U93 = ~(P3_ADD_547_U185 & P3_ADD_547_U184); 
assign P3_ADD_547_U109 = ~P3_ADD_547_U29; 
assign P3_ADD_547_U182 = ~(P3_ADD_547_U29 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_371_1212_U39 = ~P3_ADD_371_U17; 
assign P3_ADD_371_1212_U91 = ~(P3_ADD_371_1212_U233 & P3_ADD_371_1212_U232); 
assign P3_ADD_371_1212_U114 = P3_ADD_371_1212_U221 & P3_ADD_371_1212_U220; 
assign P3_ADD_371_1212_U115 = ~(P3_ADD_371_1212_U95 & P3_ADD_371_1212_U138); 
assign P3_ADD_371_1212_U155 = ~(P3_ADD_371_1212_U97 & P3_ADD_371_1212_U153); 
assign P3_ADD_371_1212_U200 = ~(P3_ADD_371_U17 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_371_1212_U214 = ~(P3_ADD_371_U17 & P3_ADD_371_1212_U38); 
assign P3_ADD_371_1212_U216 = ~(P3_ADD_371_U17 & P3_ADD_371_1212_U38); 
assign P3_ADD_371_1212_U224 = ~(P3_ADD_371_1212_U223 & P3_ADD_371_1212_U222); 
assign P3_ADD_494_U88 = ~(P3_ADD_494_U176 & P3_ADD_494_U175); 
assign P3_ADD_494_U105 = ~P3_ADD_494_U28; 
assign P3_ADD_494_U173 = ~(P3_ADD_494_U28 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_536_U88 = ~(P3_ADD_536_U176 & P3_ADD_536_U175); 
assign P3_ADD_536_U105 = ~P3_ADD_536_U28; 
assign P3_ADD_536_U173 = ~(P3_ADD_536_U28 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_402_1132_U27 = ~(P3_U2619 & P3_ADD_402_1132_U33); 
assign P3_ADD_402_1132_U38 = ~(P3_ADD_402_1132_U33 & P3_ADD_402_1132_U17); 
assign P2_R2099_U96 = ~(P2_R2099_U178 & P2_R2099_U177); 
assign P2_R2099_U115 = ~P2_R2099_U100; 
assign P2_R2099_U117 = ~(P2_R2099_U116 & P2_R2099_U100); 
assign P2_R2099_U166 = ~(P2_R2099_U99 & P2_R2099_U100); 
assign P2_ADD_402_1132_U27 = ~(P2_U2597 & P2_ADD_402_1132_U33); 
assign P2_ADD_402_1132_U38 = ~(P2_ADD_402_1132_U33 & P2_ADD_402_1132_U17); 
assign P2_R2182_U121 = ~P2_R2182_U46; 
assign P2_R2182_U125 = ~(P2_R2182_U46 & P2_R2182_U47); 
assign P2_R2182_U187 = ~(P2_R2182_U47 & P2_R2182_U46); 
assign P2_R2182_U238 = ~(P2_U2661 & P2_R2182_U60); 
assign P2_R2182_U240 = ~(P2_U2661 & P2_R2182_U60); 
assign P2_R2182_U280 = ~(P2_U2680 & P2_R2182_U46); 
assign P2_R2182_U304 = ~(P2_U2681 & P2_R2182_U44); 
assign P2_R2167_U13 = ~P2_U2710; 
assign P2_R2167_U23 = ~(P2_R2167_U21 & P2_R2167_U20 & P2_R2167_U22); 
assign P2_R2167_U27 = ~(P2_U2705 & P2_R2167_U9); 
assign P2_R2167_U31 = ~(P2_U2710 & P2_R2167_U14); 
assign P2_R2027_U93 = ~(P2_R2027_U185 & P2_R2027_U184); 
assign P2_R2027_U109 = ~P2_R2027_U29; 
assign P2_R2027_U182 = ~(P2_R2027_U29 & P2_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P2_R2337_U86 = ~(P2_R2337_U174 & P2_R2337_U173); 
assign P2_R2337_U106 = ~P2_R2337_U29; 
assign P2_R2337_U171 = ~(P2_R2337_U29 & P2_PHYADDRPOINTER_REG_15__SCAN_IN); 
assign P2_R2219_U39 = ~(P2_R2219_U64 & P2_R2219_U63); 
assign P2_R2219_U90 = ~(P2_R2219_U61 & P2_R2219_U89); 
assign P2_R2096_U74 = ~(P2_R2096_U202 & P2_R2096_U201); 
assign P2_R2096_U131 = ~P2_R2096_U105; 
assign P2_R2096_U133 = ~(P2_R2096_U132 & P2_R2096_U105); 
assign P2_R2096_U194 = ~(P2_R2096_U104 & P2_R2096_U105); 
assign P2_GTE_370_U8 = ~(P2_R2219_U26 | P2_R2219_U27 | P2_R2219_U28 | P2_GTE_370_U7); 
assign P2_R1957_U28 = ~(P2_R1957_U93 & P2_R1957_U81 & P2_R1957_U47); 
assign P2_ADD_394_U69 = ~(P2_ADD_394_U140 & P2_ADD_394_U139); 
assign P2_ADD_394_U108 = ~P2_ADD_394_U28; 
assign P2_ADD_394_U157 = ~(P2_ADD_394_U28 & P2_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P2_R2267_U43 = ~(P2_R2267_U156 & P2_R2267_U155); 
assign P2_R2267_U89 = ~P2_R2267_U23; 
assign P2_R2267_U143 = ~(P2_U3644 & P2_R2267_U23); 
assign P1_R2027_U67 = ~(P1_R2027_U174 & P1_R2027_U173); 
assign P1_R2027_U68 = ~(P1_R2027_U176 & P1_R2027_U175); 
assign P1_R2027_U116 = ~P1_R2027_U43; 
assign P1_R2027_U133 = ~P1_R2027_U103; 
assign P1_R2027_U170 = ~(P1_R2027_U43 & P1_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P1_R2027_U171 = ~(P1_R2027_U103 & P1_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P1_R2182_U24 = ~(P1_R2182_U64 & P1_R2182_U63); 
assign P1_R2182_U25 = ~(P1_R2182_U66 & P1_R2182_U65); 
assign P1_R2182_U40 = ~(P1_U2733 & P1_R2182_U56); 
assign P1_R2182_U72 = ~(P1_R2182_U56 & P1_R2182_U23); 
assign P1_R2144_U112 = ~(P1_R2144_U189 & P1_R2144_U188 & P1_R2144_U15); 
assign P1_R2144_U192 = ~(P1_R2144_U191 & P1_R2144_U190); 
assign P1_R2358_U430 = ~(P1_R2358_U429 & P1_R2358_U428); 
assign P1_R2358_U479 = ~(P1_R2358_U478 & P1_R2358_U477); 
assign P1_R2358_U480 = ~(P1_U2352 & P1_R2358_U162); 
assign P1_R2358_U482 = ~(P1_U2352 & P1_R2358_U162); 
assign P1_R2099_U39 = ~(P1_R2099_U219 & P1_R2099_U218); 
assign P1_R2099_U40 = ~(P1_R2099_U221 & P1_R2099_U220); 
assign P1_R2099_U158 = ~P1_R2099_U110; 
assign P1_R2099_U159 = ~P1_R2099_U9; 
assign P1_R2099_U215 = ~(P1_R2099_U27 & P1_R2099_U9); 
assign P1_R2099_U217 = ~(P1_R2099_U29 & P1_R2099_U110); 
assign P1_R2167_U49 = ~(P1_R2167_U45 & P1_R2167_U15); 
assign P1_R2167_U50 = ~(P1_U2356 & P1_R2167_U48); 
assign P1_R2337_U88 = ~(P1_R2337_U176 & P1_R2337_U175); 
assign P1_R2337_U105 = ~P1_R2337_U28; 
assign P1_R2337_U173 = ~(P1_R2337_U28 & P1_PHYADDRPOINTER_REG_14__SCAN_IN); 
assign P1_R2096_U88 = ~(P1_R2096_U176 & P1_R2096_U175); 
assign P1_R2096_U105 = ~P1_R2096_U28; 
assign P1_R2096_U173 = ~(P1_R2096_U28 & P1_REIP_REG_14__SCAN_IN); 
assign P1_ADD_405_U69 = ~(P1_ADD_405_U140 & P1_ADD_405_U139); 
assign P1_ADD_405_U108 = ~P1_ADD_405_U28; 
assign P1_ADD_405_U157 = ~(P1_ADD_405_U28 & P1_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P1_ADD_515_U69 = ~(P1_ADD_515_U138 & P1_ADD_515_U137); 
assign P1_ADD_515_U105 = ~P1_ADD_515_U28; 
assign P1_ADD_515_U155 = ~(P1_ADD_515_U28 & P1_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_U2601 = P3_U2392 & P3_U2352; 
assign P3_U2602 = P3_U2404 & P3_EBX_REG_31__SCAN_IN; 
assign P3_U2637 = ~(P3_U7370 & P3_U7369); 
assign P3_U2827 = ~(P3_U6432 & P3_U6431 & P3_U6430 & P3_U6429 & P3_U3957); 
assign P3_U3284 = ~(P3_U7972 & P3_U7971); 
assign P3_U4002 = P3_U6857 & P3_U6856; 
assign P3_U4003 = P3_U6861 & P3_U6860; 
assign P3_U4004 = P3_U6865 & P3_U6864; 
assign P3_U4005 = P3_U6869 & P3_U6868; 
assign P3_U4006 = P3_U6873 & P3_U6872; 
assign P3_U4007 = P3_U6877 & P3_U6876; 
assign P3_U4008 = P3_U6881 & P3_U6880; 
assign P3_U4009 = P3_U6885 & P3_U6884; 
assign P3_U4010 = P3_U6889 & P3_U6888; 
assign P3_U4011 = P3_U6893 & P3_U6892; 
assign P3_U4012 = P3_U6897 & P3_U6896; 
assign P3_U4013 = P3_U6901 & P3_U6900; 
assign P3_U4014 = P3_U6905 & P3_U6904; 
assign P3_U4015 = P3_U6907 & P3_U6909; 
assign P3_U4016 = P3_U6911 & P3_U6913; 
assign P3_U4017 = P3_U6915 & P3_U6917; 
assign P3_U4018 = P3_U6922 & P3_U6920; 
assign P3_U4019 = P3_U6927 & P3_U6925; 
assign P3_U4020 = P3_U6932 & P3_U6930; 
assign P3_U4021 = P3_U6937 & P3_U6935; 
assign P3_U4022 = P3_U6942 & P3_U6940; 
assign P3_U4023 = P3_U6947 & P3_U6945; 
assign P3_U4024 = P3_U6952 & P3_U6950; 
assign P3_U4025 = P3_U6957 & P3_U6955; 
assign P3_U4026 = P3_U6962 & P3_U6960; 
assign P3_U4027 = P3_U6967 & P3_U6965; 
assign P3_U4028 = P3_U6972 & P3_U6970; 
assign P3_U4029 = P3_U6977 & P3_U6975; 
assign P3_U4032 = P3_U7101 & P3_U7100; 
assign P3_U4036 = P3_U7111 & P3_U7110; 
assign P3_U4040 = P3_U7121 & P3_U7120; 
assign P3_U4044 = P3_U7131 & P3_U7130; 
assign P3_U4048 = P3_U7140 & P3_U7141; 
assign P3_U4053 = P3_U7150 & P3_U7151; 
assign P3_U4318 = ~P3_U3247; 
assign P3_U5542 = ~(P3_U5537 & P3_U3676); 
assign P3_U5553 = ~(P3_U7982 & P3_U7981 & P3_U3679); 
assign P3_U5566 = ~(P3_U5563 & P3_U3681); 
assign P3_U5573 = ~(P3_U7994 & P3_U7993 & P3_U5572); 
assign P3_U5653 = ~(P3_U2402 & P3_REIP_REG_0__SCAN_IN); 
assign P3_U5655 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P3_U5677 = ~(P3_U2402 & P3_REIP_REG_1__SCAN_IN); 
assign P3_U5679 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P3_U5701 = ~(P3_U2402 & P3_REIP_REG_2__SCAN_IN); 
assign P3_U5703 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P3_U5724 = ~(P3_U3715 & P3_U5706 & P3_U3718 & P3_U3714 & P3_U3721); 
assign P3_U5725 = ~(P3_U2402 & P3_REIP_REG_3__SCAN_IN); 
assign P3_U5727 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P3_U5747 = ~(P3_ADD_371_1212_U91 & P3_U2360); 
assign P3_U5749 = ~(P3_U2402 & P3_REIP_REG_4__SCAN_IN); 
assign P3_U5751 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P3_U5752 = ~(P3_ADD_360_1242_U89 & P3_U2395); 
assign P3_U5773 = ~(P3_U2402 & P3_REIP_REG_5__SCAN_IN); 
assign P3_U5775 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P3_U5797 = ~(P3_U2402 & P3_REIP_REG_6__SCAN_IN); 
assign P3_U5799 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P3_U5821 = ~(P3_U2402 & P3_REIP_REG_7__SCAN_IN); 
assign P3_U5823 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_U5845 = ~(P3_U2402 & P3_REIP_REG_8__SCAN_IN); 
assign P3_U5847 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_U5869 = ~(P3_U2402 & P3_REIP_REG_9__SCAN_IN); 
assign P3_U5871 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_U5893 = ~(P3_U2402 & P3_REIP_REG_10__SCAN_IN); 
assign P3_U5895 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P3_U5917 = ~(P3_U2402 & P3_REIP_REG_11__SCAN_IN); 
assign P3_U5919 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_U5922 = ~(P3_ADD_558_U93 & P3_U3220); 
assign P3_U5923 = ~(P3_ADD_553_U93 & P3_U4298); 
assign P3_U5924 = ~(P3_ADD_547_U93 & P3_U4299); 
assign P3_U5927 = ~(P3_ADD_531_U93 & P3_U2354); 
assign P3_U5935 = ~(P3_ADD_385_U93 & P3_U2358); 
assign P3_U5936 = ~(P3_ADD_380_U93 & P3_U2359); 
assign P3_U5937 = ~(P3_ADD_349_U93 & P3_U4306); 
assign P3_U5938 = ~(P3_ADD_344_U93 & P3_U2362); 
assign P3_U5941 = ~(P3_U2402 & P3_REIP_REG_12__SCAN_IN); 
assign P3_U5943 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P3_U5949 = ~(P3_ADD_541_U88 & P3_U4300); 
assign P3_U5950 = ~(P3_ADD_536_U88 & P3_U4301); 
assign P3_U5953 = ~(P3_ADD_515_U88 & P3_U4302); 
assign P3_U5954 = ~(P3_ADD_494_U88 & P3_U2356); 
assign P3_U5955 = ~(P3_ADD_476_U88 & P3_U4303); 
assign P3_U5956 = ~(P3_ADD_441_U88 & P3_U4304); 
assign P3_U5957 = ~(P3_ADD_405_U88 & P3_U4305); 
assign P3_U5958 = ~(P3_ADD_394_U88 & P3_U2357); 
assign P3_U5965 = ~(P3_U2402 & P3_REIP_REG_13__SCAN_IN); 
assign P3_U5967 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_U5989 = ~(P3_U2402 & P3_REIP_REG_14__SCAN_IN); 
assign P3_U5991 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_U6013 = ~(P3_U2402 & P3_REIP_REG_15__SCAN_IN); 
assign P3_U6015 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_U6037 = ~(P3_U2402 & P3_REIP_REG_16__SCAN_IN); 
assign P3_U6039 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_U6061 = ~(P3_U2402 & P3_REIP_REG_17__SCAN_IN); 
assign P3_U6063 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_U6085 = ~(P3_U2402 & P3_REIP_REG_18__SCAN_IN); 
assign P3_U6087 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_U6109 = ~(P3_U2402 & P3_REIP_REG_19__SCAN_IN); 
assign P3_U6111 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_U6133 = ~(P3_U2402 & P3_REIP_REG_20__SCAN_IN); 
assign P3_U6135 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_U6157 = ~(P3_U2402 & P3_REIP_REG_21__SCAN_IN); 
assign P3_U6159 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_U6168 = ~(P3_ADD_526_U68 & P3_U2355); 
assign P3_U6181 = ~(P3_U2402 & P3_REIP_REG_22__SCAN_IN); 
assign P3_U6183 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_U6192 = ~(P3_ADD_526_U67 & P3_U2355); 
assign P3_U6205 = ~(P3_U2402 & P3_REIP_REG_23__SCAN_IN); 
assign P3_U6207 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_U6229 = ~(P3_U2402 & P3_REIP_REG_24__SCAN_IN); 
assign P3_U6231 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_U6253 = ~(P3_U2402 & P3_REIP_REG_25__SCAN_IN); 
assign P3_U6255 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_U6277 = ~(P3_U2402 & P3_REIP_REG_26__SCAN_IN); 
assign P3_U6279 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_U6301 = ~(P3_U2402 & P3_REIP_REG_27__SCAN_IN); 
assign P3_U6303 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_U6325 = ~(P3_U2402 & P3_REIP_REG_28__SCAN_IN); 
assign P3_U6327 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_U6349 = ~(P3_U2402 & P3_REIP_REG_29__SCAN_IN); 
assign P3_U6351 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_U6373 = ~(P3_U2402 & P3_REIP_REG_30__SCAN_IN); 
assign P3_U6375 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_U6397 = ~(P3_U2402 & P3_REIP_REG_31__SCAN_IN); 
assign P3_U6398 = ~(P3_U5631 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_U6443 = ~(P3_U2387 & P3_ADD_371_1212_U91); 
assign P3_U6447 = ~(P3_U2396 & P3_ADD_360_1242_U89); 
assign P3_U6509 = ~(P3_ADD_318_U88 & P3_U2398); 
assign P3_U6514 = ~(P3_ADD_339_U88 & P3_U2388); 
assign P3_U6518 = ~(P3_ADD_315_U84 & P3_U2397); 
assign P3_U6854 = ~(P3_U2446 & BUF2_REG_0__SCAN_IN); 
assign P3_U6858 = ~(P3_U2446 & BUF2_REG_1__SCAN_IN); 
assign P3_U6862 = ~(P3_U2446 & BUF2_REG_2__SCAN_IN); 
assign P3_U6866 = ~(P3_U2446 & BUF2_REG_3__SCAN_IN); 
assign P3_U6870 = ~(P3_U2446 & BUF2_REG_4__SCAN_IN); 
assign P3_U6874 = ~(P3_U2446 & BUF2_REG_5__SCAN_IN); 
assign P3_U6878 = ~(P3_U2446 & BUF2_REG_6__SCAN_IN); 
assign P3_U6882 = ~(P3_U2446 & BUF2_REG_7__SCAN_IN); 
assign P3_U6886 = ~(P3_U2446 & BUF2_REG_8__SCAN_IN); 
assign P3_U6890 = ~(P3_U2446 & BUF2_REG_9__SCAN_IN); 
assign P3_U6894 = ~(P3_U2446 & BUF2_REG_10__SCAN_IN); 
assign P3_U6898 = ~(P3_U2446 & BUF2_REG_11__SCAN_IN); 
assign P3_U6902 = ~(P3_U2446 & BUF2_REG_12__SCAN_IN); 
assign P3_U6906 = ~(P3_U2446 & BUF2_REG_13__SCAN_IN); 
assign P3_U6910 = ~(P3_U2446 & BUF2_REG_14__SCAN_IN); 
assign P3_U6914 = ~(P3_U2446 & BUF2_REG_15__SCAN_IN); 
assign P3_U6918 = ~(P3_U2448 & BUF2_REG_0__SCAN_IN); 
assign P3_U6919 = ~(P3_U2444 & BUF2_REG_16__SCAN_IN); 
assign P3_U6923 = ~(P3_U2448 & BUF2_REG_1__SCAN_IN); 
assign P3_U6924 = ~(P3_U2444 & BUF2_REG_17__SCAN_IN); 
assign P3_U6928 = ~(P3_U2448 & BUF2_REG_2__SCAN_IN); 
assign P3_U6929 = ~(P3_U2444 & BUF2_REG_18__SCAN_IN); 
assign P3_U6933 = ~(P3_U2448 & BUF2_REG_3__SCAN_IN); 
assign P3_U6934 = ~(P3_U2444 & BUF2_REG_19__SCAN_IN); 
assign P3_U6938 = ~(P3_U2448 & BUF2_REG_4__SCAN_IN); 
assign P3_U6939 = ~(P3_U2444 & BUF2_REG_20__SCAN_IN); 
assign P3_U6943 = ~(P3_U2448 & BUF2_REG_5__SCAN_IN); 
assign P3_U6944 = ~(P3_U2444 & BUF2_REG_21__SCAN_IN); 
assign P3_U6948 = ~(P3_U2448 & BUF2_REG_6__SCAN_IN); 
assign P3_U6949 = ~(P3_U2444 & BUF2_REG_22__SCAN_IN); 
assign P3_U6951 = ~(P3_ADD_546_U68 & P3_U2400); 
assign P3_U6953 = ~(P3_U2448 & BUF2_REG_7__SCAN_IN); 
assign P3_U6954 = ~(P3_U2444 & BUF2_REG_23__SCAN_IN); 
assign P3_U6956 = ~(P3_ADD_546_U67 & P3_U2400); 
assign P3_U6958 = ~(P3_U2448 & BUF2_REG_8__SCAN_IN); 
assign P3_U6959 = ~(P3_U2444 & BUF2_REG_24__SCAN_IN); 
assign P3_U6963 = ~(P3_U2448 & BUF2_REG_9__SCAN_IN); 
assign P3_U6964 = ~(P3_U2444 & BUF2_REG_25__SCAN_IN); 
assign P3_U6968 = ~(P3_U2448 & BUF2_REG_10__SCAN_IN); 
assign P3_U6969 = ~(P3_U2444 & BUF2_REG_26__SCAN_IN); 
assign P3_U6973 = ~(P3_U2448 & BUF2_REG_11__SCAN_IN); 
assign P3_U6974 = ~(P3_U2444 & BUF2_REG_27__SCAN_IN); 
assign P3_U6978 = ~(P3_U2448 & BUF2_REG_12__SCAN_IN); 
assign P3_U6979 = ~(P3_U2444 & BUF2_REG_28__SCAN_IN); 
assign P3_U6983 = ~(P3_U2448 & BUF2_REG_13__SCAN_IN); 
assign P3_U6984 = ~(P3_U2444 & BUF2_REG_29__SCAN_IN); 
assign P3_U6988 = ~(P3_U2448 & BUF2_REG_14__SCAN_IN); 
assign P3_U6989 = ~(P3_U2444 & BUF2_REG_30__SCAN_IN); 
assign P3_U6993 = ~(P3_U2444 & BUF2_REG_31__SCAN_IN); 
assign P3_U7065 = ~(P3_ADD_552_U68 & P3_U2399); 
assign P3_U7068 = ~(P3_ADD_552_U67 & P3_U2399); 
assign P3_U7102 = ~(P3_U2405 & P3_REIP_REG_0__SCAN_IN); 
assign P3_U7112 = ~(P3_ADD_430_U4 & P3_U2405); 
assign P3_U7122 = ~(P3_ADD_430_U71 & P3_U2405); 
assign P3_U7132 = ~(P3_ADD_430_U68 & P3_U2405); 
assign P3_U7142 = ~(P3_ADD_430_U67 & P3_U2405); 
assign P3_U7152 = ~(P3_ADD_430_U66 & P3_U2405); 
assign P3_U7160 = ~(P3_ADD_430_U65 & P3_U2405); 
assign P3_U7168 = ~(P3_ADD_430_U64 & P3_U2405); 
assign P3_U7176 = ~(P3_ADD_430_U63 & P3_U2405); 
assign P3_U7184 = ~(P3_ADD_430_U62 & P3_U2405); 
assign P3_U7192 = ~(P3_ADD_430_U91 & P3_U2405); 
assign P3_U7200 = ~(P3_ADD_430_U90 & P3_U2405); 
assign P3_U7208 = ~(P3_ADD_430_U89 & P3_U2405); 
assign P3_U7216 = ~(P3_ADD_430_U88 & P3_U2405); 
assign P3_U7908 = ~(P3_U2404 & P3_U3256); 
assign P3_U7909 = ~(P3_U2392 & P3_U7096); 
assign P3_U8018 = ~(P3_U7368 & P3_U4617); 
assign P2_U2473 = P2_R2099_U94 & P2_U3324; 
assign P2_U2701 = ~(P2_U7161 & P2_U7162 & P2_U7160); 
assign P2_U3322 = ~P2_R2099_U96; 
assign P2_U3641 = ~(P2_U8336 & P2_U8335); 
assign P2_U5618 = ~(P2_R2099_U96 & P2_U5603); 
assign P2_U5629 = ~(P2_U3888 & P2_U5628); 
assign P2_U7149 = ~(P2_U4467 & P2_R2099_U96); 
assign P2_U8328 = ~(P2_U3242 & P2_R2267_U43); 
assign P2_U8409 = ~(P2_R2337_U86 & P2_U3284); 
assign P1_U2438 = P1_R2182_U42 & P1_R2182_U25; 
assign P1_U2440 = P1_R2182_U25 & P1_U3317; 
assign P1_U2441 = ~(P1_R2182_U42 | P1_R2182_U25); 
assign P1_U2667 = ~(P1_U6759 & P1_U4006); 
assign P1_U2670 = ~(P1_U6824 & P1_U6823 & P1_U4021 & P1_U6820); 
assign P1_U2766 = ~(P1_U6939 & P1_U6938 & P1_U6940); 
assign P1_U3316 = ~P1_R2182_U25; 
assign P1_U3467 = P1_U2427 & P1_U4215 & P1_R2182_U24; 
assign P1_U3488 = P1_R2182_U24 & P1_U4215; 
assign P1_U5503 = ~(P1_R2182_U25 & P1_U7509); 
assign P1_U5514 = ~(P1_U3749 & P1_U5512); 
assign P1_U5528 = ~(P1_U2427 & P1_U5525); 
assign P1_U5543 = ~(P1_R2182_U25 & P1_U5538); 
assign P1_U6763 = ~(P1_R2182_U24 & P1_U6746); 
assign P1_U6775 = ~(P1_R2182_U25 & P1_U6746); 
assign P1_U6849 = ~(P1_R2337_U88 & P1_U2352); 
assign P1_U6937 = ~(P1_R2182_U25 & P1_U3294); 
assign P3_ADD_526_U46 = ~(P3_ADD_526_U93 & P3_ADD_526_U116); 
assign P3_ADD_526_U102 = ~(P3_ADD_526_U116 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_526_U169 = ~(P3_ADD_526_U116 & P3_ADD_526_U42); 
assign P3_ADD_526_U172 = ~(P3_ADD_526_U133 & P3_ADD_526_U38); 
assign P3_ADD_552_U46 = ~(P3_ADD_552_U93 & P3_ADD_552_U116); 
assign P3_ADD_552_U102 = ~(P3_ADD_552_U116 & P3_EBX_REG_25__SCAN_IN); 
assign P3_ADD_552_U169 = ~(P3_ADD_552_U116 & P3_ADD_552_U42); 
assign P3_ADD_552_U172 = ~(P3_ADD_552_U133 & P3_ADD_552_U38); 
assign P3_ADD_546_U46 = ~(P3_ADD_546_U93 & P3_ADD_546_U116); 
assign P3_ADD_546_U102 = ~(P3_ADD_546_U116 & P3_EAX_REG_25__SCAN_IN); 
assign P3_ADD_546_U169 = ~(P3_ADD_546_U116 & P3_ADD_546_U42); 
assign P3_ADD_546_U172 = ~(P3_ADD_546_U133 & P3_ADD_546_U38); 
assign P3_ADD_391_1180_U19 = ~(P3_ADD_391_1180_U38 & P3_ADD_391_1180_U37); 
assign P3_ADD_391_1180_U34 = ~P3_ADD_391_1180_U27; 
assign P3_ADD_391_1180_U35 = ~(P3_U2620 & P3_ADD_391_1180_U27); 
assign P3_ADD_476_U30 = ~(P3_ADD_476_U105 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_476_U174 = ~(P3_ADD_476_U105 & P3_ADD_476_U29); 
assign P3_ADD_531_U31 = ~(P3_ADD_531_U109 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_531_U183 = ~(P3_ADD_531_U109 & P3_ADD_531_U30); 
assign P3_SUB_320_U7 = P3_SUB_320_U124 & P3_SUB_320_U29; 
assign P3_SUB_320_U79 = ~P3_ADD_318_U88; 
assign P3_SUB_320_U94 = ~P3_SUB_320_U29; 
assign P3_SUB_320_U156 = ~(P3_ADD_318_U88 & P3_SUB_320_U29); 
assign P3_ADD_318_U30 = ~(P3_ADD_318_U105 & P3_PHYADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_318_U174 = ~(P3_ADD_318_U105 & P3_ADD_318_U29); 
assign P3_ADD_315_U30 = ~(P3_ADD_315_U102 & P3_PHYADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_315_U166 = ~(P3_ADD_315_U102 & P3_ADD_315_U29); 
assign P3_ADD_360_1242_U110 = ~(P3_ADD_360_1242_U141 & P3_ADD_360_1242_U140); 
assign P3_ADD_360_1242_U202 = ~(P3_ADD_360_1242_U36 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_360_1242_U204 = ~(P3_ADD_360_1242_U36 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_360_1242_U214 = ~(P3_ADD_360_1242_U111 & P3_ADD_360_1242_U112); 
assign P3_ADD_360_1242_U215 = ~(P3_ADD_360_1242_U138 & P3_ADD_360_1242_U213); 
assign P3_ADD_467_U30 = ~(P3_ADD_467_U105 & P3_REIP_REG_14__SCAN_IN); 
assign P3_ADD_467_U174 = ~(P3_ADD_467_U105 & P3_ADD_467_U29); 
assign P3_ADD_430_U30 = ~(P3_ADD_430_U105 & P3_REIP_REG_14__SCAN_IN); 
assign P3_ADD_430_U174 = ~(P3_ADD_430_U105 & P3_ADD_430_U29); 
assign P3_ADD_380_U31 = ~(P3_ADD_380_U109 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_380_U183 = ~(P3_ADD_380_U109 & P3_ADD_380_U30); 
assign P3_ADD_344_U31 = ~(P3_ADD_344_U109 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_344_U183 = ~(P3_ADD_344_U109 & P3_ADD_344_U30); 
assign P3_LT_563_U28 = ~(P3_LT_563_U14 & P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P3_ADD_339_U30 = ~(P3_ADD_339_U105 & P3_PHYADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_339_U174 = ~(P3_ADD_339_U105 & P3_ADD_339_U29); 
assign P3_ADD_541_U30 = ~(P3_ADD_541_U105 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_541_U174 = ~(P3_ADD_541_U105 & P3_ADD_541_U29); 
assign P3_SUB_357_1258_U73 = ~(P3_SUB_357_1258_U333 & P3_SUB_357_1258_U332); 
assign P3_SUB_357_1258_U174 = ~P3_SUB_357_1258_U119; 
assign P3_SUB_357_1258_U300 = ~(P3_SUB_357_1258_U175 & P3_SUB_357_1258_U119); 
assign P3_SUB_357_1258_U325 = ~(P3_SUB_357_1258_U118 & P3_SUB_357_1258_U119); 
assign P3_ADD_515_U30 = ~(P3_ADD_515_U105 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_515_U174 = ~(P3_ADD_515_U105 & P3_ADD_515_U29); 
assign P3_ADD_394_U30 = ~(P3_ADD_394_U108 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_394_U178 = ~(P3_ADD_394_U108 & P3_ADD_394_U29); 
assign P3_SUB_414_U13 = P3_SUB_414_U112 & P3_SUB_414_U35; 
assign P3_SUB_414_U36 = ~(P3_SUB_414_U41 & P3_SUB_414_U65 & P3_SUB_414_U100); 
assign P3_SUB_414_U109 = ~(P3_SUB_414_U100 & P3_SUB_414_U65); 
assign P3_SUB_414_U143 = ~(P3_SUB_414_U100 & P3_SUB_414_U65); 
assign P3_ADD_441_U30 = ~(P3_ADD_441_U105 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_441_U174 = ~(P3_ADD_441_U105 & P3_ADD_441_U29); 
assign P3_ADD_349_U31 = ~(P3_ADD_349_U109 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_349_U183 = ~(P3_ADD_349_U109 & P3_ADD_349_U30); 
assign P3_ADD_405_U30 = ~(P3_ADD_405_U108 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_405_U178 = ~(P3_ADD_405_U108 & P3_ADD_405_U29); 
assign P3_ADD_553_U31 = ~(P3_ADD_553_U109 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_553_U183 = ~(P3_ADD_553_U109 & P3_ADD_553_U30); 
assign P3_ADD_558_U31 = ~(P3_ADD_558_U109 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_558_U183 = ~(P3_ADD_558_U109 & P3_ADD_558_U30); 
assign P3_ADD_385_U31 = ~(P3_ADD_385_U109 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_385_U183 = ~(P3_ADD_385_U109 & P3_ADD_385_U30); 
assign P3_ADD_547_U31 = ~(P3_ADD_547_U109 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_547_U183 = ~(P3_ADD_547_U109 & P3_ADD_547_U30); 
assign P3_ADD_371_1212_U19 = P3_ADD_371_1212_U155 & P3_ADD_371_1212_U152; 
assign P3_ADD_371_1212_U139 = ~P3_ADD_371_1212_U115; 
assign P3_ADD_371_1212_U141 = ~(P3_ADD_371_1212_U140 & P3_ADD_371_1212_U115); 
assign P3_ADD_371_1212_U213 = ~(P3_ADD_371_1212_U39 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_371_1212_U215 = ~(P3_ADD_371_1212_U39 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_371_1212_U225 = ~(P3_ADD_371_1212_U114 & P3_ADD_371_1212_U115); 
assign P3_ADD_494_U30 = ~(P3_ADD_494_U105 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_494_U174 = ~(P3_ADD_494_U105 & P3_ADD_494_U29); 
assign P3_ADD_536_U30 = ~(P3_ADD_536_U105 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_536_U174 = ~(P3_ADD_536_U105 & P3_ADD_536_U29); 
assign P3_ADD_402_1132_U19 = ~(P3_ADD_402_1132_U38 & P3_ADD_402_1132_U37); 
assign P3_ADD_402_1132_U34 = ~P3_ADD_402_1132_U27; 
assign P3_ADD_402_1132_U35 = ~(P3_U2620 & P3_ADD_402_1132_U27); 
assign P2_R2099_U97 = ~(P2_R2099_U118 & P2_R2099_U117); 
assign P2_R2099_U167 = ~(P2_R2099_U115 & P2_R2099_U165); 
assign P2_ADD_391_1196_U29 = ~P2_R2096_U74; 
assign P2_ADD_402_1132_U19 = ~(P2_ADD_402_1132_U38 & P2_ADD_402_1132_U37); 
assign P2_ADD_402_1132_U34 = ~P2_ADD_402_1132_U27; 
assign P2_ADD_402_1132_U35 = ~(P2_U2598 & P2_ADD_402_1132_U27); 
assign P2_R2182_U62 = ~P2_U2684; 
assign P2_R2182_U69 = ~(P2_R2182_U305 & P2_R2182_U304); 
assign P2_R2182_U112 = P2_R2182_U239 & P2_R2182_U238; 
assign P2_R2182_U122 = ~(P2_U2680 & P2_R2182_U121); 
assign P2_R2182_U175 = P2_U2684 | P2_U2660; 
assign P2_R2182_U177 = ~(P2_U2660 & P2_U2684); 
assign P2_R2182_U189 = ~(P2_U2680 & P2_R2182_U121); 
assign P2_R2182_U232 = ~(P2_U2684 & P2_R2182_U63); 
assign P2_R2182_U234 = ~(P2_U2684 & P2_R2182_U63); 
assign P2_R2182_U242 = ~(P2_R2182_U241 & P2_R2182_U240); 
assign P2_R2182_U279 = ~(P2_R2182_U121 & P2_R2182_U47); 
assign P2_R2167_U12 = ~P2_U2711; 
assign P2_R2167_U16 = ~P2_U2709; 
assign P2_R2167_U26 = ~(P2_R2167_U24 & P2_R2167_U25 & P2_R2167_U23); 
assign P2_R2167_U30 = ~(P2_U2711 & P2_R2167_U11); 
assign P2_R2167_U33 = ~(P2_U2703 & P2_R2167_U13); 
assign P2_R2167_U36 = ~(P2_U2709 & P2_R2167_U15); 
assign P2_R2027_U31 = ~(P2_R2027_U109 & P2_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P2_R2027_U183 = ~(P2_R2027_U109 & P2_R2027_U30); 
assign P2_R2337_U31 = ~(P2_R2337_U106 & P2_PHYADDRPOINTER_REG_15__SCAN_IN); 
assign P2_R2337_U172 = ~(P2_R2337_U106 & P2_R2337_U30); 
assign P2_R2219_U25 = ~(P2_R2219_U91 & P2_R2219_U90); 
assign P2_R2219_U65 = ~P2_R2219_U39; 
assign P2_R2219_U68 = ~(P2_R2219_U67 & P2_R2219_U39); 
assign P2_R2219_U86 = ~(P2_R2219_U32 & P2_R2219_U39); 
assign P2_R2096_U103 = ~(P2_R2096_U134 & P2_R2096_U133); 
assign P2_R2096_U195 = ~(P2_R2096_U131 & P2_R2096_U193); 
assign P2_R1957_U7 = P2_R1957_U124 & P2_R1957_U28; 
assign P2_R1957_U79 = ~P2_U3678; 
assign P2_R1957_U94 = ~P2_R1957_U28; 
assign P2_R1957_U156 = ~(P2_U3678 & P2_R1957_U28); 
assign P2_ADD_394_U30 = ~(P2_ADD_394_U108 & P2_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P2_ADD_394_U158 = ~(P2_ADD_394_U108 & P2_ADD_394_U29); 
assign P2_R2267_U29 = ~P2_U3643; 
assign P2_R2267_U59 = ~P2_U3642; 
assign P2_R2267_U100 = ~(P2_R2267_U89 & P2_R2267_U64); 
assign P2_R2267_U144 = ~(P2_R2267_U89 & P2_R2267_U64); 
assign P1_R2027_U46 = ~(P1_R2027_U93 & P1_R2027_U116); 
assign P1_R2027_U102 = ~(P1_R2027_U116 & P1_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P1_R2027_U169 = ~(P1_R2027_U116 & P1_R2027_U42); 
assign P1_R2027_U172 = ~(P1_R2027_U133 & P1_R2027_U38); 
assign P1_R2182_U27 = ~(P1_R2182_U72 & P1_R2182_U71); 
assign P1_R2182_U57 = ~P1_R2182_U40; 
assign P1_R2182_U67 = ~(P1_U2732 & P1_R2182_U40); 
assign P1_R2144_U73 = ~P1_U2767; 
assign P1_R2144_U113 = ~(P1_U2752 & P1_R2144_U192); 
assign P1_R2144_U115 = ~(P1_U2355 & P1_R2144_U112); 
assign P1_R2144_U129 = ~(P1_U2355 & P1_R2144_U112); 
assign P1_R2144_U186 = ~(P1_U2767 & P1_R2144_U12); 
assign P1_R2358_U12 = P1_R2358_U481 & P1_R2358_U480; 
assign P1_R2358_U149 = ~P1_U2671; 
assign P1_R2358_U160 = ~P1_U2616; 
assign P1_R2358_U426 = ~(P1_U2671 & P1_R2358_U23); 
assign P1_R2358_U432 = ~(P1_U2671 & P1_R2358_U23); 
assign P1_R2358_U470 = ~(P1_U2616 & P1_R2358_U23); 
assign P1_R2358_U484 = ~(P1_R2358_U483 & P1_R2358_U482); 
assign P1_R2358_U486 = ~(P1_U2616 & P1_R2358_U23); 
assign P1_R2099_U10 = ~(P1_R2099_U91 & P1_R2099_U159); 
assign P1_R2099_U109 = ~(P1_R2099_U159 & P1_R2099_U27); 
assign P1_R2099_U214 = ~(P1_R2099_U184 & P1_R2099_U159); 
assign P1_R2099_U216 = ~(P1_R2099_U158 & P1_R2099_U208); 
assign P1_R2167_U17 = ~(P1_R2167_U50 & P1_R2167_U49); 
assign P1_R2337_U30 = ~(P1_R2337_U105 & P1_PHYADDRPOINTER_REG_14__SCAN_IN); 
assign P1_R2337_U174 = ~(P1_R2337_U105 & P1_R2337_U29); 
assign P1_R2096_U30 = ~(P1_R2096_U105 & P1_REIP_REG_14__SCAN_IN); 
assign P1_R2096_U174 = ~(P1_R2096_U105 & P1_R2096_U29); 
assign P1_ADD_405_U30 = ~(P1_ADD_405_U108 & P1_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P1_ADD_405_U158 = ~(P1_ADD_405_U108 & P1_ADD_405_U29); 
assign P1_ADD_515_U30 = ~(P1_ADD_515_U105 & P1_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P1_ADD_515_U156 = ~(P1_ADD_515_U105 & P1_ADD_515_U29); 
assign P3_U2680 = ~(P3_U7069 & P3_U7067 & P3_U7068); 
assign P3_U2681 = ~(P3_U7066 & P3_U7064 & P3_U7065); 
assign P3_U2712 = ~(P3_U6954 & P3_U6953 & P3_U4025 & P3_U6956); 
assign P3_U2713 = ~(P3_U6949 & P3_U6948 & P3_U4024 & P3_U6951); 
assign P3_U2714 = ~(P3_U6944 & P3_U6943 & P3_U4023 & P3_U6946); 
assign P3_U2715 = ~(P3_U6939 & P3_U6938 & P3_U4022 & P3_U6941); 
assign P3_U2716 = ~(P3_U6934 & P3_U6933 & P3_U4021 & P3_U6936); 
assign P3_U2717 = ~(P3_U6929 & P3_U6928 & P3_U4020 & P3_U6931); 
assign P3_U2718 = ~(P3_U6924 & P3_U6923 & P3_U4019 & P3_U6926); 
assign P3_U2719 = ~(P3_U6919 & P3_U6918 & P3_U4018 & P3_U6921); 
assign P3_U2720 = ~(P3_U6914 & P3_U4017 & P3_U6916); 
assign P3_U2721 = ~(P3_U6910 & P3_U4016 & P3_U6912); 
assign P3_U2722 = ~(P3_U6906 & P3_U4015 & P3_U6908); 
assign P3_U2723 = ~(P3_U6903 & P3_U6902 & P3_U4014); 
assign P3_U2724 = ~(P3_U6899 & P3_U6898 & P3_U4013); 
assign P3_U2725 = ~(P3_U6895 & P3_U6894 & P3_U4012); 
assign P3_U2726 = ~(P3_U6891 & P3_U6890 & P3_U4011); 
assign P3_U2727 = ~(P3_U6887 & P3_U6886 & P3_U4010); 
assign P3_U2728 = ~(P3_U6883 & P3_U6882 & P3_U4009); 
assign P3_U2729 = ~(P3_U6879 & P3_U6878 & P3_U4008); 
assign P3_U2730 = ~(P3_U6875 & P3_U6874 & P3_U4007); 
assign P3_U2731 = ~(P3_U6871 & P3_U6870 & P3_U4006); 
assign P3_U2732 = ~(P3_U6867 & P3_U6866 & P3_U4005); 
assign P3_U2733 = ~(P3_U6863 & P3_U6862 & P3_U4004); 
assign P3_U2734 = ~(P3_U6859 & P3_U6858 & P3_U4003); 
assign P3_U2735 = ~(P3_U6855 & P3_U6854 & P3_U4002); 
assign P3_U3295 = ~(P3_U8019 & P3_U8018); 
assign P3_U3729 = P3_U3728 & P3_U3727 & P3_U5747; 
assign P3_U3730 = P3_U3731 & P3_U5752; 
assign P3_U3783 = P3_U5924 & P3_U5923; 
assign P3_U3785 = P3_U5926 & P3_U5925 & P3_U5927 & P3_U3784; 
assign P3_U3787 = P3_U5938 & P3_U5937 & P3_U5936 & P3_U5935; 
assign P3_U3791 = P3_U5953 & P3_U5952; 
assign P3_U3793 = P3_U5955 & P3_U5954 & P3_U5956 & P3_U5958 & P3_U5957; 
assign P3_U3803 = P3_U5991 & P3_U5989; 
assign P3_U3811 = P3_U6015 & P3_U6013; 
assign P3_U3845 = P3_U6135 & P3_U6133; 
assign P3_U3853 = P3_U6159 & P3_U6157; 
assign P3_U3863 = P3_U6183 & P3_U6181; 
assign P3_U3873 = P3_U6207 & P3_U6205; 
assign P3_U3883 = P3_U6231 & P3_U6229; 
assign P3_U3893 = P3_U6255 & P3_U6253; 
assign P3_U3939 = P3_U6398 & P3_U3247; 
assign P3_U3958 = P3_U6442 & P3_U6441 & P3_U6444 & P3_U6443; 
assign P3_U5545 = ~(P3_U4340 & P3_U5542); 
assign P3_U5556 = ~(P3_U4340 & P3_U5553); 
assign P3_U5569 = ~(P3_U4340 & P3_U5566); 
assign P3_U5575 = ~(P3_U4340 & P3_U5573); 
assign P3_U5654 = ~(P3_U4318 & P3_U5652); 
assign P3_U5678 = ~(P3_U4318 & P3_U5676); 
assign P3_U5702 = ~(P3_U4318 & P3_U5700); 
assign P3_U5726 = ~(P3_U4318 & P3_U5724); 
assign P3_U5771 = ~(P3_ADD_371_1212_U19 & P3_U2360); 
assign P3_U5777 = ~(P3_SUB_357_1258_U73 & P3_U2393); 
assign P3_U6451 = ~(P3_U2387 & P3_ADD_371_1212_U19); 
assign P3_U6456 = ~(P3_U2394 & P3_SUB_357_1258_U73); 
assign P3_U6985 = ~(P3_ADD_391_1180_U19 & P3_U2411); 
assign P3_U7085 = ~(P3_ADD_402_1132_U19 & P3_U2408); 
assign P3_U7097 = ~(P3_U2602 & P3_EBX_REG_0__SCAN_IN); 
assign P3_U7098 = ~(P3_U2601 & P3_REIP_REG_0__SCAN_IN); 
assign P3_U7107 = ~(P3_SUB_414_U50 & P3_U2602); 
assign P3_U7108 = ~(P3_ADD_467_U4 & P3_U2601); 
assign P3_U7117 = ~(P3_SUB_414_U17 & P3_U2602); 
assign P3_U7118 = ~(P3_ADD_467_U71 & P3_U2601); 
assign P3_U7127 = ~(P3_SUB_414_U59 & P3_U2602); 
assign P3_U7128 = ~(P3_ADD_467_U68 & P3_U2601); 
assign P3_U7137 = ~(P3_SUB_414_U18 & P3_U2602); 
assign P3_U7138 = ~(P3_ADD_467_U67 & P3_U2601); 
assign P3_U7147 = ~(P3_SUB_414_U57 & P3_U2602); 
assign P3_U7148 = ~(P3_ADD_467_U66 & P3_U2601); 
assign P3_U7157 = ~(P3_SUB_414_U19 & P3_U2602); 
assign P3_U7158 = ~(P3_ADD_467_U65 & P3_U2601); 
assign P3_U7165 = ~(P3_SUB_414_U55 & P3_U2602); 
assign P3_U7166 = ~(P3_ADD_467_U64 & P3_U2601); 
assign P3_U7173 = ~(P3_SUB_414_U20 & P3_U2602); 
assign P3_U7174 = ~(P3_ADD_467_U63 & P3_U2601); 
assign P3_U7181 = ~(P3_SUB_414_U53 & P3_U2602); 
assign P3_U7182 = ~(P3_ADD_467_U62 & P3_U2601); 
assign P3_U7189 = ~(P3_SUB_414_U6 & P3_U2602); 
assign P3_U7190 = ~(P3_ADD_467_U91 & P3_U2601); 
assign P3_U7197 = ~(P3_SUB_414_U82 & P3_U2602); 
assign P3_U7198 = ~(P3_ADD_467_U90 & P3_U2601); 
assign P3_U7205 = ~(P3_SUB_414_U7 & P3_U2602); 
assign P3_U7206 = ~(P3_ADD_467_U89 & P3_U2601); 
assign P3_U7213 = ~(P3_SUB_414_U80 & P3_U2602); 
assign P3_U7214 = ~(P3_ADD_467_U88 & P3_U2601); 
assign P3_U7221 = ~(P3_SUB_414_U8 & P3_U2602); 
assign P3_U7229 = ~(P3_SUB_414_U78 & P3_U2602); 
assign P3_U7237 = ~(P3_SUB_414_U9 & P3_U2602); 
assign P3_U7245 = ~(P3_SUB_414_U76 & P3_U2602); 
assign P3_U7253 = ~(P3_SUB_414_U10 & P3_U2602); 
assign P3_U7261 = ~(P3_SUB_414_U74 & P3_U2602); 
assign P3_U7269 = ~(P3_SUB_414_U11 & P3_U2602); 
assign P3_U7277 = ~(P3_SUB_414_U70 & P3_U2602); 
assign P3_U7285 = ~(P3_SUB_414_U12 & P3_U2602); 
assign P3_U7293 = ~(P3_SUB_414_U68 & P3_U2602); 
assign P3_U7301 = ~(P3_SUB_414_U13 & P3_U2602); 
assign P3_U7910 = ~(P3_U7908 & P3_U4317 & P3_U7909); 
assign P3_U8047 = ~(P3_U5542 & P3_U4290); 
assign P3_U8049 = ~(P3_U5553 & P3_U4290); 
assign P3_U8051 = ~(P3_U5566 & P3_U4290); 
assign P3_U8053 = ~(P3_U5573 & P3_U4290); 
assign P2_U2683 = P2_ADD_402_1132_U19 & P2_U2355; 
assign P2_U2700 = ~(P2_U7150 & P2_U7151 & P2_U7149); 
assign P2_U2708 = P2_R2219_U25 & P2_U7723; 
assign P2_U3314 = ~P2_R2182_U69; 
assign P2_U3677 = ~(P2_U8410 & P2_U8409); 
assign P2_U5619 = ~(P2_U3885 & P2_U5618); 
assign P2_U5632 = ~(P2_U4466 & P2_U5629); 
assign P2_U5662 = ~(P2_R2182_U69 & P2_U5661); 
assign P2_U8333 = ~(P2_R2219_U25 & P2_U2617); 
assign P1_U2357 = P1_U5959 & P1_U3865 & P1_R2167_U17; 
assign P1_U2439 = P1_R2182_U42 & P1_U3316; 
assign P1_U2448 = P1_R2167_U17 & P1_U3284; 
assign P1_U2613 = ~(P1_U6847 & P1_U6848 & P1_U6849); 
assign P1_U2668 = ~(P1_U6767 & P1_U6766 & P1_U4008 & P1_U6763); 
assign P1_U2669 = ~(P1_U6779 & P1_U6778 & P1_U4010 & P1_U6775); 
assign P1_U2765 = ~(P1_U6936 & P1_U6935 & P1_U6937); 
assign P1_U3273 = ~P1_R2167_U17; 
assign P1_U3281 = ~(P1_R2167_U17 & P1_U4497); 
assign P1_U3299 = ~(P1_R2167_U17 & P1_STATE2_REG_3__SCAN_IN); 
assign P1_U4535 = ~(P1_U2438 & P1_U2442); 
assign P1_U4603 = ~(P1_U2443 & P1_U2438); 
assign P1_U4661 = ~(P1_U2444 & P1_U2438); 
assign P1_U4719 = ~(P1_U2445 & P1_U2438); 
assign P1_U4776 = ~(P1_U2440 & P1_U2442); 
assign P1_U4834 = ~(P1_U2440 & P1_U2443); 
assign P1_U4891 = ~(P1_U2440 & P1_U2444); 
assign P1_U4949 = ~(P1_U2440 & P1_U2445); 
assign P1_U5234 = ~(P1_U2441 & P1_U2442); 
assign P1_U5292 = ~(P1_U2441 & P1_U2443); 
assign P1_U5349 = ~(P1_U2441 & P1_U2444); 
assign P1_U5407 = ~(P1_U2441 & P1_U2445); 
assign P1_U5506 = ~(P1_U5503 & P1_U3747); 
assign P1_U5517 = ~(P1_U2427 & P1_U5514); 
assign P1_U6151 = ~(P1_U4200 & P1_U3283 & P1_R2167_U17); 
assign P1_U6361 = ~(P1_U4202 & P1_R2167_U17); 
assign P1_U6780 = ~(P1_R2182_U27 & P1_U6746); 
assign P1_U7501 = ~(P1_U7493 & P1_R2167_U17); 
assign P1_U7502 = ~(P1_U7493 & P1_U4201 & P1_R2167_U17); 
assign P1_U7681 = ~(P1_U4216 & P1_R2167_U17); 
assign P1_U7698 = ~(P1_R2167_U17 & P1_U7497); 
assign P1_U7743 = ~(P1_R2167_U17 & P1_U7611 & P1_U4432); 
assign P3_ADD_526_U65 = ~(P3_ADD_526_U170 & P3_ADD_526_U169); 
assign P3_ADD_526_U66 = ~(P3_ADD_526_U172 & P3_ADD_526_U171); 
assign P3_ADD_526_U122 = ~P3_ADD_526_U46; 
assign P3_ADD_526_U132 = ~P3_ADD_526_U102; 
assign P3_ADD_526_U166 = ~(P3_ADD_526_U46 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_526_U167 = ~(P3_ADD_526_U102 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_552_U65 = ~(P3_ADD_552_U170 & P3_ADD_552_U169); 
assign P3_ADD_552_U66 = ~(P3_ADD_552_U172 & P3_ADD_552_U171); 
assign P3_ADD_552_U122 = ~P3_ADD_552_U46; 
assign P3_ADD_552_U132 = ~P3_ADD_552_U102; 
assign P3_ADD_552_U166 = ~(P3_ADD_552_U46 & P3_EBX_REG_27__SCAN_IN); 
assign P3_ADD_552_U167 = ~(P3_ADD_552_U102 & P3_EBX_REG_26__SCAN_IN); 
assign P3_ADD_546_U65 = ~(P3_ADD_546_U170 & P3_ADD_546_U169); 
assign P3_ADD_546_U66 = ~(P3_ADD_546_U172 & P3_ADD_546_U171); 
assign P3_ADD_546_U122 = ~P3_ADD_546_U46; 
assign P3_ADD_546_U132 = ~P3_ADD_546_U102; 
assign P3_ADD_546_U166 = ~(P3_ADD_546_U46 & P3_EAX_REG_27__SCAN_IN); 
assign P3_ADD_546_U167 = ~(P3_ADD_546_U102 & P3_EAX_REG_26__SCAN_IN); 
assign P3_ADD_391_1180_U36 = ~(P3_ADD_391_1180_U34 & P3_ADD_391_1180_U26); 
assign P3_ADD_476_U87 = ~(P3_ADD_476_U174 & P3_ADD_476_U173); 
assign P3_ADD_476_U106 = ~P3_ADD_476_U30; 
assign P3_ADD_476_U171 = ~(P3_ADD_476_U30 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_531_U92 = ~(P3_ADD_531_U183 & P3_ADD_531_U182); 
assign P3_ADD_531_U110 = ~P3_ADD_531_U31; 
assign P3_ADD_531_U180 = ~(P3_ADD_531_U31 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_SUB_320_U121 = ~(P3_SUB_320_U94 & P3_SUB_320_U79); 
assign P3_SUB_320_U157 = ~(P3_SUB_320_U94 & P3_SUB_320_U79); 
assign P3_ADD_318_U87 = ~(P3_ADD_318_U174 & P3_ADD_318_U173); 
assign P3_ADD_318_U106 = ~P3_ADD_318_U30; 
assign P3_ADD_318_U171 = ~(P3_ADD_318_U30 & P3_PHYADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_315_U83 = ~(P3_ADD_315_U166 & P3_ADD_315_U165); 
assign P3_ADD_315_U103 = ~P3_ADD_315_U30; 
assign P3_ADD_315_U163 = ~(P3_ADD_315_U30 & P3_PHYADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_360_1242_U88 = ~(P3_ADD_360_1242_U215 & P3_ADD_360_1242_U214); 
assign P3_ADD_360_1242_U109 = P3_ADD_360_1242_U203 & P3_ADD_360_1242_U202; 
assign P3_ADD_360_1242_U120 = ~(P3_ADD_360_1242_U110 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_360_1242_U142 = ~P3_ADD_360_1242_U110; 
assign P3_ADD_360_1242_U143 = ~(P3_ADD_360_U16 & P3_ADD_360_1242_U110); 
assign P3_ADD_360_1242_U206 = ~(P3_ADD_360_1242_U205 & P3_ADD_360_1242_U204); 
assign P3_ADD_467_U87 = ~(P3_ADD_467_U174 & P3_ADD_467_U173); 
assign P3_ADD_467_U106 = ~P3_ADD_467_U30; 
assign P3_ADD_467_U171 = ~(P3_ADD_467_U30 & P3_REIP_REG_15__SCAN_IN); 
assign P3_ADD_430_U87 = ~(P3_ADD_430_U174 & P3_ADD_430_U173); 
assign P3_ADD_430_U106 = ~P3_ADD_430_U30; 
assign P3_ADD_430_U171 = ~(P3_ADD_430_U30 & P3_REIP_REG_15__SCAN_IN); 
assign P3_ADD_380_U92 = ~(P3_ADD_380_U183 & P3_ADD_380_U182); 
assign P3_ADD_380_U110 = ~P3_ADD_380_U31; 
assign P3_ADD_380_U180 = ~(P3_ADD_380_U31 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_344_U92 = ~(P3_ADD_344_U183 & P3_ADD_344_U182); 
assign P3_ADD_344_U110 = ~P3_ADD_344_U31; 
assign P3_ADD_344_U180 = ~(P3_ADD_344_U31 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_339_U87 = ~(P3_ADD_339_U174 & P3_ADD_339_U173); 
assign P3_ADD_339_U106 = ~P3_ADD_339_U30; 
assign P3_ADD_339_U171 = ~(P3_ADD_339_U30 & P3_PHYADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_541_U87 = ~(P3_ADD_541_U174 & P3_ADD_541_U173); 
assign P3_ADD_541_U106 = ~P3_ADD_541_U30; 
assign P3_ADD_541_U171 = ~(P3_ADD_541_U30 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_SUB_357_1258_U117 = ~(P3_SUB_357_1258_U300 & P3_SUB_357_1258_U267); 
assign P3_SUB_357_1258_U326 = ~(P3_SUB_357_1258_U174 & P3_SUB_357_1258_U324); 
assign P3_ADD_515_U87 = ~(P3_ADD_515_U174 & P3_ADD_515_U173); 
assign P3_ADD_515_U106 = ~P3_ADD_515_U30; 
assign P3_ADD_515_U171 = ~(P3_ADD_515_U30 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_394_U87 = ~(P3_ADD_394_U178 & P3_ADD_394_U177); 
assign P3_ADD_394_U109 = ~P3_ADD_394_U30; 
assign P3_ADD_394_U175 = ~(P3_ADD_394_U30 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_SUB_414_U66 = P3_SUB_414_U143 & P3_SUB_414_U142; 
assign P3_SUB_414_U101 = ~P3_SUB_414_U36; 
assign P3_SUB_414_U110 = ~(P3_SUB_414_U109 & P3_EBX_REG_26__SCAN_IN); 
assign P3_SUB_414_U140 = ~(P3_SUB_414_U36 & P3_EBX_REG_27__SCAN_IN); 
assign P3_ADD_441_U87 = ~(P3_ADD_441_U174 & P3_ADD_441_U173); 
assign P3_ADD_441_U106 = ~P3_ADD_441_U30; 
assign P3_ADD_441_U171 = ~(P3_ADD_441_U30 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_349_U92 = ~(P3_ADD_349_U183 & P3_ADD_349_U182); 
assign P3_ADD_349_U110 = ~P3_ADD_349_U31; 
assign P3_ADD_349_U180 = ~(P3_ADD_349_U31 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_405_U87 = ~(P3_ADD_405_U178 & P3_ADD_405_U177); 
assign P3_ADD_405_U109 = ~P3_ADD_405_U30; 
assign P3_ADD_405_U175 = ~(P3_ADD_405_U30 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_553_U92 = ~(P3_ADD_553_U183 & P3_ADD_553_U182); 
assign P3_ADD_553_U110 = ~P3_ADD_553_U31; 
assign P3_ADD_553_U180 = ~(P3_ADD_553_U31 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_558_U92 = ~(P3_ADD_558_U183 & P3_ADD_558_U182); 
assign P3_ADD_558_U110 = ~P3_ADD_558_U31; 
assign P3_ADD_558_U180 = ~(P3_ADD_558_U31 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_385_U92 = ~(P3_ADD_385_U183 & P3_ADD_385_U182); 
assign P3_ADD_385_U110 = ~P3_ADD_385_U31; 
assign P3_ADD_385_U180 = ~(P3_ADD_385_U31 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_547_U92 = ~(P3_ADD_547_U183 & P3_ADD_547_U182); 
assign P3_ADD_547_U110 = ~P3_ADD_547_U31; 
assign P3_ADD_547_U180 = ~(P3_ADD_547_U31 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_371_1212_U112 = P3_ADD_371_1212_U214 & P3_ADD_371_1212_U213; 
assign P3_ADD_371_1212_U113 = ~(P3_ADD_371_1212_U142 & P3_ADD_371_1212_U141); 
assign P3_ADD_371_1212_U217 = ~(P3_ADD_371_1212_U216 & P3_ADD_371_1212_U215); 
assign P3_ADD_371_1212_U226 = ~(P3_ADD_371_1212_U139 & P3_ADD_371_1212_U224); 
assign P3_ADD_494_U87 = ~(P3_ADD_494_U174 & P3_ADD_494_U173); 
assign P3_ADD_494_U106 = ~P3_ADD_494_U30; 
assign P3_ADD_494_U171 = ~(P3_ADD_494_U30 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_536_U87 = ~(P3_ADD_536_U174 & P3_ADD_536_U173); 
assign P3_ADD_536_U106 = ~P3_ADD_536_U30; 
assign P3_ADD_536_U171 = ~(P3_ADD_536_U30 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_402_1132_U36 = ~(P3_ADD_402_1132_U34 & P3_ADD_402_1132_U26); 
assign P2_R2099_U15 = ~(P2_U2743 & P2_R2099_U97); 
assign P2_R2099_U95 = ~(P2_R2099_U167 & P2_R2099_U166); 
assign P2_R2099_U119 = ~P2_R2099_U97; 
assign P2_R2099_U159 = ~(P2_U2743 & P2_R2099_U97); 
assign P2_ADD_391_1196_U20 = ~P2_R2182_U69; 
assign P2_ADD_391_1196_U22 = ~(P2_R2182_U69 & P2_R2096_U68); 
assign P2_ADD_391_1196_U477 = ~(P2_R2182_U69 & P2_ADD_391_1196_U19); 
assign P2_ADD_402_1132_U36 = ~(P2_ADD_402_1132_U34 & P2_ADD_402_1132_U26); 
assign P2_R2182_U67 = ~P2_U2701; 
assign P2_R2182_U101 = ~(P2_R2182_U280 & P2_R2182_U279); 
assign P2_R2182_U188 = ~(P2_U2701 & P2_R2182_U187); 
assign P2_R2182_U231 = ~(P2_U2660 & P2_R2182_U62); 
assign P2_R2182_U233 = ~(P2_U2660 & P2_R2182_U62); 
assign P2_R2167_U28 = ~(P2_U2704 & P2_R2167_U12); 
assign P2_R2167_U34 = ~(P2_U2361 & P2_R2167_U16); 
assign P2_R2027_U92 = ~(P2_R2027_U183 & P2_R2027_U182); 
assign P2_R2027_U110 = ~P2_R2027_U31; 
assign P2_R2027_U180 = ~(P2_R2027_U31 & P2_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P2_R2337_U85 = ~(P2_R2337_U172 & P2_R2337_U171); 
assign P2_R2337_U107 = ~P2_R2337_U31; 
assign P2_R2337_U169 = ~(P2_R2337_U31 & P2_PHYADDRPOINTER_REG_16__SCAN_IN); 
assign P2_R2219_U7 = P2_R2219_U68 & P2_R2219_U66; 
assign P2_R2219_U85 = ~(P2_R2219_U65 & P2_R2219_U84); 
assign P2_R2096_U73 = ~(P2_R2096_U195 & P2_R2096_U194); 
assign P2_R2096_U135 = ~P2_R2096_U103; 
assign P2_R2096_U137 = ~(P2_R2096_U136 & P2_R2096_U103); 
assign P2_R2096_U187 = ~(P2_R2096_U102 & P2_R2096_U103); 
assign P2_GTE_370_U6 = ~(P2_R2219_U25 | P2_GTE_370_U8); 
assign P2_R1957_U121 = ~(P2_R1957_U94 & P2_R1957_U79); 
assign P2_R1957_U157 = ~(P2_R1957_U94 & P2_R1957_U79); 
assign P2_ADD_394_U78 = ~(P2_ADD_394_U158 & P2_ADD_394_U157); 
assign P2_ADD_394_U109 = ~P2_ADD_394_U30; 
assign P2_ADD_394_U151 = ~(P2_ADD_394_U30 & P2_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P2_R2267_U24 = ~(P2_R2267_U89 & P2_R2267_U64 & P2_R2267_U29); 
assign P2_R2267_U28 = ~P2_U3641; 
assign P2_R2267_U65 = P2_R2267_U144 & P2_R2267_U143; 
assign P2_R2267_U101 = ~(P2_U3643 & P2_R2267_U100); 
assign P1_R2027_U65 = ~(P1_R2027_U170 & P1_R2027_U169); 
assign P1_R2027_U66 = ~(P1_R2027_U172 & P1_R2027_U171); 
assign P1_R2027_U122 = ~P1_R2027_U46; 
assign P1_R2027_U132 = ~P1_R2027_U102; 
assign P1_R2027_U166 = ~(P1_R2027_U46 & P1_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P1_R2027_U167 = ~(P1_R2027_U102 & P1_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P1_R2182_U68 = ~(P1_R2182_U57 & P1_R2182_U39); 
assign P1_R2144_U72 = ~P1_U2766; 
assign P1_R2144_U93 = ~(P1_R2144_U129 & P1_R2144_U113); 
assign P1_R2144_U98 = ~(P1_R2144_U113 & P1_R2144_U112); 
assign P1_R2144_U183 = ~(P1_U2766 & P1_R2144_U12); 
assign P1_R2144_U185 = ~(P1_U2355 & P1_R2144_U73); 
assign P1_R2144_U194 = ~(P1_U2766 & P1_R2144_U12); 
assign P1_R2358_U146 = ~P1_U2667; 
assign P1_R2358_U148 = ~P1_U2670; 
assign P1_R2358_U410 = ~(P1_U2667 & P1_R2358_U23); 
assign P1_R2358_U415 = ~(P1_U2667 & P1_R2358_U23); 
assign P1_R2358_U423 = ~(P1_U2670 & P1_R2358_U23); 
assign P1_R2358_U425 = ~(P1_U2352 & P1_R2358_U149); 
assign P1_R2358_U431 = ~(P1_U2352 & P1_R2358_U149); 
assign P1_R2358_U436 = ~(P1_U2670 & P1_R2358_U23); 
assign P1_R2358_U469 = ~(P1_U2352 & P1_R2358_U160); 
assign P1_R2358_U485 = ~(P1_U2352 & P1_R2358_U160); 
assign P1_R2099_U37 = ~(P1_R2099_U215 & P1_R2099_U214); 
assign P1_R2099_U38 = ~(P1_R2099_U217 & P1_R2099_U216); 
assign P1_R2099_U160 = ~P1_R2099_U109; 
assign P1_R2099_U161 = ~P1_R2099_U10; 
assign P1_R2099_U213 = ~(P1_R2099_U26 & P1_R2099_U109); 
assign P1_R2099_U344 = ~(P1_R2099_U62 & P1_R2099_U10); 
assign P1_R2337_U87 = ~(P1_R2337_U174 & P1_R2337_U173); 
assign P1_R2337_U106 = ~P1_R2337_U30; 
assign P1_R2337_U171 = ~(P1_R2337_U30 & P1_PHYADDRPOINTER_REG_15__SCAN_IN); 
assign P1_R2096_U87 = ~(P1_R2096_U174 & P1_R2096_U173); 
assign P1_R2096_U106 = ~P1_R2096_U30; 
assign P1_R2096_U171 = ~(P1_R2096_U30 & P1_REIP_REG_15__SCAN_IN); 
assign P1_ADD_405_U78 = ~(P1_ADD_405_U158 & P1_ADD_405_U157); 
assign P1_ADD_405_U109 = ~P1_ADD_405_U30; 
assign P1_ADD_405_U151 = ~(P1_ADD_405_U30 & P1_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P1_ADD_515_U78 = ~(P1_ADD_515_U156 & P1_ADD_515_U155); 
assign P1_ADD_515_U106 = ~P1_ADD_515_U30; 
assign P1_ADD_515_U149 = ~(P1_ADD_515_U30 & P1_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_U2826 = ~(P3_U6438 & P3_U6437 & P3_U6439 & P3_U6440 & P3_U3958); 
assign P3_U2859 = ~(P3_U5727 & P3_U5725 & P3_U5726); 
assign P3_U2860 = ~(P3_U5703 & P3_U5701 & P3_U5702); 
assign P3_U2861 = ~(P3_U5679 & P3_U5677 & P3_U5678); 
assign P3_U2862 = ~(P3_U5654 & P3_U5653 & P3_U5655); 
assign P3_U3305 = ~(P3_U8047 & P3_U8046); 
assign P3_U3306 = ~(P3_U8049 & P3_U8048); 
assign P3_U3307 = ~(P3_U8051 & P3_U8050); 
assign P3_U3308 = ~(P3_U8053 & P3_U8052); 
assign P3_U3737 = P3_U3736 & P3_U3735 & P3_U5771; 
assign P3_U3959 = P3_U6450 & P3_U6449 & P3_U6452 & P3_U6451; 
assign P3_U4031 = P3_U7098 & P3_U7097 & P3_U4032; 
assign P3_U4035 = P3_U7108 & P3_U7107 & P3_U4036; 
assign P3_U4039 = P3_U7118 & P3_U7117 & P3_U4040; 
assign P3_U4043 = P3_U7128 & P3_U7127 & P3_U4044; 
assign P3_U4047 = P3_U7137 & P3_U4316 & P3_U7138; 
assign P3_U4052 = P3_U7147 & P3_U4316 & P3_U7148; 
assign P3_U4057 = P3_U7157 & P3_U4316 & P3_U7158; 
assign P3_U4060 = P3_U7165 & P3_U4316 & P3_U7166; 
assign P3_U4063 = P3_U7173 & P3_U4316 & P3_U7174; 
assign P3_U4066 = P3_U7181 & P3_U4316 & P3_U7182; 
assign P3_U4069 = P3_U7189 & P3_U4316 & P3_U7190; 
assign P3_U4072 = P3_U7197 & P3_U4316 & P3_U7198; 
assign P3_U4075 = P3_U7205 & P3_U4316 & P3_U7206; 
assign P3_U4078 = P3_U7213 & P3_U4316 & P3_U7214; 
assign P3_U5546 = ~(P3_U5545 & P3_U5544); 
assign P3_U5557 = ~(P3_U3680 & P3_U5556); 
assign P3_U5570 = ~(P3_U3683 & P3_U5569); 
assign P3_U5577 = ~(P3_U3684 & P3_U5575); 
assign P3_U5748 = ~(P3_U5730 & P3_U3726 & P3_U5728 & P3_U3722 & P3_U3729); 
assign P3_U5776 = ~(P3_ADD_360_1242_U88 & P3_U2395); 
assign P3_U5946 = ~(P3_ADD_558_U92 & P3_U3220); 
assign P3_U5947 = ~(P3_ADD_553_U92 & P3_U4298); 
assign P3_U5948 = ~(P3_ADD_547_U92 & P3_U4299); 
assign P3_U5951 = ~(P3_ADD_531_U92 & P3_U2354); 
assign P3_U5959 = ~(P3_ADD_385_U92 & P3_U2358); 
assign P3_U5960 = ~(P3_ADD_380_U92 & P3_U2359); 
assign P3_U5961 = ~(P3_ADD_349_U92 & P3_U4306); 
assign P3_U5962 = ~(P3_ADD_344_U92 & P3_U2362); 
assign P3_U5973 = ~(P3_ADD_541_U87 & P3_U4300); 
assign P3_U5974 = ~(P3_ADD_536_U87 & P3_U4301); 
assign P3_U5977 = ~(P3_ADD_515_U87 & P3_U4302); 
assign P3_U5978 = ~(P3_ADD_494_U87 & P3_U2356); 
assign P3_U5979 = ~(P3_ADD_476_U87 & P3_U4303); 
assign P3_U5980 = ~(P3_ADD_441_U87 & P3_U4304); 
assign P3_U5981 = ~(P3_ADD_405_U87 & P3_U4305); 
assign P3_U5982 = ~(P3_ADD_394_U87 & P3_U2357); 
assign P3_U6216 = ~(P3_ADD_526_U66 & P3_U2355); 
assign P3_U6240 = ~(P3_ADD_526_U65 & P3_U2355); 
assign P3_U6455 = ~(P3_U2396 & P3_ADD_360_1242_U88); 
assign P3_U6517 = ~(P3_ADD_318_U87 & P3_U2398); 
assign P3_U6522 = ~(P3_ADD_339_U87 & P3_U2388); 
assign P3_U6526 = ~(P3_ADD_315_U83 & P3_U2397); 
assign P3_U6961 = ~(P3_ADD_546_U66 & P3_U2400); 
assign P3_U6966 = ~(P3_ADD_546_U65 & P3_U2400); 
assign P3_U7071 = ~(P3_ADD_552_U66 & P3_U2399); 
assign P3_U7074 = ~(P3_ADD_552_U65 & P3_U2399); 
assign P3_U7099 = ~(P3_U7910 & P3_EBX_REG_0__SCAN_IN); 
assign P3_U7109 = ~(P3_U7910 & P3_EBX_REG_1__SCAN_IN); 
assign P3_U7119 = ~(P3_U7910 & P3_EBX_REG_2__SCAN_IN); 
assign P3_U7129 = ~(P3_U7910 & P3_EBX_REG_3__SCAN_IN); 
assign P3_U7139 = ~(P3_U7910 & P3_EBX_REG_4__SCAN_IN); 
assign P3_U7149 = ~(P3_U7910 & P3_EBX_REG_5__SCAN_IN); 
assign P3_U7159 = ~(P3_U7910 & P3_EBX_REG_6__SCAN_IN); 
assign P3_U7167 = ~(P3_U7910 & P3_EBX_REG_7__SCAN_IN); 
assign P3_U7175 = ~(P3_U7910 & P3_EBX_REG_8__SCAN_IN); 
assign P3_U7183 = ~(P3_U7910 & P3_EBX_REG_9__SCAN_IN); 
assign P3_U7191 = ~(P3_U7910 & P3_EBX_REG_10__SCAN_IN); 
assign P3_U7199 = ~(P3_U7910 & P3_EBX_REG_11__SCAN_IN); 
assign P3_U7207 = ~(P3_U7910 & P3_EBX_REG_12__SCAN_IN); 
assign P3_U7215 = ~(P3_U7910 & P3_EBX_REG_13__SCAN_IN); 
assign P3_U7222 = ~(P3_ADD_467_U87 & P3_U2601); 
assign P3_U7223 = ~(P3_U7910 & P3_EBX_REG_14__SCAN_IN); 
assign P3_U7224 = ~(P3_ADD_430_U87 & P3_U2405); 
assign P3_U7231 = ~(P3_U7910 & P3_EBX_REG_15__SCAN_IN); 
assign P3_U7239 = ~(P3_U7910 & P3_EBX_REG_16__SCAN_IN); 
assign P3_U7247 = ~(P3_U7910 & P3_EBX_REG_17__SCAN_IN); 
assign P3_U7255 = ~(P3_U7910 & P3_EBX_REG_18__SCAN_IN); 
assign P3_U7263 = ~(P3_U7910 & P3_EBX_REG_19__SCAN_IN); 
assign P3_U7271 = ~(P3_U7910 & P3_EBX_REG_20__SCAN_IN); 
assign P3_U7279 = ~(P3_U7910 & P3_EBX_REG_21__SCAN_IN); 
assign P3_U7287 = ~(P3_U7910 & P3_EBX_REG_22__SCAN_IN); 
assign P3_U7295 = ~(P3_U7910 & P3_EBX_REG_23__SCAN_IN); 
assign P3_U7303 = ~(P3_U7910 & P3_EBX_REG_24__SCAN_IN); 
assign P3_U7309 = ~(P3_SUB_414_U66 & P3_U2602); 
assign P3_U7311 = ~(P3_U7910 & P3_EBX_REG_25__SCAN_IN); 
assign P3_U7319 = ~(P3_U7910 & P3_EBX_REG_26__SCAN_IN); 
assign P3_U7327 = ~(P3_U7910 & P3_EBX_REG_27__SCAN_IN); 
assign P3_U7335 = ~(P3_U7910 & P3_EBX_REG_28__SCAN_IN); 
assign P3_U7343 = ~(P3_U7910 & P3_EBX_REG_29__SCAN_IN); 
assign P3_U7351 = ~(P3_U7910 & P3_EBX_REG_30__SCAN_IN); 
assign P3_U7360 = ~(P3_U7910 & P3_EBX_REG_31__SCAN_IN); 
assign P3_U7906 = ~(P3_U3939 & P3_U6397); 
assign P2_U2466 = P2_R2099_U96 & P2_R2099_U95; 
assign P2_U2483 = P2_R2099_U95 & P2_U3322; 
assign P2_U2504 = ~(P2_R2099_U95 | P2_R2099_U96); 
assign P2_U3287 = ~P2_GTE_370_U6; 
assign P2_U3321 = ~P2_R2099_U95; 
assign P2_U3640 = ~(P2_U8334 & P2_U8333); 
assign P2_U4447 = ~(P2_R2219_U7 & P2_U2617); 
assign P2_U4612 = ~(P2_GTE_370_U6 & P2_U4417); 
assign P2_U5610 = ~(P2_R2099_U95 & P2_U5603); 
assign P2_U5622 = ~(P2_U4466 & P2_U5619); 
assign P2_U5666 = ~(P2_GTE_370_U6 & P2_U4417); 
assign P2_U7138 = ~(P2_U4467 & P2_R2099_U95); 
assign P2_U8326 = ~(P2_U3242 & P2_R2267_U65); 
assign P2_U8407 = ~(P2_R2337_U85 & P2_U3284); 
assign P1_U2381 = P1_U2357 & P1_U3271; 
assign P1_U2382 = P1_U2357 & P1_U4477; 
assign P1_U2425 = P1_U2368 & P1_U2448; 
assign P1_U3321 = ~(P1_U3306 & P1_U4535); 
assign P1_U3328 = ~(P1_U3324 & P1_U4603); 
assign P1_U3335 = ~(P1_U3330 & P1_U4661); 
assign P1_U3339 = ~(P1_U3337 & P1_U4719); 
assign P1_U3344 = ~(P1_U3341 & P1_U4776); 
assign P1_U3348 = ~(P1_U3346 & P1_U4834); 
assign P1_U3351 = ~(P1_U3349 & P1_U4891); 
assign P1_U3355 = ~(P1_U3353 & P1_U4949); 
assign P1_U3375 = ~(P1_U3373 & P1_U5234); 
assign P1_U3379 = ~(P1_U3377 & P1_U5292); 
assign P1_U3382 = ~(P1_U3380 & P1_U5349); 
assign P1_U3386 = ~(P1_U3384 & P1_U5407); 
assign P1_U3406 = ~(P1_U3271 & P1_U3273); 
assign P1_U3883 = P1_U6151 & P1_U6150; 
assign P1_U4248 = ~(P1_U2451 & P1_U2353 & P1_U3862 & P1_U2448); 
assign P1_U4252 = ~P1_U3299; 
assign P1_U4259 = ~P1_U3281; 
assign P1_U4509 = ~(P1_U2448 & P1_U4262); 
assign P1_U4547 = ~(P1_U4546 & P1_U3297 & P1_U3299); 
assign P1_U5005 = ~(P1_U2439 & P1_U2442); 
assign P1_U5062 = ~(P1_U2439 & P1_U2443); 
assign P1_U5119 = ~(P1_U2439 & P1_U2444); 
assign P1_U5177 = ~(P1_U2439 & P1_U2445); 
assign P1_U5508 = ~(P1_U2427 & P1_U5506); 
assign P1_U6263 = ~(P1_U4198 & P1_U3273); 
assign P1_U6846 = ~(P1_R2337_U87 & P1_U2352); 
assign P1_U7503 = ~(P1_U7502 & P1_U6149); 
assign P1_U7541 = ~(P1_U2357 & P1_U7493); 
assign P1_U7543 = ~(P1_U2357 & P1_U7493); 
assign P1_U7545 = ~(P1_U2357 & P1_U7493); 
assign P1_U7547 = ~(P1_U2357 & P1_U7493); 
assign P1_U7549 = ~(P1_U2357 & P1_U7493); 
assign P1_U7551 = ~(P1_U2357 & P1_U7493); 
assign P1_U7553 = ~(P1_U2357 & P1_U7493); 
assign P1_U7555 = ~(P1_U2357 & P1_U7493); 
assign P1_U7557 = ~(P1_U2357 & P1_U7493); 
assign P1_U7559 = ~(P1_U2357 & P1_U7493); 
assign P1_U7561 = ~(P1_U2357 & P1_U7493); 
assign P1_U7563 = ~(P1_U2357 & P1_U7493); 
assign P1_U7565 = ~(P1_U2357 & P1_U7493); 
assign P1_U7567 = ~(P1_U2357 & P1_U7493); 
assign P1_U7569 = ~(P1_U2357 & P1_U7493); 
assign P1_U7571 = ~(P1_U2357 & P1_U7493); 
assign P1_U7573 = ~(P1_U2357 & P1_U7493); 
assign P1_U7575 = ~(P1_U2357 & P1_U7493); 
assign P1_U7577 = ~(P1_U2357 & P1_U7493); 
assign P1_U7579 = ~(P1_U2357 & P1_U7493); 
assign P1_U7581 = ~(P1_U2357 & P1_U7493); 
assign P1_U7583 = ~(P1_U2357 & P1_U7493); 
assign P1_U7585 = ~(P1_U2357 & P1_U7493); 
assign P1_U7587 = ~(P1_U2357 & P1_U7493); 
assign P1_U7589 = ~(P1_U2357 & P1_U7493); 
assign P1_U7591 = ~(P1_U2357 & P1_U7493); 
assign P1_U7593 = ~(P1_U2357 & P1_U7493); 
assign P1_U7595 = ~(P1_U2357 & P1_U7493); 
assign P1_U7597 = ~(P1_U2357 & P1_U7493); 
assign P1_U7599 = ~(P1_U2357 & P1_U7493); 
assign P1_U7601 = ~(P1_U2357 & P1_U7493); 
assign P1_U7680 = ~(P1_U7501 & P1_U3284); 
assign P1_U7682 = ~(P1_U4506 & P1_U3273); 
assign P1_U7697 = ~(P1_U4216 & P1_U3273); 
assign P1_U7741 = ~(P1_U3271 & P1_U3281); 
assign P3_ADD_526_U48 = ~(P3_ADD_526_U94 & P3_ADD_526_U122); 
assign P3_ADD_526_U101 = ~(P3_ADD_526_U122 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_526_U165 = ~(P3_ADD_526_U122 & P3_ADD_526_U44); 
assign P3_ADD_526_U168 = ~(P3_ADD_526_U132 & P3_ADD_526_U41); 
assign P3_ADD_552_U48 = ~(P3_ADD_552_U94 & P3_ADD_552_U122); 
assign P3_ADD_552_U101 = ~(P3_ADD_552_U122 & P3_EBX_REG_27__SCAN_IN); 
assign P3_ADD_552_U165 = ~(P3_ADD_552_U122 & P3_ADD_552_U44); 
assign P3_ADD_552_U168 = ~(P3_ADD_552_U132 & P3_ADD_552_U41); 
assign P3_ADD_546_U48 = ~(P3_ADD_546_U94 & P3_ADD_546_U122); 
assign P3_ADD_546_U101 = ~(P3_ADD_546_U122 & P3_EAX_REG_27__SCAN_IN); 
assign P3_ADD_546_U165 = ~(P3_ADD_546_U122 & P3_ADD_546_U44); 
assign P3_ADD_546_U168 = ~(P3_ADD_546_U132 & P3_ADD_546_U41); 
assign P3_ADD_391_1180_U18 = ~(P3_ADD_391_1180_U36 & P3_ADD_391_1180_U35); 
assign P3_ADD_476_U32 = ~(P3_ADD_476_U106 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_476_U172 = ~(P3_ADD_476_U106 & P3_ADD_476_U31); 
assign P3_ADD_531_U33 = ~(P3_ADD_531_U110 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_531_U181 = ~(P3_ADD_531_U110 & P3_ADD_531_U32); 
assign P3_SUB_320_U47 = ~P3_ADD_318_U87; 
assign P3_SUB_320_U80 = P3_SUB_320_U157 & P3_SUB_320_U156; 
assign P3_SUB_320_U122 = ~(P3_ADD_318_U87 & P3_SUB_320_U121); 
assign P3_ADD_318_U32 = ~(P3_ADD_318_U106 & P3_PHYADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_318_U172 = ~(P3_ADD_318_U106 & P3_ADD_318_U31); 
assign P3_ADD_315_U32 = ~(P3_ADD_315_U103 & P3_PHYADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_315_U164 = ~(P3_ADD_315_U103 & P3_ADD_315_U31); 
assign P3_ADD_360_1242_U108 = ~(P3_ADD_360_1242_U143 & P3_ADD_360_1242_U120 & P3_ADD_360_1242_U189); 
assign P3_ADD_360_1242_U207 = ~(P3_ADD_360_1242_U109 & P3_ADD_360_1242_U110); 
assign P3_ADD_360_1242_U208 = ~(P3_ADD_360_1242_U142 & P3_ADD_360_1242_U206); 
assign P3_ADD_467_U32 = ~(P3_ADD_467_U106 & P3_REIP_REG_15__SCAN_IN); 
assign P3_ADD_467_U172 = ~(P3_ADD_467_U106 & P3_ADD_467_U31); 
assign P3_ADD_430_U32 = ~(P3_ADD_430_U106 & P3_REIP_REG_15__SCAN_IN); 
assign P3_ADD_430_U172 = ~(P3_ADD_430_U106 & P3_ADD_430_U31); 
assign P3_ADD_380_U33 = ~(P3_ADD_380_U110 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_380_U181 = ~(P3_ADD_380_U110 & P3_ADD_380_U32); 
assign P3_ADD_344_U33 = ~(P3_ADD_344_U110 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_344_U181 = ~(P3_ADD_344_U110 & P3_ADD_344_U32); 
assign P3_ADD_339_U32 = ~(P3_ADD_339_U106 & P3_PHYADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_339_U172 = ~(P3_ADD_339_U106 & P3_ADD_339_U31); 
assign P3_ADD_541_U32 = ~(P3_ADD_541_U106 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_541_U172 = ~(P3_ADD_541_U106 & P3_ADD_541_U31); 
assign P3_SUB_357_1258_U72 = ~(P3_SUB_357_1258_U326 & P3_SUB_357_1258_U325); 
assign P3_SUB_357_1258_U152 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U117); 
assign P3_SUB_357_1258_U176 = ~(P3_SUB_357_1258_U117 & P3_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P3_SUB_357_1258_U301 = ~P3_SUB_357_1258_U117; 
assign P3_SUB_357_1258_U318 = ~(P3_SUB_357_1258_U116 & P3_SUB_357_1258_U117); 
assign P3_ADD_515_U32 = ~(P3_ADD_515_U106 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_515_U172 = ~(P3_ADD_515_U106 & P3_ADD_515_U31); 
assign P3_ADD_394_U32 = ~(P3_ADD_394_U109 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_394_U176 = ~(P3_ADD_394_U109 & P3_ADD_394_U31); 
assign P3_SUB_414_U14 = P3_SUB_414_U110 & P3_SUB_414_U36; 
assign P3_SUB_414_U37 = ~(P3_SUB_414_U40 & P3_SUB_414_U63 & P3_SUB_414_U101); 
assign P3_SUB_414_U107 = ~(P3_SUB_414_U101 & P3_SUB_414_U63); 
assign P3_SUB_414_U141 = ~(P3_SUB_414_U101 & P3_SUB_414_U63); 
assign P3_ADD_441_U32 = ~(P3_ADD_441_U106 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_441_U172 = ~(P3_ADD_441_U106 & P3_ADD_441_U31); 
assign P3_ADD_349_U33 = ~(P3_ADD_349_U110 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_349_U181 = ~(P3_ADD_349_U110 & P3_ADD_349_U32); 
assign P3_ADD_405_U32 = ~(P3_ADD_405_U109 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_405_U176 = ~(P3_ADD_405_U109 & P3_ADD_405_U31); 
assign P3_ADD_553_U33 = ~(P3_ADD_553_U110 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_553_U181 = ~(P3_ADD_553_U110 & P3_ADD_553_U32); 
assign P3_ADD_558_U33 = ~(P3_ADD_558_U110 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_558_U181 = ~(P3_ADD_558_U110 & P3_ADD_558_U32); 
assign P3_ADD_385_U33 = ~(P3_ADD_385_U110 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_385_U181 = ~(P3_ADD_385_U110 & P3_ADD_385_U32); 
assign P3_ADD_547_U33 = ~(P3_ADD_547_U110 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_547_U181 = ~(P3_ADD_547_U110 & P3_ADD_547_U32); 
assign P3_ADD_371_1212_U90 = ~(P3_ADD_371_1212_U226 & P3_ADD_371_1212_U225); 
assign P3_ADD_371_1212_U118 = ~(P3_ADD_371_1212_U113 & P3_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P3_ADD_371_1212_U143 = ~P3_ADD_371_1212_U113; 
assign P3_ADD_371_1212_U144 = ~(P3_ADD_371_U17 & P3_ADD_371_1212_U113); 
assign P3_ADD_371_1212_U218 = ~(P3_ADD_371_1212_U112 & P3_ADD_371_1212_U113); 
assign P3_ADD_494_U32 = ~(P3_ADD_494_U106 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_494_U172 = ~(P3_ADD_494_U106 & P3_ADD_494_U31); 
assign P3_ADD_536_U32 = ~(P3_ADD_536_U106 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_536_U172 = ~(P3_ADD_536_U106 & P3_ADD_536_U31); 
assign P3_ADD_402_1132_U18 = ~(P3_ADD_402_1132_U36 & P3_ADD_402_1132_U35); 
assign P2_R2099_U120 = ~P2_R2099_U15; 
assign P2_R2099_U157 = ~(P2_U2742 & P2_R2099_U15); 
assign P2_R2099_U160 = ~(P2_R2099_U119 & P2_R2099_U14); 
assign P2_ADD_391_1196_U18 = ~P2_R2096_U73; 
assign P2_ADD_391_1196_U162 = ~P2_ADD_391_1196_U22; 
assign P2_ADD_391_1196_U163 = ~(P2_ADD_391_1196_U23 & P2_ADD_391_1196_U22); 
assign P2_ADD_391_1196_U478 = ~(P2_R2096_U68 & P2_ADD_391_1196_U20); 
assign P2_ADD_402_1132_U18 = ~(P2_ADD_402_1132_U36 & P2_ADD_402_1132_U35); 
assign P2_R2182_U42 = ~P2_U2700; 
assign P2_R2182_U64 = ~P2_U2683; 
assign P2_R2182_U110 = P2_R2182_U232 & P2_R2182_U231; 
assign P2_R2182_U123 = ~(P2_R2182_U122 & P2_R2182_U67); 
assign P2_R2182_U124 = P2_U2679 | P2_U2700; 
assign P2_R2182_U127 = ~(P2_U2679 & P2_U2700); 
assign P2_R2182_U179 = P2_U2683 | P2_U2659; 
assign P2_R2182_U181 = ~(P2_U2659 & P2_U2683); 
assign P2_R2182_U183 = ~(P2_U2659 & P2_U2683); 
assign P2_R2182_U185 = P2_U2659 | P2_U2683; 
assign P2_R2182_U191 = ~(P2_U2679 & P2_U2700); 
assign P2_R2182_U223 = ~(P2_U2700 & P2_R2182_U43); 
assign P2_R2182_U225 = ~(P2_U2683 & P2_R2182_U65); 
assign P2_R2182_U227 = ~(P2_U2683 & P2_R2182_U65); 
assign P2_R2182_U235 = ~(P2_R2182_U234 & P2_R2182_U233); 
assign P2_R2182_U281 = ~P2_R2182_U101; 
assign P2_R2182_U283 = ~(P2_R2182_U101 & P2_R2182_U67); 
assign P2_R2167_U18 = ~P2_U2708; 
assign P2_R2167_U29 = ~(P2_R2167_U27 & P2_R2167_U28 & P2_R2167_U26); 
assign P2_R2167_U40 = ~(P2_U2708 & P2_R2167_U15); 
assign P2_R2167_U42 = ~(P2_R2167_U17 & P2_R2167_U15 & P2_U2708); 
assign P2_R2027_U33 = ~(P2_R2027_U110 & P2_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P2_R2027_U181 = ~(P2_R2027_U110 & P2_R2027_U32); 
assign P2_R2337_U33 = ~(P2_R2337_U107 & P2_PHYADDRPOINTER_REG_16__SCAN_IN); 
assign P2_R2337_U170 = ~(P2_R2337_U107 & P2_R2337_U32); 
assign P2_R2219_U24 = ~(P2_R2219_U86 & P2_R2219_U85); 
assign P2_R2096_U101 = ~(P2_R2096_U138 & P2_R2096_U137); 
assign P2_R2096_U188 = ~(P2_R2096_U135 & P2_R2096_U186); 
assign P2_R1957_U46 = ~P2_U3677; 
assign P2_R1957_U80 = P2_R1957_U157 & P2_R1957_U156; 
assign P2_R1957_U122 = ~(P2_U3677 & P2_R1957_U121); 
assign P2_ADD_394_U32 = ~(P2_ADD_394_U109 & P2_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P2_ADD_394_U152 = ~(P2_ADD_394_U109 & P2_ADD_394_U31); 
assign P2_R2267_U17 = P2_R2267_U101 & P2_R2267_U24; 
assign P2_R2267_U90 = ~P2_R2267_U24; 
assign P2_R2267_U139 = ~(P2_U3642 & P2_R2267_U24); 
assign P1_R2027_U48 = ~(P1_R2027_U94 & P1_R2027_U122); 
assign P1_R2027_U101 = ~(P1_R2027_U122 & P1_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P1_R2027_U165 = ~(P1_R2027_U122 & P1_R2027_U44); 
assign P1_R2027_U168 = ~(P1_R2027_U132 & P1_R2027_U41); 
assign P1_R2182_U26 = ~(P1_R2182_U68 & P1_R2182_U67); 
assign P1_R2144_U28 = ~(P1_R2144_U186 & P1_R2144_U185); 
assign P1_R2144_U75 = ~P1_U2765; 
assign P1_R2144_U130 = ~P1_R2144_U93; 
assign P1_R2144_U148 = ~P1_R2144_U98; 
assign P1_R2144_U182 = ~(P1_U2355 & P1_R2144_U72); 
assign P1_R2144_U193 = ~(P1_U2355 & P1_R2144_U72); 
assign P1_R2144_U196 = ~(P1_U2765 & P1_R2144_U12); 
assign P1_R2144_U198 = ~(P1_U2765 & P1_R2144_U12); 
assign P1_R2144_U259 = ~(P1_U2355 & P1_R2144_U98); 
assign P1_R2358_U147 = ~P1_U2668; 
assign P1_R2358_U151 = ~P1_U2669; 
assign P1_R2358_U159 = ~P1_U2613; 
assign P1_R2358_U409 = ~(P1_U2352 & P1_R2358_U146); 
assign P1_R2358_U412 = ~(P1_U2668 & P1_R2358_U23); 
assign P1_R2358_U414 = ~(P1_U2352 & P1_R2358_U146); 
assign P1_R2358_U422 = ~(P1_U2352 & P1_R2358_U148); 
assign P1_R2358_U427 = ~(P1_R2358_U426 & P1_R2358_U425); 
assign P1_R2358_U435 = ~(P1_U2352 & P1_R2358_U148); 
assign P1_R2358_U438 = ~(P1_U2669 & P1_R2358_U23); 
assign P1_R2358_U440 = ~(P1_U2669 & P1_R2358_U23); 
assign P1_R2358_U443 = ~(P1_U2668 & P1_R2358_U23); 
assign P1_R2358_U462 = ~(P1_U2613 & P1_R2358_U23); 
assign P1_R2358_U468 = ~(P1_U2613 & P1_R2358_U23); 
assign P1_R2358_U471 = ~(P1_R2358_U470 & P1_R2358_U469); 
assign P1_R2099_U11 = ~(P1_R2099_U92 & P1_R2099_U161); 
assign P1_R2099_U144 = ~(P1_R2099_U161 & P1_R2099_U62); 
assign P1_R2099_U212 = ~(P1_R2099_U160 & P1_R2099_U211); 
assign P1_R2099_U343 = ~(P1_R2099_U261 & P1_R2099_U161); 
assign P1_R2337_U32 = ~(P1_R2337_U106 & P1_PHYADDRPOINTER_REG_15__SCAN_IN); 
assign P1_R2337_U172 = ~(P1_R2337_U106 & P1_R2337_U31); 
assign P1_R2096_U32 = ~(P1_R2096_U106 & P1_REIP_REG_15__SCAN_IN); 
assign P1_R2096_U172 = ~(P1_R2096_U106 & P1_R2096_U31); 
assign P1_ADD_405_U32 = ~(P1_ADD_405_U109 & P1_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P1_ADD_405_U152 = ~(P1_ADD_405_U109 & P1_ADD_405_U31); 
assign P1_ADD_515_U32 = ~(P1_ADD_515_U106 & P1_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P1_ADD_515_U150 = ~(P1_ADD_515_U106 & P1_ADD_515_U31); 
assign P3_U2678 = ~(P3_U7075 & P3_U7073 & P3_U7074); 
assign P3_U2679 = ~(P3_U7072 & P3_U7070 & P3_U7071); 
assign P3_U2710 = ~(P3_U6964 & P3_U6963 & P3_U4027 & P3_U6966); 
assign P3_U2711 = ~(P3_U6959 & P3_U6958 & P3_U4026 & P3_U6961); 
assign P3_U2825 = ~(P3_U6446 & P3_U6445 & P3_U6448 & P3_U6447 & P3_U3959); 
assign P3_U3738 = P3_U3739 & P3_U5776; 
assign P3_U3790 = P3_U5948 & P3_U5947; 
assign P3_U3792 = P3_U5950 & P3_U5949 & P3_U5951 & P3_U3791; 
assign P3_U3794 = P3_U5962 & P3_U5961 & P3_U5960 & P3_U5959; 
assign P3_U3797 = P3_U5977 & P3_U5976; 
assign P3_U3800 = P3_U5979 & P3_U5978 & P3_U5980 & P3_U5982 & P3_U5981; 
assign P3_U4081 = P3_U7221 & P3_U4316 & P3_U7222; 
assign P3_U5750 = ~(P3_U4318 & P3_U5748); 
assign P3_U5772 = ~(P3_U3734 & P3_U5754 & P3_U5753 & P3_U3730 & P3_U3737); 
assign P3_U5795 = ~(P3_ADD_371_1212_U90 & P3_U2360); 
assign P3_U5801 = ~(P3_SUB_357_1258_U72 & P3_U2393); 
assign P3_U6459 = ~(P3_U2387 & P3_ADD_371_1212_U90); 
assign P3_U6464 = ~(P3_U2394 & P3_SUB_357_1258_U72); 
assign P3_U6990 = ~(P3_ADD_391_1180_U18 & P3_U2411); 
assign P3_U7088 = ~(P3_ADD_402_1132_U18 & P3_U2408); 
assign P3_U7317 = ~(P3_SUB_414_U14 & P3_U2602); 
assign P3_U7980 = ~(P3_U5546 & P3_U4283); 
assign P3_U7990 = ~(P3_U5557 & P3_U4283); 
assign P3_U7992 = ~(P3_U5570 & P3_U4283); 
assign P3_U7996 = ~(P3_U5577 & P3_U4283); 
assign P2_U2492 = P2_R2099_U96 & P2_U3321; 
assign P2_U2682 = P2_U2355 & P2_ADD_402_1132_U18; 
assign P2_U2699 = ~(P2_U7139 & P2_U7140 & P2_U7138); 
assign P2_U2766 = ~(P2_U4447 & P2_U7539); 
assign P2_U2767 = ~(P2_U4447 & P2_U7540); 
assign P2_U2768 = ~(P2_U4447 & P2_U7541); 
assign P2_U2769 = ~(P2_U4447 & P2_U7542); 
assign P2_U2770 = ~(P2_U4447 & P2_U7543); 
assign P2_U2771 = ~(P2_U4447 & P2_U7544); 
assign P2_U2772 = ~(P2_U4447 & P2_U7545); 
assign P2_U2773 = ~(P2_U4447 & P2_U7546); 
assign P2_U2774 = ~(P2_U4447 & P2_U7547); 
assign P2_U2775 = ~(P2_U4447 & P2_U7548); 
assign P2_U2776 = ~(P2_U4447 & P2_U7549); 
assign P2_U2777 = ~(P2_U4447 & P2_U7550); 
assign P2_U2778 = ~(P2_U4447 & P2_U7551); 
assign P2_U2779 = ~(P2_U4447 & P2_U7552); 
assign P2_U2780 = ~(P2_U4447 & P2_U7553); 
assign P2_U2781 = ~(P2_U4447 & P2_U7554); 
assign P2_U2782 = ~(P2_U4447 & P2_U7555); 
assign P2_U2783 = ~(P2_U4447 & P2_U7556); 
assign P2_U2784 = ~(P2_U4447 & P2_U7557); 
assign P2_U2785 = ~(P2_U4447 & P2_U7558); 
assign P2_U2786 = ~(P2_U4447 & P2_U7559); 
assign P2_U2787 = ~(P2_U4447 & P2_U7560); 
assign P2_U2788 = ~(P2_U4447 & P2_U7537); 
assign P2_U2789 = ~(P2_U4447 & P2_U7538); 
assign P2_U3555 = ~(P2_U2504 & P2_U2479); 
assign P2_U3556 = ~(P2_U2504 & P2_U2473); 
assign P2_U3557 = ~(P2_U2504 & P2_U2470); 
assign P2_U3558 = ~(P2_U2504 & P2_U2467); 
assign P2_U3563 = ~(P2_U2483 & P2_U2479); 
assign P2_U3564 = ~(P2_U2483 & P2_U2473); 
assign P2_U3565 = ~(P2_U2483 & P2_U2470); 
assign P2_U3566 = ~(P2_U2483 & P2_U2467); 
assign P2_U3567 = ~(P2_U2479 & P2_U2466); 
assign P2_U3568 = ~(P2_U2473 & P2_U2466); 
assign P2_U3569 = ~(P2_U2470 & P2_U2466); 
assign P2_U3570 = ~(P2_U2466 & P2_U2467); 
assign P2_U3676 = ~(P2_U8408 & P2_U8407); 
assign P2_U4606 = ~(P2_U4417 & P2_U3287); 
assign P2_U5611 = ~(P2_U3884 & P2_U5610); 
assign P2_U8131 = ~(P2_U3287 & P2_U7873); 
assign P2_U8324 = ~(P2_U3242 & P2_R2267_U17); 
assign P2_U8331 = ~(P2_R2219_U24 & P2_U2617); 
assign P1_U2473 = P1_U7680 & P1_U7679 & P1_U3406; 
assign P1_U2612 = ~(P1_U6844 & P1_U6845 & P1_U6846); 
assign P1_U3300 = ~(P1_U4547 & P1_U3294); 
assign P1_U3361 = ~(P1_U3356 & P1_U5005); 
assign P1_U3365 = ~(P1_U3363 & P1_U5062); 
assign P1_U3368 = ~(P1_U3366 & P1_U5119); 
assign P1_U3372 = ~(P1_U3370 & P1_U5177); 
assign P1_U3416 = ~(P1_U3863 & P1_U4248); 
assign P1_U4182 = ~(P1_U7698 & P1_U7697 & P1_U3738); 
assign P1_U4260 = ~P1_U3406; 
assign P1_U4508 = ~(P1_U7682 & P1_U7681 & P1_U4507); 
assign P1_U4521 = ~(P1_U4252 & P1_U4261); 
assign P1_U4536 = ~P1_U3321; 
assign P1_U4604 = ~P1_U3328; 
assign P1_U4662 = ~P1_U3335; 
assign P1_U4720 = ~P1_U3339; 
assign P1_U4777 = ~P1_U3344; 
assign P1_U4835 = ~P1_U3348; 
assign P1_U4892 = ~P1_U3351; 
assign P1_U4950 = ~P1_U3355; 
assign P1_U5235 = ~P1_U3375; 
assign P1_U5293 = ~P1_U3379; 
assign P1_U5350 = ~P1_U3382; 
assign P1_U5408 = ~P1_U3386; 
assign P1_U5507 = ~(P1_U4252 & P1_U3438); 
assign P1_U5516 = ~(P1_U4252 & P1_U3401); 
assign P1_U5527 = ~(P1_U5519 & P1_U4252); 
assign P1_U5532 = ~(P1_U4252 & P1_U3266); 
assign P1_U5960 = ~(P1_U2382 & P1_EAX_REG_15__SCAN_IN); 
assign P1_U5961 = ~(U340 & P1_U2381); 
assign P1_U5963 = ~(P1_U2382 & P1_EAX_REG_14__SCAN_IN); 
assign P1_U5964 = ~(U341 & P1_U2381); 
assign P1_U5966 = ~(P1_U2382 & P1_EAX_REG_13__SCAN_IN); 
assign P1_U5967 = ~(U342 & P1_U2381); 
assign P1_U5969 = ~(P1_U2382 & P1_EAX_REG_12__SCAN_IN); 
assign P1_U5970 = ~(U343 & P1_U2381); 
assign P1_U5972 = ~(P1_U2382 & P1_EAX_REG_11__SCAN_IN); 
assign P1_U5973 = ~(U344 & P1_U2381); 
assign P1_U5975 = ~(P1_U2382 & P1_EAX_REG_10__SCAN_IN); 
assign P1_U5976 = ~(U345 & P1_U2381); 
assign P1_U5978 = ~(P1_U2382 & P1_EAX_REG_9__SCAN_IN); 
assign P1_U5979 = ~(U315 & P1_U2381); 
assign P1_U5981 = ~(P1_U2382 & P1_EAX_REG_8__SCAN_IN); 
assign P1_U5982 = ~(U316 & P1_U2381); 
assign P1_U5984 = ~(P1_U2382 & P1_EAX_REG_7__SCAN_IN); 
assign P1_U5985 = ~(P1_U2381 & U317); 
assign P1_U5987 = ~(P1_U2382 & P1_EAX_REG_6__SCAN_IN); 
assign P1_U5988 = ~(P1_U2381 & U318); 
assign P1_U5990 = ~(P1_U2382 & P1_EAX_REG_5__SCAN_IN); 
assign P1_U5991 = ~(P1_U2381 & U319); 
assign P1_U5993 = ~(P1_U2382 & P1_EAX_REG_4__SCAN_IN); 
assign P1_U5994 = ~(P1_U2381 & U320); 
assign P1_U5996 = ~(P1_U2382 & P1_EAX_REG_3__SCAN_IN); 
assign P1_U5997 = ~(P1_U2381 & U321); 
assign P1_U5999 = ~(P1_U2382 & P1_EAX_REG_2__SCAN_IN); 
assign P1_U6000 = ~(P1_U2381 & U324); 
assign P1_U6002 = ~(P1_U2382 & P1_EAX_REG_1__SCAN_IN); 
assign P1_U6003 = ~(P1_U2381 & U335); 
assign P1_U6005 = ~(P1_U2382 & P1_EAX_REG_0__SCAN_IN); 
assign P1_U6006 = ~(P1_U2381 & U346); 
assign P1_U6008 = ~(P1_U2382 & P1_EAX_REG_30__SCAN_IN); 
assign P1_U6009 = ~(U341 & P1_U2381); 
assign P1_U6011 = ~(P1_U2382 & P1_EAX_REG_29__SCAN_IN); 
assign P1_U6012 = ~(U342 & P1_U2381); 
assign P1_U6014 = ~(P1_U2382 & P1_EAX_REG_28__SCAN_IN); 
assign P1_U6015 = ~(U343 & P1_U2381); 
assign P1_U6017 = ~(P1_U2382 & P1_EAX_REG_27__SCAN_IN); 
assign P1_U6018 = ~(U344 & P1_U2381); 
assign P1_U6020 = ~(P1_U2382 & P1_EAX_REG_26__SCAN_IN); 
assign P1_U6021 = ~(U345 & P1_U2381); 
assign P1_U6023 = ~(P1_U2382 & P1_EAX_REG_25__SCAN_IN); 
assign P1_U6024 = ~(U315 & P1_U2381); 
assign P1_U6026 = ~(P1_U2382 & P1_EAX_REG_24__SCAN_IN); 
assign P1_U6027 = ~(U316 & P1_U2381); 
assign P1_U6029 = ~(P1_U2382 & P1_EAX_REG_23__SCAN_IN); 
assign P1_U6030 = ~(P1_U2381 & U317); 
assign P1_U6032 = ~(P1_U2382 & P1_EAX_REG_22__SCAN_IN); 
assign P1_U6033 = ~(P1_U2381 & U318); 
assign P1_U6035 = ~(P1_U2382 & P1_EAX_REG_21__SCAN_IN); 
assign P1_U6036 = ~(P1_U2381 & U319); 
assign P1_U6038 = ~(P1_U2382 & P1_EAX_REG_20__SCAN_IN); 
assign P1_U6039 = ~(P1_U2381 & U320); 
assign P1_U6041 = ~(P1_U2382 & P1_EAX_REG_19__SCAN_IN); 
assign P1_U6042 = ~(P1_U2381 & U321); 
assign P1_U6044 = ~(P1_U2382 & P1_EAX_REG_18__SCAN_IN); 
assign P1_U6045 = ~(P1_U2381 & U324); 
assign P1_U6047 = ~(P1_U2382 & P1_EAX_REG_17__SCAN_IN); 
assign P1_U6048 = ~(P1_U2381 & U335); 
assign P1_U6050 = ~(P1_U2382 & P1_EAX_REG_16__SCAN_IN); 
assign P1_U6051 = ~(P1_U2381 & U346); 
assign P1_U6053 = ~(P1_U4235 & P1_U7606 & P1_U4259); 
assign P1_U6152 = ~(P1_U7503 & P1_U3257); 
assign P1_U6264 = ~(P1_U4205 & P1_U6263); 
assign P1_U6616 = ~(P1_U4499 & P1_U3969 & P1_U3406); 
assign P1_U6771 = ~(P1_R2182_U26 & P1_U6746); 
assign P1_U7498 = ~(P1_U2425 & P1_U7493); 
assign P1_U7499 = ~(P1_U2425 & P1_U7493); 
assign P1_U7542 = ~(P1_U7541 & P1_UWORD_REG_0__SCAN_IN); 
assign P1_U7544 = ~(P1_U7543 & P1_UWORD_REG_1__SCAN_IN); 
assign P1_U7546 = ~(P1_U7545 & P1_UWORD_REG_2__SCAN_IN); 
assign P1_U7548 = ~(P1_U7547 & P1_UWORD_REG_3__SCAN_IN); 
assign P1_U7550 = ~(P1_U7549 & P1_UWORD_REG_4__SCAN_IN); 
assign P1_U7552 = ~(P1_U7551 & P1_UWORD_REG_5__SCAN_IN); 
assign P1_U7554 = ~(P1_U7553 & P1_UWORD_REG_6__SCAN_IN); 
assign P1_U7556 = ~(P1_U7555 & P1_UWORD_REG_7__SCAN_IN); 
assign P1_U7558 = ~(P1_U7557 & P1_UWORD_REG_8__SCAN_IN); 
assign P1_U7560 = ~(P1_U7559 & P1_UWORD_REG_9__SCAN_IN); 
assign P1_U7562 = ~(P1_U7561 & P1_UWORD_REG_10__SCAN_IN); 
assign P1_U7564 = ~(P1_U7563 & P1_UWORD_REG_11__SCAN_IN); 
assign P1_U7566 = ~(P1_U7565 & P1_UWORD_REG_12__SCAN_IN); 
assign P1_U7568 = ~(P1_U7567 & P1_UWORD_REG_13__SCAN_IN); 
assign P1_U7570 = ~(P1_U7569 & P1_UWORD_REG_14__SCAN_IN); 
assign P1_U7572 = ~(P1_U7571 & P1_LWORD_REG_0__SCAN_IN); 
assign P1_U7574 = ~(P1_U7573 & P1_LWORD_REG_1__SCAN_IN); 
assign P1_U7576 = ~(P1_U7575 & P1_LWORD_REG_2__SCAN_IN); 
assign P1_U7578 = ~(P1_U7577 & P1_LWORD_REG_3__SCAN_IN); 
assign P1_U7580 = ~(P1_U7579 & P1_LWORD_REG_4__SCAN_IN); 
assign P1_U7582 = ~(P1_U7581 & P1_LWORD_REG_5__SCAN_IN); 
assign P1_U7584 = ~(P1_U7583 & P1_LWORD_REG_6__SCAN_IN); 
assign P1_U7586 = ~(P1_U7585 & P1_LWORD_REG_7__SCAN_IN); 
assign P1_U7588 = ~(P1_U7587 & P1_LWORD_REG_8__SCAN_IN); 
assign P1_U7590 = ~(P1_U7589 & P1_LWORD_REG_9__SCAN_IN); 
assign P1_U7592 = ~(P1_U7591 & P1_LWORD_REG_10__SCAN_IN); 
assign P1_U7594 = ~(P1_U7593 & P1_LWORD_REG_11__SCAN_IN); 
assign P1_U7596 = ~(P1_U7595 & P1_LWORD_REG_12__SCAN_IN); 
assign P1_U7598 = ~(P1_U7597 & P1_LWORD_REG_13__SCAN_IN); 
assign P1_U7600 = ~(P1_U7599 & P1_LWORD_REG_14__SCAN_IN); 
assign P1_U7602 = ~(P1_U7601 & P1_LWORD_REG_15__SCAN_IN); 
assign P1_U7603 = ~(P1_U7493 & P1_U3568 & P1_U4259); 
assign P1_U7742 = ~(P1_U7741 & P1_U7740 & P1_U3257 & P1_U4171); 
assign P3_ADD_526_U63 = ~(P3_ADD_526_U166 & P3_ADD_526_U165); 
assign P3_ADD_526_U64 = ~(P3_ADD_526_U168 & P3_ADD_526_U167); 
assign P3_ADD_526_U123 = ~P3_ADD_526_U48; 
assign P3_ADD_526_U131 = ~P3_ADD_526_U101; 
assign P3_ADD_526_U162 = ~(P3_ADD_526_U48 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_526_U163 = ~(P3_ADD_526_U101 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_552_U63 = ~(P3_ADD_552_U166 & P3_ADD_552_U165); 
assign P3_ADD_552_U64 = ~(P3_ADD_552_U168 & P3_ADD_552_U167); 
assign P3_ADD_552_U123 = ~P3_ADD_552_U48; 
assign P3_ADD_552_U131 = ~P3_ADD_552_U101; 
assign P3_ADD_552_U162 = ~(P3_ADD_552_U48 & P3_EBX_REG_29__SCAN_IN); 
assign P3_ADD_552_U163 = ~(P3_ADD_552_U101 & P3_EBX_REG_28__SCAN_IN); 
assign P3_ADD_546_U63 = ~(P3_ADD_546_U166 & P3_ADD_546_U165); 
assign P3_ADD_546_U64 = ~(P3_ADD_546_U168 & P3_ADD_546_U167); 
assign P3_ADD_546_U123 = ~P3_ADD_546_U48; 
assign P3_ADD_546_U131 = ~P3_ADD_546_U101; 
assign P3_ADD_546_U162 = ~(P3_ADD_546_U48 & P3_EAX_REG_29__SCAN_IN); 
assign P3_ADD_546_U163 = ~(P3_ADD_546_U101 & P3_EAX_REG_28__SCAN_IN); 
assign P3_ADD_476_U86 = ~(P3_ADD_476_U172 & P3_ADD_476_U171); 
assign P3_ADD_476_U107 = ~P3_ADD_476_U32; 
assign P3_ADD_476_U169 = ~(P3_ADD_476_U32 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_531_U91 = ~(P3_ADD_531_U181 & P3_ADD_531_U180); 
assign P3_ADD_531_U111 = ~P3_ADD_531_U33; 
assign P3_ADD_531_U178 = ~(P3_ADD_531_U33 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_SUB_320_U30 = ~(P3_SUB_320_U47 & P3_SUB_320_U79 & P3_SUB_320_U94); 
assign P3_ADD_318_U86 = ~(P3_ADD_318_U172 & P3_ADD_318_U171); 
assign P3_ADD_318_U107 = ~P3_ADD_318_U32; 
assign P3_ADD_318_U169 = ~(P3_ADD_318_U32 & P3_PHYADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_315_U82 = ~(P3_ADD_315_U164 & P3_ADD_315_U163); 
assign P3_ADD_315_U104 = ~P3_ADD_315_U32; 
assign P3_ADD_315_U161 = ~(P3_ADD_315_U32 & P3_PHYADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_360_1242_U87 = ~(P3_ADD_360_1242_U208 & P3_ADD_360_1242_U207); 
assign P3_ADD_360_1242_U144 = ~P3_ADD_360_1242_U108; 
assign P3_ADD_360_1242_U146 = ~(P3_ADD_360_1242_U145 & P3_ADD_360_1242_U108); 
assign P3_ADD_360_1242_U200 = ~(P3_ADD_360_1242_U107 & P3_ADD_360_1242_U108); 
assign P3_ADD_467_U86 = ~(P3_ADD_467_U172 & P3_ADD_467_U171); 
assign P3_ADD_467_U107 = ~P3_ADD_467_U32; 
assign P3_ADD_467_U169 = ~(P3_ADD_467_U32 & P3_REIP_REG_16__SCAN_IN); 
assign P3_ADD_430_U86 = ~(P3_ADD_430_U172 & P3_ADD_430_U171); 
assign P3_ADD_430_U107 = ~P3_ADD_430_U32; 
assign P3_ADD_430_U169 = ~(P3_ADD_430_U32 & P3_REIP_REG_16__SCAN_IN); 
assign P3_ADD_380_U91 = ~(P3_ADD_380_U181 & P3_ADD_380_U180); 
assign P3_ADD_380_U111 = ~P3_ADD_380_U33; 
assign P3_ADD_380_U178 = ~(P3_ADD_380_U33 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_344_U91 = ~(P3_ADD_344_U181 & P3_ADD_344_U180); 
assign P3_ADD_344_U111 = ~P3_ADD_344_U33; 
assign P3_ADD_344_U178 = ~(P3_ADD_344_U33 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_LT_563_U10 = ~P3_U3306; 
assign P3_LT_563_U13 = ~P3_U3305; 
assign P3_LT_563_U15 = ~P3_U3308; 
assign P3_LT_563_U20 = ~(P3_U3306 & P3_LT_563_U11); 
assign P3_LT_563_U25 = ~(P3_U3305 & P3_LT_563_U12); 
assign P3_ADD_339_U86 = ~(P3_ADD_339_U172 & P3_ADD_339_U171); 
assign P3_ADD_339_U107 = ~P3_ADD_339_U32; 
assign P3_ADD_339_U169 = ~(P3_ADD_339_U32 & P3_PHYADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_541_U86 = ~(P3_ADD_541_U172 & P3_ADD_541_U171); 
assign P3_ADD_541_U107 = ~P3_ADD_541_U32; 
assign P3_ADD_541_U169 = ~(P3_ADD_541_U32 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_SUB_357_1258_U115 = ~(P3_SUB_357_1258_U176 & P3_SUB_357_1258_U152 & P3_SUB_357_1258_U268); 
assign P3_SUB_357_1258_U319 = ~(P3_SUB_357_1258_U301 & P3_SUB_357_1258_U317); 
assign P3_SUB_563_U6 = ~P3_U3305; 
assign P3_SUB_563_U7 = ~P3_U3306; 
assign P3_ADD_515_U86 = ~(P3_ADD_515_U172 & P3_ADD_515_U171); 
assign P3_ADD_515_U107 = ~P3_ADD_515_U32; 
assign P3_ADD_515_U169 = ~(P3_ADD_515_U32 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_394_U86 = ~(P3_ADD_394_U176 & P3_ADD_394_U175); 
assign P3_ADD_394_U110 = ~P3_ADD_394_U32; 
assign P3_ADD_394_U173 = ~(P3_ADD_394_U32 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_SUB_414_U64 = P3_SUB_414_U141 & P3_SUB_414_U140; 
assign P3_SUB_414_U102 = ~P3_SUB_414_U37; 
assign P3_SUB_414_U106 = ~(P3_SUB_414_U37 & P3_EBX_REG_29__SCAN_IN); 
assign P3_SUB_414_U108 = ~(P3_SUB_414_U107 & P3_EBX_REG_28__SCAN_IN); 
assign P3_ADD_441_U86 = ~(P3_ADD_441_U172 & P3_ADD_441_U171); 
assign P3_ADD_441_U107 = ~P3_ADD_441_U32; 
assign P3_ADD_441_U169 = ~(P3_ADD_441_U32 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_349_U91 = ~(P3_ADD_349_U181 & P3_ADD_349_U180); 
assign P3_ADD_349_U111 = ~P3_ADD_349_U33; 
assign P3_ADD_349_U178 = ~(P3_ADD_349_U33 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_405_U86 = ~(P3_ADD_405_U176 & P3_ADD_405_U175); 
assign P3_ADD_405_U110 = ~P3_ADD_405_U32; 
assign P3_ADD_405_U173 = ~(P3_ADD_405_U32 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_553_U91 = ~(P3_ADD_553_U181 & P3_ADD_553_U180); 
assign P3_ADD_553_U111 = ~P3_ADD_553_U33; 
assign P3_ADD_553_U178 = ~(P3_ADD_553_U33 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_558_U91 = ~(P3_ADD_558_U181 & P3_ADD_558_U180); 
assign P3_ADD_558_U111 = ~P3_ADD_558_U33; 
assign P3_ADD_558_U178 = ~(P3_ADD_558_U33 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_385_U91 = ~(P3_ADD_385_U181 & P3_ADD_385_U180); 
assign P3_ADD_385_U111 = ~P3_ADD_385_U33; 
assign P3_ADD_385_U178 = ~(P3_ADD_385_U33 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_547_U91 = ~(P3_ADD_547_U181 & P3_ADD_547_U180); 
assign P3_ADD_547_U111 = ~P3_ADD_547_U33; 
assign P3_ADD_547_U178 = ~(P3_ADD_547_U33 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_371_1212_U111 = ~(P3_ADD_371_1212_U144 & P3_ADD_371_1212_U118 & P3_ADD_371_1212_U200); 
assign P3_ADD_371_1212_U219 = ~(P3_ADD_371_1212_U143 & P3_ADD_371_1212_U217); 
assign P3_ADD_494_U86 = ~(P3_ADD_494_U172 & P3_ADD_494_U171); 
assign P3_ADD_494_U107 = ~P3_ADD_494_U32; 
assign P3_ADD_494_U169 = ~(P3_ADD_494_U32 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_536_U86 = ~(P3_ADD_536_U172 & P3_ADD_536_U171); 
assign P3_ADD_536_U107 = ~P3_ADD_536_U32; 
assign P3_ADD_536_U169 = ~(P3_ADD_536_U32 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P2_R2099_U17 = ~(P2_U2742 & P2_R2099_U120); 
assign P2_R2099_U98 = P2_R2099_U160 & P2_R2099_U159; 
assign P2_R2099_U158 = ~(P2_R2099_U120 & P2_R2099_U16); 
assign P2_ADD_391_1196_U87 = ~(P2_ADD_391_1196_U478 & P2_ADD_391_1196_U477); 
assign P2_ADD_391_1196_U143 = ~(P2_R2096_U51 & P2_ADD_391_1196_U162); 
assign P2_R2182_U100 = P2_R2182_U191 & P2_R2182_U125; 
assign P2_R2182_U126 = ~(P2_R2182_U125 & P2_R2182_U123 & P2_R2182_U124); 
assign P2_R2182_U222 = ~(P2_U2679 & P2_R2182_U42); 
assign P2_R2182_U224 = ~(P2_U2659 & P2_R2182_U64); 
assign P2_R2182_U226 = ~(P2_U2659 & P2_R2182_U64); 
assign P2_R2182_U282 = ~(P2_R2182_U281 & P2_U2701); 
assign P2_R2167_U32 = ~(P2_R2167_U30 & P2_R2167_U29 & P2_R2167_U31); 
assign P2_R2167_U39 = ~(P2_U2361 & P2_R2167_U18); 
assign P2_R2167_U41 = ~(P2_U2361 & P2_R2167_U18 & P2_STATE2_REG_0__SCAN_IN); 
assign P2_R2027_U91 = ~(P2_R2027_U181 & P2_R2027_U180); 
assign P2_R2027_U111 = ~P2_R2027_U33; 
assign P2_R2027_U178 = ~(P2_R2027_U33 & P2_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P2_R2337_U84 = ~(P2_R2337_U170 & P2_R2337_U169); 
assign P2_R2337_U108 = ~P2_R2337_U33; 
assign P2_R2337_U167 = ~(P2_R2337_U33 & P2_PHYADDRPOINTER_REG_17__SCAN_IN); 
assign P2_R2096_U72 = ~(P2_R2096_U188 & P2_R2096_U187); 
assign P2_R2096_U139 = ~P2_R2096_U101; 
assign P2_R2096_U141 = ~(P2_R2096_U140 & P2_R2096_U101); 
assign P2_R2096_U180 = ~(P2_R2096_U100 & P2_R2096_U101); 
assign P2_R1957_U29 = ~(P2_R1957_U94 & P2_R1957_U79 & P2_R1957_U46); 
assign P2_ADD_394_U75 = ~(P2_ADD_394_U152 & P2_ADD_394_U151); 
assign P2_ADD_394_U110 = ~P2_ADD_394_U32; 
assign P2_ADD_394_U185 = ~(P2_ADD_394_U32 & P2_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P2_R2267_U25 = ~(P2_R2267_U90 & P2_R2267_U59 & P2_R2267_U28); 
assign P2_R2267_U57 = ~P2_U3640; 
assign P2_R2267_U98 = ~(P2_R2267_U90 & P2_R2267_U59); 
assign P2_R2267_U140 = ~(P2_R2267_U90 & P2_R2267_U59); 
assign P1_R2027_U63 = ~(P1_R2027_U166 & P1_R2027_U165); 
assign P1_R2027_U64 = ~(P1_R2027_U168 & P1_R2027_U167); 
assign P1_R2027_U123 = ~P1_R2027_U48; 
assign P1_R2027_U131 = ~P1_R2027_U101; 
assign P1_R2027_U162 = ~(P1_R2027_U48 & P1_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P1_R2027_U163 = ~(P1_R2027_U101 & P1_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P1_R2144_U100 = ~(P1_U2751 & P1_R2144_U28); 
assign P1_R2144_U109 = ~(P1_R2144_U194 & P1_R2144_U193 & P1_R2144_U13); 
assign P1_R2144_U184 = ~(P1_R2144_U183 & P1_R2144_U182); 
assign P1_R2144_U187 = ~P1_R2144_U28; 
assign P1_R2144_U195 = ~(P1_U2355 & P1_R2144_U75); 
assign P1_R2144_U197 = ~(P1_U2355 & P1_R2144_U75); 
assign P1_R2144_U241 = ~(P1_R2144_U28 & P1_R2144_U14); 
assign P1_R2144_U243 = ~(P1_R2144_U28 & P1_R2144_U14); 
assign P1_R2144_U260 = ~(P1_R2144_U148 & P1_R2144_U12); 
assign P1_R2358_U411 = ~(P1_U2352 & P1_R2358_U147); 
assign P1_R2358_U416 = ~(P1_R2358_U415 & P1_R2358_U414); 
assign P1_R2358_U424 = ~(P1_R2358_U423 & P1_R2358_U422); 
assign P1_R2358_U437 = ~(P1_U2352 & P1_R2358_U151); 
assign P1_R2358_U439 = ~(P1_U2352 & P1_R2358_U151); 
assign P1_R2358_U442 = ~(P1_U2352 & P1_R2358_U147); 
assign P1_R2358_U461 = ~(P1_U2352 & P1_R2358_U159); 
assign P1_R2358_U467 = ~(P1_U2352 & P1_R2358_U159); 
assign P1_R2099_U36 = ~(P1_R2099_U213 & P1_R2099_U212); 
assign P1_R2099_U85 = ~(P1_R2099_U344 & P1_R2099_U343); 
assign P1_R2099_U162 = ~P1_R2099_U144; 
assign P1_R2099_U163 = ~P1_R2099_U11; 
assign P1_R2099_U340 = ~(P1_R2099_U60 & P1_R2099_U11); 
assign P1_R2099_U342 = ~(P1_R2099_U63 & P1_R2099_U144); 
assign P1_R2337_U86 = ~(P1_R2337_U172 & P1_R2337_U171); 
assign P1_R2337_U107 = ~P1_R2337_U32; 
assign P1_R2337_U169 = ~(P1_R2337_U32 & P1_PHYADDRPOINTER_REG_16__SCAN_IN); 
assign P1_R2096_U86 = ~(P1_R2096_U172 & P1_R2096_U171); 
assign P1_R2096_U107 = ~P1_R2096_U32; 
assign P1_R2096_U169 = ~(P1_R2096_U32 & P1_REIP_REG_16__SCAN_IN); 
assign P1_ADD_405_U75 = ~(P1_ADD_405_U152 & P1_ADD_405_U151); 
assign P1_ADD_405_U110 = ~P1_ADD_405_U32; 
assign P1_ADD_405_U185 = ~(P1_ADD_405_U32 & P1_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P1_ADD_515_U75 = ~(P1_ADD_515_U150 & P1_ADD_515_U149); 
assign P1_ADD_515_U107 = ~P1_ADD_515_U32; 
assign P1_ADD_515_U181 = ~(P1_ADD_515_U32 & P1_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_U2858 = ~(P3_U5751 & P3_U5749 & P3_U5750); 
assign P3_U3285 = ~(P3_U7980 & P3_U7979); 
assign P3_U3288 = ~(P3_U7990 & P3_U7989); 
assign P3_U3289 = ~(P3_U7992 & P3_U7991); 
assign P3_U3290 = ~(P3_U7996 & P3_U7995); 
assign P3_U3745 = P3_U3744 & P3_U3743 & P3_U5795; 
assign P3_U3960 = P3_U6458 & P3_U6457 & P3_U6460 & P3_U6459; 
assign P3_U5774 = ~(P3_U4318 & P3_U5772); 
assign P3_U5800 = ~(P3_ADD_360_1242_U87 & P3_U2395); 
assign P3_U5970 = ~(P3_ADD_558_U91 & P3_U3220); 
assign P3_U5971 = ~(P3_ADD_553_U91 & P3_U4298); 
assign P3_U5972 = ~(P3_ADD_547_U91 & P3_U4299); 
assign P3_U5975 = ~(P3_ADD_531_U91 & P3_U2354); 
assign P3_U5983 = ~(P3_ADD_385_U91 & P3_U2358); 
assign P3_U5984 = ~(P3_ADD_380_U91 & P3_U2359); 
assign P3_U5985 = ~(P3_ADD_349_U91 & P3_U4306); 
assign P3_U5986 = ~(P3_ADD_344_U91 & P3_U2362); 
assign P3_U5997 = ~(P3_ADD_541_U86 & P3_U4300); 
assign P3_U5998 = ~(P3_ADD_536_U86 & P3_U4301); 
assign P3_U6001 = ~(P3_ADD_515_U86 & P3_U4302); 
assign P3_U6002 = ~(P3_ADD_494_U86 & P3_U2356); 
assign P3_U6003 = ~(P3_ADD_476_U86 & P3_U4303); 
assign P3_U6004 = ~(P3_ADD_441_U86 & P3_U4304); 
assign P3_U6005 = ~(P3_ADD_405_U86 & P3_U4305); 
assign P3_U6006 = ~(P3_ADD_394_U86 & P3_U2357); 
assign P3_U6264 = ~(P3_ADD_526_U64 & P3_U2355); 
assign P3_U6288 = ~(P3_ADD_526_U63 & P3_U2355); 
assign P3_U6463 = ~(P3_U2396 & P3_ADD_360_1242_U87); 
assign P3_U6525 = ~(P3_ADD_318_U86 & P3_U2398); 
assign P3_U6530 = ~(P3_ADD_339_U86 & P3_U2388); 
assign P3_U6534 = ~(P3_ADD_315_U82 & P3_U2397); 
assign P3_U6971 = ~(P3_ADD_546_U64 & P3_U2400); 
assign P3_U6976 = ~(P3_ADD_546_U63 & P3_U2400); 
assign P3_U7077 = ~(P3_ADD_552_U64 & P3_U2399); 
assign P3_U7080 = ~(P3_ADD_552_U63 & P3_U2399); 
assign P3_U7230 = ~(P3_ADD_467_U86 & P3_U2601); 
assign P3_U7232 = ~(P3_ADD_430_U86 & P3_U2405); 
assign P3_U7325 = ~(P3_SUB_414_U64 & P3_U2602); 
assign P2_U3326 = ~(P2_U3570 & P2_U3312); 
assign P2_U3340 = ~(P2_U3569 & P2_U3336); 
assign P2_U3356 = ~(P2_U3568 & P2_U3350); 
assign P2_U3367 = ~(P2_U3567 & P2_U3365); 
assign P2_U3381 = ~(P2_U3566 & P2_U3377); 
assign P2_U3392 = ~(P2_U3565 & P2_U3390); 
assign P2_U3404 = ~(P2_U3564 & P2_U3401); 
assign P2_U3415 = ~(P2_U3563 & P2_U3413); 
assign P2_U3476 = ~(P2_U3558 & P2_U3473); 
assign P2_U3487 = ~(P2_U3557 & P2_U3485); 
assign P2_U3499 = ~(P2_U3556 & P2_U3496); 
assign P2_U3510 = ~(P2_U3555 & P2_U3508); 
assign P2_U3559 = ~(P2_U2492 & P2_U2479); 
assign P2_U3560 = ~(P2_U2492 & P2_U2473); 
assign P2_U3561 = ~(P2_U2492 & P2_U2470); 
assign P2_U3562 = ~(P2_U2492 & P2_U2467); 
assign P2_U3639 = ~(P2_U8332 & P2_U8331); 
assign P2_U4653 = ~P2_U3570; 
assign P2_U4713 = ~P2_U3569; 
assign P2_U4772 = ~P2_U3568; 
assign P2_U4829 = ~P2_U3567; 
assign P2_U4887 = ~P2_U3566; 
assign P2_U4944 = ~P2_U3565; 
assign P2_U5002 = ~P2_U3564; 
assign P2_U5059 = ~P2_U3563; 
assign P2_U5345 = ~P2_U3558; 
assign P2_U5402 = ~P2_U3557; 
assign P2_U5460 = ~P2_U3556; 
assign P2_U5517 = ~P2_U3555; 
assign P2_U5613 = ~(P2_U4466 & P2_U5611); 
assign P2_U8405 = ~(P2_R2337_U84 & P2_U3284); 
assign P1_U2364 = P1_U3864 & P1_U3416; 
assign P1_U2365 = P1_U4261 & P1_U3416; 
assign P1_U2372 = P1_U3416 & P1_STATE2_REG_0__SCAN_IN; 
assign P1_U2376 = P1_U5798 & P1_U3416; 
assign P1_U3285 = ~(P1_U2473 & P1_U4501); 
assign P1_U3417 = ~(P1_U6054 & P1_U6053); 
assign P1_U3426 = ~(P1_U4235 & P1_U6264); 
assign P1_U3581 = P1_U7603 & P1_STATE2_REG_2__SCAN_IN; 
assign P1_U4178 = ~(P1_U4508 & P1_U3391); 
assign P1_U4224 = ~P1_U3300; 
assign P1_U5006 = ~P1_U3361; 
assign P1_U5063 = ~P1_U3365; 
assign P1_U5120 = ~P1_U3368; 
assign P1_U5178 = ~P1_U3372; 
assign P1_U5473 = ~P1_U4182; 
assign P1_U5474 = ~(P1_U2368 & P1_U4182); 
assign P1_U5509 = ~(P1_U5508 & P1_U5507); 
assign P1_U5518 = ~(P1_U5517 & P1_U5515 & P1_U5516); 
assign P1_U5529 = ~(P1_U5528 & P1_U5526 & P1_U5527); 
assign P1_U5535 = ~(P1_U5533 & P1_U5534 & P1_U5532); 
assign P1_U5559 = ~(P1_U4260 & P1_U2431); 
assign P1_U5795 = ~P1_U3416; 
assign P1_U5962 = ~(P1_U5961 & P1_U5960); 
assign P1_U5965 = ~(P1_U5964 & P1_U5963); 
assign P1_U5968 = ~(P1_U5967 & P1_U5966); 
assign P1_U5971 = ~(P1_U5970 & P1_U5969); 
assign P1_U5974 = ~(P1_U5973 & P1_U5972); 
assign P1_U5977 = ~(P1_U5976 & P1_U5975); 
assign P1_U5980 = ~(P1_U5979 & P1_U5978); 
assign P1_U5983 = ~(P1_U5982 & P1_U5981); 
assign P1_U5986 = ~(P1_U5985 & P1_U5984); 
assign P1_U5989 = ~(P1_U5988 & P1_U5987); 
assign P1_U5992 = ~(P1_U5991 & P1_U5990); 
assign P1_U5995 = ~(P1_U5994 & P1_U5993); 
assign P1_U5998 = ~(P1_U5997 & P1_U5996); 
assign P1_U6001 = ~(P1_U6000 & P1_U5999); 
assign P1_U6004 = ~(P1_U6003 & P1_U6002); 
assign P1_U6007 = ~(P1_U6006 & P1_U6005); 
assign P1_U6010 = ~(P1_U6009 & P1_U6008); 
assign P1_U6013 = ~(P1_U6012 & P1_U6011); 
assign P1_U6016 = ~(P1_U6015 & P1_U6014); 
assign P1_U6019 = ~(P1_U6018 & P1_U6017); 
assign P1_U6022 = ~(P1_U6021 & P1_U6020); 
assign P1_U6025 = ~(P1_U6024 & P1_U6023); 
assign P1_U6028 = ~(P1_U6027 & P1_U6026); 
assign P1_U6031 = ~(P1_U6030 & P1_U6029); 
assign P1_U6034 = ~(P1_U6033 & P1_U6032); 
assign P1_U6037 = ~(P1_U6036 & P1_U6035); 
assign P1_U6040 = ~(P1_U6039 & P1_U6038); 
assign P1_U6043 = ~(P1_U6042 & P1_U6041); 
assign P1_U6046 = ~(P1_U6045 & P1_U6044); 
assign P1_U6049 = ~(P1_U6048 & P1_U6047); 
assign P1_U6052 = ~(P1_U6051 & P1_U6050); 
assign P1_U6153 = ~(P1_U3883 & P1_U6152); 
assign P1_U6610 = ~(P1_U2368 & P1_U2473); 
assign P1_U6617 = ~(P1_U6616 & P1_MEMORYFETCH_REG_SCAN_IN); 
assign P1_U6843 = ~(P1_R2337_U86 & P1_U2352); 
assign P1_U7500 = ~(P1_U6361 & P1_U6360 & P1_U7499); 
assign P1_U7774 = ~(P1_U3488 & P1_U4182); 
assign P1_U7777 = ~(P1_U5506 & P1_U4182); 
assign P1_U7779 = ~(P1_U5514 & P1_U4182); 
assign P1_U7781 = ~(P1_U5525 & P1_U4182); 
assign P1_U7783 = ~(P1_U5531 & P1_U4182); 
assign P3_ADD_526_U49 = ~(P3_ADD_526_U123 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_526_U161 = ~(P3_ADD_526_U123 & P3_ADD_526_U47); 
assign P3_ADD_526_U164 = ~(P3_ADD_526_U131 & P3_ADD_526_U45); 
assign P3_ADD_552_U49 = ~(P3_ADD_552_U123 & P3_EBX_REG_29__SCAN_IN); 
assign P3_ADD_552_U161 = ~(P3_ADD_552_U123 & P3_ADD_552_U47); 
assign P3_ADD_552_U164 = ~(P3_ADD_552_U131 & P3_ADD_552_U45); 
assign P3_ADD_546_U49 = ~(P3_ADD_546_U123 & P3_EAX_REG_29__SCAN_IN); 
assign P3_ADD_546_U161 = ~(P3_ADD_546_U123 & P3_ADD_546_U47); 
assign P3_ADD_546_U164 = ~(P3_ADD_546_U131 & P3_ADD_546_U45); 
assign P3_ADD_476_U34 = ~(P3_ADD_476_U107 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_476_U170 = ~(P3_ADD_476_U107 & P3_ADD_476_U33); 
assign P3_ADD_531_U35 = ~(P3_ADD_531_U111 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_531_U179 = ~(P3_ADD_531_U111 & P3_ADD_531_U34); 
assign P3_SUB_320_U8 = P3_SUB_320_U122 & P3_SUB_320_U30; 
assign P3_SUB_320_U77 = ~P3_ADD_318_U86; 
assign P3_SUB_320_U95 = ~P3_SUB_320_U30; 
assign P3_SUB_320_U154 = ~(P3_ADD_318_U86 & P3_SUB_320_U30); 
assign P3_ADD_318_U34 = ~(P3_ADD_318_U107 & P3_PHYADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_318_U170 = ~(P3_ADD_318_U107 & P3_ADD_318_U33); 
assign P3_ADD_315_U34 = ~(P3_ADD_315_U104 & P3_PHYADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_315_U162 = ~(P3_ADD_315_U104 & P3_ADD_315_U33); 
assign P3_ADD_360_1242_U105 = ~(P3_ADD_360_1242_U147 & P3_ADD_360_1242_U146); 
assign P3_ADD_360_1242_U201 = ~(P3_ADD_360_1242_U144 & P3_ADD_360_1242_U199); 
assign P3_LT_563_1260_U7 = ~(P3_SUB_563_U7 | P3_SUB_563_U6); 
assign P3_ADD_467_U34 = ~(P3_ADD_467_U107 & P3_REIP_REG_16__SCAN_IN); 
assign P3_ADD_467_U170 = ~(P3_ADD_467_U107 & P3_ADD_467_U33); 
assign P3_ADD_430_U34 = ~(P3_ADD_430_U107 & P3_REIP_REG_16__SCAN_IN); 
assign P3_ADD_430_U170 = ~(P3_ADD_430_U107 & P3_ADD_430_U33); 
assign P3_ADD_380_U35 = ~(P3_ADD_380_U111 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_380_U179 = ~(P3_ADD_380_U111 & P3_ADD_380_U34); 
assign P3_ADD_344_U35 = ~(P3_ADD_344_U111 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_344_U179 = ~(P3_ADD_344_U111 & P3_ADD_344_U34); 
assign P3_LT_563_U8 = ~(P3_LT_563_U15 & P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P3_LT_563_U22 = ~(P3_LT_563_U10 & P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P3_LT_563_U23 = ~(P3_LT_563_U13 & P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P3_ADD_339_U34 = ~(P3_ADD_339_U107 & P3_PHYADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_339_U170 = ~(P3_ADD_339_U107 & P3_ADD_339_U33); 
assign P3_ADD_541_U34 = ~(P3_ADD_541_U107 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_541_U170 = ~(P3_ADD_541_U107 & P3_ADD_541_U33); 
assign P3_SUB_357_1258_U71 = ~(P3_SUB_357_1258_U319 & P3_SUB_357_1258_U318); 
assign P3_SUB_357_1258_U177 = ~P3_SUB_357_1258_U115; 
assign P3_SUB_357_1258_U286 = ~(P3_SUB_357_1258_U178 & P3_SUB_357_1258_U115); 
assign P3_SUB_357_1258_U288 = ~(P3_SUB_357_1258_U6 & P3_SUB_357_1258_U115); 
assign P3_SUB_357_1258_U290 = ~(P3_SUB_357_1258_U7 & P3_SUB_357_1258_U115); 
assign P3_SUB_357_1258_U292 = ~(P3_SUB_357_1258_U98 & P3_SUB_357_1258_U115); 
assign P3_SUB_357_1258_U311 = ~(P3_SUB_357_1258_U258 & P3_SUB_357_1258_U115); 
assign P3_ADD_515_U34 = ~(P3_ADD_515_U107 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_515_U170 = ~(P3_ADD_515_U107 & P3_ADD_515_U33); 
assign P3_ADD_394_U34 = ~(P3_ADD_394_U110 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_394_U174 = ~(P3_ADD_394_U110 & P3_ADD_394_U33); 
assign P3_SUB_414_U15 = P3_SUB_414_U108 & P3_SUB_414_U37; 
assign P3_SUB_414_U38 = ~(P3_SUB_414_U102 & P3_SUB_414_U39); 
assign P3_ADD_441_U34 = ~(P3_ADD_441_U107 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_441_U170 = ~(P3_ADD_441_U107 & P3_ADD_441_U33); 
assign P3_ADD_349_U35 = ~(P3_ADD_349_U111 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_349_U179 = ~(P3_ADD_349_U111 & P3_ADD_349_U34); 
assign P3_ADD_405_U34 = ~(P3_ADD_405_U110 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_405_U174 = ~(P3_ADD_405_U110 & P3_ADD_405_U33); 
assign P3_ADD_553_U35 = ~(P3_ADD_553_U111 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_553_U179 = ~(P3_ADD_553_U111 & P3_ADD_553_U34); 
assign P3_ADD_558_U35 = ~(P3_ADD_558_U111 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_558_U179 = ~(P3_ADD_558_U111 & P3_ADD_558_U34); 
assign P3_ADD_385_U35 = ~(P3_ADD_385_U111 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_385_U179 = ~(P3_ADD_385_U111 & P3_ADD_385_U34); 
assign P3_ADD_547_U35 = ~(P3_ADD_547_U111 & P3_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P3_ADD_547_U179 = ~(P3_ADD_547_U111 & P3_ADD_547_U34); 
assign P3_ADD_371_1212_U89 = ~(P3_ADD_371_1212_U219 & P3_ADD_371_1212_U218); 
assign P3_ADD_371_1212_U145 = ~P3_ADD_371_1212_U111; 
assign P3_ADD_371_1212_U147 = ~(P3_ADD_371_1212_U146 & P3_ADD_371_1212_U111); 
assign P3_ADD_371_1212_U211 = ~(P3_ADD_371_1212_U110 & P3_ADD_371_1212_U111); 
assign P3_ADD_494_U34 = ~(P3_ADD_494_U107 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_494_U170 = ~(P3_ADD_494_U107 & P3_ADD_494_U33); 
assign P3_ADD_536_U34 = ~(P3_ADD_536_U107 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_536_U170 = ~(P3_ADD_536_U107 & P3_ADD_536_U33); 
assign P2_R2099_U71 = ~(P2_R2099_U158 & P2_R2099_U157); 
assign P2_R2099_U121 = ~P2_R2099_U17; 
assign P2_R2099_U155 = ~(P2_U2741 & P2_R2099_U17); 
assign P2_ADD_391_1196_U16 = ~P2_R2096_U72; 
assign P2_ADD_391_1196_U160 = ~P2_ADD_391_1196_U143; 
assign P2_R2182_U48 = ~P2_U2699; 
assign P2_R2182_U68 = ~(P2_R2182_U283 & P2_R2182_U282); 
assign P2_R2182_U99 = P2_R2182_U223 & P2_R2182_U222 & P2_R2182_U189; 
assign P2_R2182_U106 = ~(P2_R2182_U126 & P2_R2182_U127); 
assign P2_R2182_U108 = ~P2_U2682; 
assign P2_R2182_U109 = P2_R2182_U225 & P2_R2182_U224; 
assign P2_R2182_U129 = P2_U2699 | P2_U2678; 
assign P2_R2182_U131 = ~(P2_U2678 & P2_U2699); 
assign P2_R2182_U192 = ~(P2_R2182_U124 & P2_R2182_U123 & P2_R2182_U100); 
assign P2_R2182_U211 = ~(P2_U2699 & P2_R2182_U49); 
assign P2_R2182_U213 = ~(P2_U2699 & P2_R2182_U49); 
assign P2_R2182_U218 = ~(P2_U2682 & P2_R2182_U107); 
assign P2_R2182_U220 = ~(P2_U2682 & P2_R2182_U107); 
assign P2_R2182_U228 = ~(P2_R2182_U227 & P2_R2182_U226); 
assign P2_R2167_U35 = ~(P2_R2167_U33 & P2_R2167_U32 & P2_R2167_U34); 
assign P2_R2027_U35 = ~(P2_R2027_U111 & P2_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P2_R2027_U179 = ~(P2_R2027_U111 & P2_R2027_U34); 
assign P2_R2337_U35 = ~(P2_R2337_U108 & P2_PHYADDRPOINTER_REG_17__SCAN_IN); 
assign P2_R2337_U168 = ~(P2_R2337_U108 & P2_R2337_U34); 
assign P2_R2096_U99 = ~(P2_R2096_U142 & P2_R2096_U141); 
assign P2_R2096_U181 = ~(P2_R2096_U139 & P2_R2096_U179); 
assign P2_R1957_U8 = P2_R1957_U122 & P2_R1957_U29; 
assign P2_R1957_U77 = ~P2_U3676; 
assign P2_R1957_U95 = ~P2_R1957_U29; 
assign P2_R1957_U154 = ~(P2_U3676 & P2_R1957_U29); 
assign P2_ADD_394_U34 = ~(P2_ADD_394_U110 & P2_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P2_ADD_394_U186 = ~(P2_ADD_394_U110 & P2_ADD_394_U33); 
assign P2_R2267_U41 = ~P2_U2767; 
assign P2_R2267_U44 = ~(P2_U2789 | P2_U2788); 
assign P2_R2267_U45 = ~(P2_U2787 | P2_U2786); 
assign P2_R2267_U46 = ~(P2_U2785 | P2_U2784); 
assign P2_R2267_U47 = ~(P2_U2783 | P2_U2782); 
assign P2_R2267_U48 = ~(P2_U2781 | P2_U2780); 
assign P2_R2267_U49 = ~(P2_U2779 | P2_U2778); 
assign P2_R2267_U50 = ~(P2_U2777 | P2_U2776); 
assign P2_R2267_U51 = ~(P2_U2775 | P2_U2774); 
assign P2_R2267_U52 = ~(P2_U2773 | P2_U2772); 
assign P2_R2267_U53 = ~(P2_U2771 | P2_U2770); 
assign P2_R2267_U54 = ~(P2_U2769 | P2_U2768); 
assign P2_R2267_U55 = ~P2_U2789; 
assign P2_R2267_U60 = P2_R2267_U140 & P2_R2267_U139; 
assign P2_R2267_U61 = ~P2_U2766; 
assign P2_R2267_U66 = ~P2_U2769; 
assign P2_R2267_U68 = ~P2_U2771; 
assign P2_R2267_U70 = ~P2_U2773; 
assign P2_R2267_U72 = ~P2_U2775; 
assign P2_R2267_U74 = ~P2_U2777; 
assign P2_R2267_U78 = ~P2_U2779; 
assign P2_R2267_U80 = ~P2_U2781; 
assign P2_R2267_U82 = ~P2_U2783; 
assign P2_R2267_U84 = ~P2_U2785; 
assign P2_R2267_U86 = ~P2_U2787; 
assign P2_R2267_U91 = ~P2_R2267_U25; 
assign P2_R2267_U99 = ~(P2_U3641 & P2_R2267_U98); 
assign P2_R2267_U137 = ~(P2_U3640 & P2_R2267_U25); 
assign P1_R2027_U49 = ~(P1_R2027_U123 & P1_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P1_R2027_U161 = ~(P1_R2027_U123 & P1_R2027_U47); 
assign P1_R2027_U164 = ~(P1_R2027_U131 & P1_R2027_U45); 
assign P1_R2144_U43 = ~(P1_R2144_U260 & P1_R2144_U259); 
assign P1_R2144_U55 = P1_R2144_U109 & P1_R2144_U106; 
assign P1_R2144_U110 = ~(P1_R2144_U196 & P1_R2144_U195 & P1_R2144_U16); 
assign P1_R2144_U114 = ~(P1_R2144_U187 & P1_R2144_U14); 
assign P1_R2144_U116 = ~(P1_U2750 & P1_R2144_U184); 
assign P1_R2144_U131 = ~(P1_R2144_U187 & P1_R2144_U14); 
assign P1_R2144_U154 = ~(P1_R2144_U113 & P1_R2144_U115 & P1_R2144_U100); 
assign P1_R2144_U157 = ~(P1_U2750 & P1_R2144_U184); 
assign P1_R2144_U162 = ~(P1_U2750 & P1_R2144_U184); 
assign P1_R2144_U199 = ~(P1_R2144_U198 & P1_R2144_U197); 
assign P1_R2144_U240 = ~(P1_R2144_U187 & P1_U2751); 
assign P1_R2144_U242 = ~(P1_R2144_U187 & P1_U2751); 
assign P1_R2358_U158 = ~P1_U2612; 
assign P1_R2358_U413 = ~(P1_R2358_U412 & P1_R2358_U411); 
assign P1_R2358_U441 = ~(P1_R2358_U440 & P1_R2358_U439); 
assign P1_R2358_U460 = ~(P1_U2612 & P1_R2358_U23); 
assign P1_R2358_U463 = ~(P1_R2358_U462 & P1_R2358_U461); 
assign P1_R2358_U465 = ~(P1_U2612 & P1_R2358_U23); 
assign P1_R2099_U12 = ~(P1_R2099_U93 & P1_R2099_U163); 
assign P1_R2099_U143 = ~(P1_R2099_U163 & P1_R2099_U60); 
assign P1_R2099_U339 = ~(P1_R2099_U267 & P1_R2099_U163); 
assign P1_R2099_U341 = ~(P1_R2099_U162 & P1_R2099_U264); 
assign P1_R2337_U34 = ~(P1_R2337_U107 & P1_PHYADDRPOINTER_REG_16__SCAN_IN); 
assign P1_R2337_U170 = ~(P1_R2337_U107 & P1_R2337_U33); 
assign P1_R2096_U34 = ~(P1_R2096_U107 & P1_REIP_REG_16__SCAN_IN); 
assign P1_R2096_U170 = ~(P1_R2096_U107 & P1_R2096_U33); 
assign P1_ADD_405_U34 = ~(P1_ADD_405_U110 & P1_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P1_ADD_405_U186 = ~(P1_ADD_405_U110 & P1_ADD_405_U33); 
assign P1_ADD_515_U34 = ~(P1_ADD_515_U107 & P1_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P1_ADD_515_U182 = ~(P1_ADD_515_U107 & P1_ADD_515_U33); 
assign P3_U2676 = ~(P3_U7081 & P3_U7079 & P3_U7080); 
assign P3_U2677 = ~(P3_U7078 & P3_U7076 & P3_U7077); 
assign P3_U2708 = ~(P3_U6974 & P3_U6973 & P3_U4029 & P3_U6976); 
assign P3_U2709 = ~(P3_U6969 & P3_U6968 & P3_U4028 & P3_U6971); 
assign P3_U2824 = ~(P3_U6454 & P3_U6453 & P3_U6456 & P3_U6455 & P3_U3960); 
assign P3_U2857 = ~(P3_U5775 & P3_U5773 & P3_U5774); 
assign P3_U3746 = P3_U3747 & P3_U5800; 
assign P3_U3796 = P3_U5972 & P3_U5971; 
assign P3_U3798 = P3_U5974 & P3_U5973 & P3_U5975 & P3_U3797; 
assign P3_U3801 = P3_U5986 & P3_U5985 & P3_U5984 & P3_U5983; 
assign P3_U3805 = P3_U6001 & P3_U6000; 
assign P3_U3808 = P3_U6003 & P3_U6002 & P3_U6004 & P3_U6006 & P3_U6005; 
assign P3_U4084 = P3_U7229 & P3_U4316 & P3_U7230; 
assign P3_U5796 = ~(P3_U3742 & P3_U5778 & P3_U5777 & P3_U3738 & P3_U3745); 
assign P3_U5819 = ~(P3_ADD_371_1212_U89 & P3_U2360); 
assign P3_U5825 = ~(P3_SUB_357_1258_U71 & P3_U2393); 
assign P3_U6467 = ~(P3_U2387 & P3_ADD_371_1212_U89); 
assign P3_U6472 = ~(P3_U2394 & P3_SUB_357_1258_U71); 
assign P3_U7333 = ~(P3_SUB_414_U15 & P3_U2602); 
assign P2_U2476 = ~(P2_R2182_U69 | P2_R2182_U68); 
assign P2_U3315 = ~P2_R2182_U68; 
assign P2_U3318 = ~(P2_R2182_U68 & P2_R2182_U69); 
assign P2_U3337 = ~(P2_R2182_U68 & P2_U3314); 
assign P2_U3430 = ~(P2_U3562 & P2_U3424); 
assign P2_U3441 = ~(P2_U3561 & P2_U3439); 
assign P2_U3453 = ~(P2_U3560 & P2_U3450); 
assign P2_U3464 = ~(P2_U3559 & P2_U3462); 
assign P2_U3675 = ~(P2_U8406 & P2_U8405); 
assign P2_U4654 = ~P2_U3326; 
assign P2_U4667 = ~(P2_U3326 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U4714 = ~P2_U3340; 
assign P2_U4725 = ~(P2_U3340 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U4773 = ~P2_U3356; 
assign P2_U4784 = ~(P2_U3356 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U4830 = ~P2_U3367; 
assign P2_U4841 = ~(P2_U3367 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U4888 = ~P2_U3381; 
assign P2_U4899 = ~(P2_U3381 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U4945 = ~P2_U3392; 
assign P2_U4956 = ~(P2_U3392 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5003 = ~P2_U3404; 
assign P2_U5014 = ~(P2_U3404 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5060 = ~P2_U3415; 
assign P2_U5071 = ~(P2_U3415 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5116 = ~P2_U3562; 
assign P2_U5172 = ~P2_U3561; 
assign P2_U5230 = ~P2_U3560; 
assign P2_U5287 = ~P2_U3559; 
assign P2_U5346 = ~P2_U3476; 
assign P2_U5357 = ~(P2_U3476 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5403 = ~P2_U3487; 
assign P2_U5414 = ~(P2_U3487 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5461 = ~P2_U3499; 
assign P2_U5472 = ~(P2_U3499 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5518 = ~P2_U3510; 
assign P2_U5529 = ~(P2_U3510 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5658 = ~(P2_R2182_U68 & P2_U5644); 
assign P2_U7167 = ~(P2_U5517 & P2_INSTQUEUE_REG_0__7__SCAN_IN); 
assign P2_U7168 = ~(P2_U5460 & P2_INSTQUEUE_REG_1__7__SCAN_IN); 
assign P2_U7169 = ~(P2_U5402 & P2_INSTQUEUE_REG_2__7__SCAN_IN); 
assign P2_U7170 = ~(P2_U5345 & P2_INSTQUEUE_REG_3__7__SCAN_IN); 
assign P2_U7175 = ~(P2_U5059 & P2_INSTQUEUE_REG_8__7__SCAN_IN); 
assign P2_U7176 = ~(P2_U5002 & P2_INSTQUEUE_REG_9__7__SCAN_IN); 
assign P2_U7177 = ~(P2_U4944 & P2_INSTQUEUE_REG_10__7__SCAN_IN); 
assign P2_U7178 = ~(P2_U4887 & P2_INSTQUEUE_REG_11__7__SCAN_IN); 
assign P2_U7179 = ~(P2_U4829 & P2_INSTQUEUE_REG_12__7__SCAN_IN); 
assign P2_U7180 = ~(P2_U4772 & P2_INSTQUEUE_REG_13__7__SCAN_IN); 
assign P2_U7181 = ~(P2_U4713 & P2_INSTQUEUE_REG_14__7__SCAN_IN); 
assign P2_U7182 = ~(P2_U4653 & P2_INSTQUEUE_REG_15__7__SCAN_IN); 
assign P2_U7184 = ~(P2_U5517 & P2_INSTQUEUE_REG_0__6__SCAN_IN); 
assign P2_U7185 = ~(P2_U5460 & P2_INSTQUEUE_REG_1__6__SCAN_IN); 
assign P2_U7186 = ~(P2_U5402 & P2_INSTQUEUE_REG_2__6__SCAN_IN); 
assign P2_U7187 = ~(P2_U5345 & P2_INSTQUEUE_REG_3__6__SCAN_IN); 
assign P2_U7192 = ~(P2_U5059 & P2_INSTQUEUE_REG_8__6__SCAN_IN); 
assign P2_U7193 = ~(P2_U5002 & P2_INSTQUEUE_REG_9__6__SCAN_IN); 
assign P2_U7194 = ~(P2_U4944 & P2_INSTQUEUE_REG_10__6__SCAN_IN); 
assign P2_U7195 = ~(P2_U4887 & P2_INSTQUEUE_REG_11__6__SCAN_IN); 
assign P2_U7196 = ~(P2_U4829 & P2_INSTQUEUE_REG_12__6__SCAN_IN); 
assign P2_U7197 = ~(P2_U4772 & P2_INSTQUEUE_REG_13__6__SCAN_IN); 
assign P2_U7198 = ~(P2_U4713 & P2_INSTQUEUE_REG_14__6__SCAN_IN); 
assign P2_U7199 = ~(P2_U4653 & P2_INSTQUEUE_REG_15__6__SCAN_IN); 
assign P2_U7218 = ~(P2_U5517 & P2_INSTQUEUE_REG_0__5__SCAN_IN); 
assign P2_U7219 = ~(P2_U5460 & P2_INSTQUEUE_REG_1__5__SCAN_IN); 
assign P2_U7220 = ~(P2_U5402 & P2_INSTQUEUE_REG_2__5__SCAN_IN); 
assign P2_U7221 = ~(P2_U5345 & P2_INSTQUEUE_REG_3__5__SCAN_IN); 
assign P2_U7226 = ~(P2_U5059 & P2_INSTQUEUE_REG_8__5__SCAN_IN); 
assign P2_U7227 = ~(P2_U5002 & P2_INSTQUEUE_REG_9__5__SCAN_IN); 
assign P2_U7228 = ~(P2_U4944 & P2_INSTQUEUE_REG_10__5__SCAN_IN); 
assign P2_U7229 = ~(P2_U4887 & P2_INSTQUEUE_REG_11__5__SCAN_IN); 
assign P2_U7230 = ~(P2_U4829 & P2_INSTQUEUE_REG_12__5__SCAN_IN); 
assign P2_U7231 = ~(P2_U4772 & P2_INSTQUEUE_REG_13__5__SCAN_IN); 
assign P2_U7232 = ~(P2_U4713 & P2_INSTQUEUE_REG_14__5__SCAN_IN); 
assign P2_U7233 = ~(P2_U4653 & P2_INSTQUEUE_REG_15__5__SCAN_IN); 
assign P2_U7252 = ~(P2_U5517 & P2_INSTQUEUE_REG_0__4__SCAN_IN); 
assign P2_U7253 = ~(P2_U5460 & P2_INSTQUEUE_REG_1__4__SCAN_IN); 
assign P2_U7254 = ~(P2_U5402 & P2_INSTQUEUE_REG_2__4__SCAN_IN); 
assign P2_U7255 = ~(P2_U5345 & P2_INSTQUEUE_REG_3__4__SCAN_IN); 
assign P2_U7260 = ~(P2_U5059 & P2_INSTQUEUE_REG_8__4__SCAN_IN); 
assign P2_U7261 = ~(P2_U5002 & P2_INSTQUEUE_REG_9__4__SCAN_IN); 
assign P2_U7262 = ~(P2_U4944 & P2_INSTQUEUE_REG_10__4__SCAN_IN); 
assign P2_U7263 = ~(P2_U4887 & P2_INSTQUEUE_REG_11__4__SCAN_IN); 
assign P2_U7264 = ~(P2_U4829 & P2_INSTQUEUE_REG_12__4__SCAN_IN); 
assign P2_U7265 = ~(P2_U4772 & P2_INSTQUEUE_REG_13__4__SCAN_IN); 
assign P2_U7266 = ~(P2_U4713 & P2_INSTQUEUE_REG_14__4__SCAN_IN); 
assign P2_U7267 = ~(P2_U4653 & P2_INSTQUEUE_REG_15__4__SCAN_IN); 
assign P2_U7286 = ~(P2_U5517 & P2_INSTQUEUE_REG_0__3__SCAN_IN); 
assign P2_U7287 = ~(P2_U5460 & P2_INSTQUEUE_REG_1__3__SCAN_IN); 
assign P2_U7288 = ~(P2_U5402 & P2_INSTQUEUE_REG_2__3__SCAN_IN); 
assign P2_U7289 = ~(P2_U5345 & P2_INSTQUEUE_REG_3__3__SCAN_IN); 
assign P2_U7294 = ~(P2_U5059 & P2_INSTQUEUE_REG_8__3__SCAN_IN); 
assign P2_U7295 = ~(P2_U5002 & P2_INSTQUEUE_REG_9__3__SCAN_IN); 
assign P2_U7296 = ~(P2_U4944 & P2_INSTQUEUE_REG_10__3__SCAN_IN); 
assign P2_U7297 = ~(P2_U4887 & P2_INSTQUEUE_REG_11__3__SCAN_IN); 
assign P2_U7298 = ~(P2_U4829 & P2_INSTQUEUE_REG_12__3__SCAN_IN); 
assign P2_U7299 = ~(P2_U4772 & P2_INSTQUEUE_REG_13__3__SCAN_IN); 
assign P2_U7300 = ~(P2_U4713 & P2_INSTQUEUE_REG_14__3__SCAN_IN); 
assign P2_U7301 = ~(P2_U4653 & P2_INSTQUEUE_REG_15__3__SCAN_IN); 
assign P2_U7320 = ~(P2_U5517 & P2_INSTQUEUE_REG_0__2__SCAN_IN); 
assign P2_U7321 = ~(P2_U5460 & P2_INSTQUEUE_REG_1__2__SCAN_IN); 
assign P2_U7322 = ~(P2_U5402 & P2_INSTQUEUE_REG_2__2__SCAN_IN); 
assign P2_U7323 = ~(P2_U5345 & P2_INSTQUEUE_REG_3__2__SCAN_IN); 
assign P2_U7328 = ~(P2_U5059 & P2_INSTQUEUE_REG_8__2__SCAN_IN); 
assign P2_U7329 = ~(P2_U5002 & P2_INSTQUEUE_REG_9__2__SCAN_IN); 
assign P2_U7330 = ~(P2_U4944 & P2_INSTQUEUE_REG_10__2__SCAN_IN); 
assign P2_U7331 = ~(P2_U4887 & P2_INSTQUEUE_REG_11__2__SCAN_IN); 
assign P2_U7332 = ~(P2_U4829 & P2_INSTQUEUE_REG_12__2__SCAN_IN); 
assign P2_U7333 = ~(P2_U4772 & P2_INSTQUEUE_REG_13__2__SCAN_IN); 
assign P2_U7334 = ~(P2_U4713 & P2_INSTQUEUE_REG_14__2__SCAN_IN); 
assign P2_U7335 = ~(P2_U4653 & P2_INSTQUEUE_REG_15__2__SCAN_IN); 
assign P2_U7354 = ~(P2_U5517 & P2_INSTQUEUE_REG_0__1__SCAN_IN); 
assign P2_U7355 = ~(P2_U5460 & P2_INSTQUEUE_REG_1__1__SCAN_IN); 
assign P2_U7356 = ~(P2_U5402 & P2_INSTQUEUE_REG_2__1__SCAN_IN); 
assign P2_U7357 = ~(P2_U5345 & P2_INSTQUEUE_REG_3__1__SCAN_IN); 
assign P2_U7362 = ~(P2_U5059 & P2_INSTQUEUE_REG_8__1__SCAN_IN); 
assign P2_U7363 = ~(P2_U5002 & P2_INSTQUEUE_REG_9__1__SCAN_IN); 
assign P2_U7364 = ~(P2_U4944 & P2_INSTQUEUE_REG_10__1__SCAN_IN); 
assign P2_U7365 = ~(P2_U4887 & P2_INSTQUEUE_REG_11__1__SCAN_IN); 
assign P2_U7366 = ~(P2_U4829 & P2_INSTQUEUE_REG_12__1__SCAN_IN); 
assign P2_U7367 = ~(P2_U4772 & P2_INSTQUEUE_REG_13__1__SCAN_IN); 
assign P2_U7368 = ~(P2_U4713 & P2_INSTQUEUE_REG_14__1__SCAN_IN); 
assign P2_U7369 = ~(P2_U4653 & P2_INSTQUEUE_REG_15__1__SCAN_IN); 
assign P2_U7388 = ~(P2_U5517 & P2_INSTQUEUE_REG_0__0__SCAN_IN); 
assign P2_U7389 = ~(P2_U5460 & P2_INSTQUEUE_REG_1__0__SCAN_IN); 
assign P2_U7390 = ~(P2_U5402 & P2_INSTQUEUE_REG_2__0__SCAN_IN); 
assign P2_U7391 = ~(P2_U5345 & P2_INSTQUEUE_REG_3__0__SCAN_IN); 
assign P2_U7396 = ~(P2_U5059 & P2_INSTQUEUE_REG_8__0__SCAN_IN); 
assign P2_U7397 = ~(P2_U5002 & P2_INSTQUEUE_REG_9__0__SCAN_IN); 
assign P2_U7398 = ~(P2_U4944 & P2_INSTQUEUE_REG_10__0__SCAN_IN); 
assign P2_U7399 = ~(P2_U4887 & P2_INSTQUEUE_REG_11__0__SCAN_IN); 
assign P2_U7400 = ~(P2_U4829 & P2_INSTQUEUE_REG_12__0__SCAN_IN); 
assign P2_U7401 = ~(P2_U4772 & P2_INSTQUEUE_REG_13__0__SCAN_IN); 
assign P2_U7402 = ~(P2_U4713 & P2_INSTQUEUE_REG_14__0__SCAN_IN); 
assign P2_U7403 = ~(P2_U4653 & P2_INSTQUEUE_REG_15__0__SCAN_IN); 
assign P2_U8322 = ~(P2_U3242 & P2_R2267_U60); 
assign P1_U2358 = P1_U2388 & P1_U4224; 
assign P1_U2361 = P1_U4224 & P1_STATE2_REG_3__SCAN_IN; 
assign P1_U2384 = P1_U3417 & P1_STATE2_REG_0__SCAN_IN; 
assign P1_U2385 = P1_U3417 & P1_U3294; 
assign P1_U2390 = U346 & P1_U4224; 
assign P1_U2391 = U335 & P1_U4224; 
assign P1_U2392 = U324 & P1_U4224; 
assign P1_U2393 = U321 & P1_U4224; 
assign P1_U2394 = U320 & P1_U4224; 
assign P1_U2395 = U319 & P1_U4224; 
assign P1_U2396 = U318 & P1_U4224; 
assign P1_U2397 = U317 & P1_U4224; 
assign P1_U2611 = ~(P1_U6841 & P1_U6842 & P1_U6843); 
assign P1_U2801 = ~(P1_U6617 & P1_U3432 & P1_U7498); 
assign P1_U3309 = ~P1_R2144_U43; 
assign P1_U3424 = ~(P1_U4235 & P1_U6153); 
assign P1_U3587 = P1_U4552 & P1_U4553 & P1_U4224; 
assign P1_U3596 = P1_U4610 & P1_U4611 & P1_U4224; 
assign P1_U3605 = P1_U4669 & P1_U4670 & P1_U4224; 
assign P1_U3614 = P1_U4726 & P1_U4727 & P1_U4224; 
assign P1_U3623 = P1_U4784 & P1_U4785 & P1_U4224; 
assign P1_U3632 = P1_U4841 & P1_U4842 & P1_U4224; 
assign P1_U3641 = P1_U4899 & P1_U4900 & P1_U4224; 
assign P1_U3650 = P1_U4956 & P1_U4957 & P1_U4224; 
assign P1_U3659 = P1_U5012 & P1_U5013 & P1_U4224; 
assign P1_U3668 = P1_U5069 & P1_U5070 & P1_U4224; 
assign P1_U3677 = P1_U5127 & P1_U5128 & P1_U4224; 
assign P1_U3686 = P1_U5184 & P1_U5185 & P1_U4224; 
assign P1_U3695 = P1_U5242 & P1_U5243 & P1_U4224; 
assign P1_U3704 = P1_U5299 & P1_U5300 & P1_U4224; 
assign P1_U3713 = P1_U5357 & P1_U5358 & P1_U4224; 
assign P1_U3722 = P1_U5414 & P1_U5415 & P1_U4224; 
assign P1_U4172 = ~(P1_U3739 & P1_U5474); 
assign P1_U4177 = ~(P1_U2368 & P1_U3285); 
assign P1_U4222 = ~P1_U3426; 
assign P1_U4228 = ~(P1_U4235 & P1_U7500); 
assign P1_U4237 = ~P1_U4178; 
assign P1_U4502 = ~P1_U3285; 
assign P1_U5556 = ~(P1_R2144_U43 & P1_U4209); 
assign P1_U5560 = ~(P1_U2518 & P1_U5559 & P1_U7743 & P1_U7742); 
assign P1_U5799 = ~(P1_U2376 & P1_PHYADDRPOINTER_REG_0__SCAN_IN); 
assign P1_U5801 = ~(P1_U2365 & P1_REIP_REG_0__SCAN_IN); 
assign P1_U5803 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_0__SCAN_IN); 
assign P1_U5804 = ~(P1_R2337_U4 & P1_U2376); 
assign P1_U5806 = ~(P1_U2365 & P1_REIP_REG_1__SCAN_IN); 
assign P1_U5808 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_1__SCAN_IN); 
assign P1_U5809 = ~(P1_R2337_U71 & P1_U2376); 
assign P1_U5811 = ~(P1_U2365 & P1_REIP_REG_2__SCAN_IN); 
assign P1_U5813 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_2__SCAN_IN); 
assign P1_U5814 = ~(P1_R2337_U68 & P1_U2376); 
assign P1_U5816 = ~(P1_U2365 & P1_REIP_REG_3__SCAN_IN); 
assign P1_U5818 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_3__SCAN_IN); 
assign P1_U5819 = ~(P1_R2337_U67 & P1_U2376); 
assign P1_U5821 = ~(P1_U2365 & P1_REIP_REG_4__SCAN_IN); 
assign P1_U5823 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_4__SCAN_IN); 
assign P1_U5824 = ~(P1_R2337_U66 & P1_U2376); 
assign P1_U5826 = ~(P1_U2365 & P1_REIP_REG_5__SCAN_IN); 
assign P1_U5828 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_5__SCAN_IN); 
assign P1_U5829 = ~(P1_R2337_U65 & P1_U2376); 
assign P1_U5831 = ~(P1_U2365 & P1_REIP_REG_6__SCAN_IN); 
assign P1_U5833 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_6__SCAN_IN); 
assign P1_U5834 = ~(P1_R2337_U64 & P1_U2376); 
assign P1_U5836 = ~(P1_U2365 & P1_REIP_REG_7__SCAN_IN); 
assign P1_U5838 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_7__SCAN_IN); 
assign P1_U5839 = ~(P1_R2337_U63 & P1_U2376); 
assign P1_U5841 = ~(P1_U2365 & P1_REIP_REG_8__SCAN_IN); 
assign P1_U5843 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_8__SCAN_IN); 
assign P1_U5844 = ~(P1_R2337_U62 & P1_U2376); 
assign P1_U5846 = ~(P1_U2365 & P1_REIP_REG_9__SCAN_IN); 
assign P1_U5848 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_9__SCAN_IN); 
assign P1_U5849 = ~(P1_R2337_U91 & P1_U2376); 
assign P1_U5851 = ~(P1_U2365 & P1_REIP_REG_10__SCAN_IN); 
assign P1_U5853 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_10__SCAN_IN); 
assign P1_U5854 = ~(P1_R2337_U90 & P1_U2376); 
assign P1_U5856 = ~(P1_U2365 & P1_REIP_REG_11__SCAN_IN); 
assign P1_U5858 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_11__SCAN_IN); 
assign P1_U5859 = ~(P1_R2337_U89 & P1_U2376); 
assign P1_U5861 = ~(P1_U2365 & P1_REIP_REG_12__SCAN_IN); 
assign P1_U5863 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_12__SCAN_IN); 
assign P1_U5864 = ~(P1_R2337_U88 & P1_U2376); 
assign P1_U5866 = ~(P1_U2365 & P1_REIP_REG_13__SCAN_IN); 
assign P1_U5868 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_13__SCAN_IN); 
assign P1_U5869 = ~(P1_R2337_U87 & P1_U2376); 
assign P1_U5871 = ~(P1_U2365 & P1_REIP_REG_14__SCAN_IN); 
assign P1_U5873 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_14__SCAN_IN); 
assign P1_U5874 = ~(P1_R2337_U86 & P1_U2376); 
assign P1_U5876 = ~(P1_U2365 & P1_REIP_REG_15__SCAN_IN); 
assign P1_U5878 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_15__SCAN_IN); 
assign P1_U5881 = ~(P1_U2365 & P1_REIP_REG_16__SCAN_IN); 
assign P1_U5883 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_16__SCAN_IN); 
assign P1_U5886 = ~(P1_U2365 & P1_REIP_REG_17__SCAN_IN); 
assign P1_U5888 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_17__SCAN_IN); 
assign P1_U5891 = ~(P1_U2365 & P1_REIP_REG_18__SCAN_IN); 
assign P1_U5893 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_18__SCAN_IN); 
assign P1_U5896 = ~(P1_U2365 & P1_REIP_REG_19__SCAN_IN); 
assign P1_U5898 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_19__SCAN_IN); 
assign P1_U5901 = ~(P1_U2365 & P1_REIP_REG_20__SCAN_IN); 
assign P1_U5903 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_20__SCAN_IN); 
assign P1_U5906 = ~(P1_U2365 & P1_REIP_REG_21__SCAN_IN); 
assign P1_U5908 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_21__SCAN_IN); 
assign P1_U5911 = ~(P1_U2365 & P1_REIP_REG_22__SCAN_IN); 
assign P1_U5913 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_22__SCAN_IN); 
assign P1_U5916 = ~(P1_U2365 & P1_REIP_REG_23__SCAN_IN); 
assign P1_U5918 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_23__SCAN_IN); 
assign P1_U5921 = ~(P1_U2365 & P1_REIP_REG_24__SCAN_IN); 
assign P1_U5923 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_24__SCAN_IN); 
assign P1_U5926 = ~(P1_U2365 & P1_REIP_REG_25__SCAN_IN); 
assign P1_U5928 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_25__SCAN_IN); 
assign P1_U5931 = ~(P1_U2365 & P1_REIP_REG_26__SCAN_IN); 
assign P1_U5933 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_26__SCAN_IN); 
assign P1_U5936 = ~(P1_U2365 & P1_REIP_REG_27__SCAN_IN); 
assign P1_U5938 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_27__SCAN_IN); 
assign P1_U5941 = ~(P1_U2365 & P1_REIP_REG_28__SCAN_IN); 
assign P1_U5943 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_28__SCAN_IN); 
assign P1_U5946 = ~(P1_U2365 & P1_REIP_REG_29__SCAN_IN); 
assign P1_U5948 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_29__SCAN_IN); 
assign P1_U5951 = ~(P1_U2365 & P1_REIP_REG_30__SCAN_IN); 
assign P1_U5953 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_30__SCAN_IN); 
assign P1_U5956 = ~(P1_U2365 & P1_REIP_REG_31__SCAN_IN); 
assign P1_U5958 = ~(P1_U5795 & P1_PHYADDRPOINTER_REG_31__SCAN_IN); 
assign P1_U6055 = ~P1_U3417; 
assign P1_U6267 = ~(P1_U3426 & P1_EBX_REG_0__SCAN_IN); 
assign P1_U6270 = ~(P1_U3426 & P1_EBX_REG_1__SCAN_IN); 
assign P1_U6273 = ~(P1_U3426 & P1_EBX_REG_2__SCAN_IN); 
assign P1_U6276 = ~(P1_U3426 & P1_EBX_REG_3__SCAN_IN); 
assign P1_U6279 = ~(P1_U3426 & P1_EBX_REG_4__SCAN_IN); 
assign P1_U6282 = ~(P1_U3426 & P1_EBX_REG_5__SCAN_IN); 
assign P1_U6285 = ~(P1_U3426 & P1_EBX_REG_6__SCAN_IN); 
assign P1_U6288 = ~(P1_U3426 & P1_EBX_REG_7__SCAN_IN); 
assign P1_U6291 = ~(P1_U3426 & P1_EBX_REG_8__SCAN_IN); 
assign P1_U6294 = ~(P1_U3426 & P1_EBX_REG_9__SCAN_IN); 
assign P1_U6297 = ~(P1_U3426 & P1_EBX_REG_10__SCAN_IN); 
assign P1_U6300 = ~(P1_U3426 & P1_EBX_REG_11__SCAN_IN); 
assign P1_U6303 = ~(P1_U3426 & P1_EBX_REG_12__SCAN_IN); 
assign P1_U6306 = ~(P1_U3426 & P1_EBX_REG_13__SCAN_IN); 
assign P1_U6309 = ~(P1_U3426 & P1_EBX_REG_14__SCAN_IN); 
assign P1_U6312 = ~(P1_U3426 & P1_EBX_REG_15__SCAN_IN); 
assign P1_U6315 = ~(P1_U3426 & P1_EBX_REG_16__SCAN_IN); 
assign P1_U6318 = ~(P1_U3426 & P1_EBX_REG_17__SCAN_IN); 
assign P1_U6321 = ~(P1_U3426 & P1_EBX_REG_18__SCAN_IN); 
assign P1_U6324 = ~(P1_U3426 & P1_EBX_REG_19__SCAN_IN); 
assign P1_U6327 = ~(P1_U3426 & P1_EBX_REG_20__SCAN_IN); 
assign P1_U6330 = ~(P1_U3426 & P1_EBX_REG_21__SCAN_IN); 
assign P1_U6333 = ~(P1_U3426 & P1_EBX_REG_22__SCAN_IN); 
assign P1_U6336 = ~(P1_U3426 & P1_EBX_REG_23__SCAN_IN); 
assign P1_U6339 = ~(P1_U3426 & P1_EBX_REG_24__SCAN_IN); 
assign P1_U6342 = ~(P1_U3426 & P1_EBX_REG_25__SCAN_IN); 
assign P1_U6345 = ~(P1_U3426 & P1_EBX_REG_26__SCAN_IN); 
assign P1_U6348 = ~(P1_U3426 & P1_EBX_REG_27__SCAN_IN); 
assign P1_U6351 = ~(P1_U3426 & P1_EBX_REG_28__SCAN_IN); 
assign P1_U6354 = ~(P1_U3426 & P1_EBX_REG_29__SCAN_IN); 
assign P1_U6357 = ~(P1_U3426 & P1_EBX_REG_30__SCAN_IN); 
assign P1_U6359 = ~(P1_U3426 & P1_EBX_REG_31__SCAN_IN); 
assign P1_U6611 = ~(P1_U6610 & P1_CODEFETCH_REG_SCAN_IN); 
assign P1_U6889 = ~(P1_U4159 & P1_R2144_U43); 
assign P1_U7510 = ~(P1_U7493 & P1_U5962); 
assign P1_U7511 = ~(P1_U7493 & P1_U5965); 
assign P1_U7512 = ~(P1_U7493 & P1_U5968); 
assign P1_U7513 = ~(P1_U7493 & P1_U5971); 
assign P1_U7514 = ~(P1_U7493 & P1_U5974); 
assign P1_U7515 = ~(P1_U7493 & P1_U5977); 
assign P1_U7516 = ~(P1_U7493 & P1_U5980); 
assign P1_U7517 = ~(P1_U7493 & P1_U5983); 
assign P1_U7518 = ~(P1_U7493 & P1_U5986); 
assign P1_U7519 = ~(P1_U7493 & P1_U5989); 
assign P1_U7520 = ~(P1_U7493 & P1_U5992); 
assign P1_U7521 = ~(P1_U7493 & P1_U5995); 
assign P1_U7522 = ~(P1_U7493 & P1_U5998); 
assign P1_U7523 = ~(P1_U7493 & P1_U6001); 
assign P1_U7524 = ~(P1_U7493 & P1_U6004); 
assign P1_U7525 = ~(P1_U7493 & P1_U6007); 
assign P1_U7526 = ~(P1_U7493 & P1_U6010); 
assign P1_U7527 = ~(P1_U7493 & P1_U6013); 
assign P1_U7528 = ~(P1_U7493 & P1_U6016); 
assign P1_U7529 = ~(P1_U7493 & P1_U6019); 
assign P1_U7530 = ~(P1_U7493 & P1_U6022); 
assign P1_U7531 = ~(P1_U7493 & P1_U6025); 
assign P1_U7532 = ~(P1_U7493 & P1_U6028); 
assign P1_U7533 = ~(P1_U7493 & P1_U6031); 
assign P1_U7534 = ~(P1_U7493 & P1_U6034); 
assign P1_U7535 = ~(P1_U7493 & P1_U6037); 
assign P1_U7536 = ~(P1_U7493 & P1_U6040); 
assign P1_U7537 = ~(P1_U7493 & P1_U6043); 
assign P1_U7538 = ~(P1_U7493 & P1_U6046); 
assign P1_U7539 = ~(P1_U7493 & P1_U6049); 
assign P1_U7540 = ~(P1_U7493 & P1_U6052); 
assign P1_U7775 = ~(P1_U5473 & P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P1_U7776 = ~(P1_U5473 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P1_U7778 = ~(P1_U5473 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_U7780 = ~(P1_U5473 & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U7782 = ~(P1_U5473 & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P3_ADD_526_U61 = ~(P3_ADD_526_U162 & P3_ADD_526_U161); 
assign P3_ADD_526_U62 = ~(P3_ADD_526_U164 & P3_ADD_526_U163); 
assign P3_ADD_526_U128 = ~P3_ADD_526_U49; 
assign P3_ADD_526_U157 = ~(P3_ADD_526_U49 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_552_U61 = ~(P3_ADD_552_U162 & P3_ADD_552_U161); 
assign P3_ADD_552_U62 = ~(P3_ADD_552_U164 & P3_ADD_552_U163); 
assign P3_ADD_552_U128 = ~P3_ADD_552_U49; 
assign P3_ADD_552_U157 = ~(P3_ADD_552_U49 & P3_EBX_REG_30__SCAN_IN); 
assign P3_ADD_546_U61 = ~(P3_ADD_546_U162 & P3_ADD_546_U161); 
assign P3_ADD_546_U62 = ~(P3_ADD_546_U164 & P3_ADD_546_U163); 
assign P3_ADD_546_U128 = ~P3_ADD_546_U49; 
assign P3_ADD_546_U157 = ~(P3_ADD_546_U49 & P3_EAX_REG_30__SCAN_IN); 
assign P3_ADD_476_U85 = ~(P3_ADD_476_U170 & P3_ADD_476_U169); 
assign P3_ADD_476_U108 = ~P3_ADD_476_U34; 
assign P3_ADD_476_U167 = ~(P3_ADD_476_U34 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_531_U90 = ~(P3_ADD_531_U179 & P3_ADD_531_U178); 
assign P3_ADD_531_U112 = ~P3_ADD_531_U35; 
assign P3_ADD_531_U176 = ~(P3_ADD_531_U35 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_SUB_320_U119 = ~(P3_SUB_320_U95 & P3_SUB_320_U77); 
assign P3_SUB_320_U155 = ~(P3_SUB_320_U95 & P3_SUB_320_U77); 
assign P3_ADD_318_U85 = ~(P3_ADD_318_U170 & P3_ADD_318_U169); 
assign P3_ADD_318_U108 = ~P3_ADD_318_U34; 
assign P3_ADD_318_U167 = ~(P3_ADD_318_U34 & P3_PHYADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_315_U81 = ~(P3_ADD_315_U162 & P3_ADD_315_U161); 
assign P3_ADD_315_U105 = ~P3_ADD_315_U34; 
assign P3_ADD_315_U159 = ~(P3_ADD_315_U34 & P3_PHYADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_360_1242_U45 = ~(P3_ADD_360_1242_U97 & P3_ADD_360_1242_U105); 
assign P3_ADD_360_1242_U86 = ~(P3_ADD_360_1242_U201 & P3_ADD_360_1242_U200); 
assign P3_ADD_360_1242_U148 = ~P3_ADD_360_1242_U105; 
assign P3_ADD_360_1242_U185 = ~(P3_ADD_360_1242_U105 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_360_1242_U193 = ~(P3_ADD_360_1242_U105 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_LT_563_1260_U6 = P3_LT_563_1260_U7 | P3_U3304; 
assign P3_ADD_467_U85 = ~(P3_ADD_467_U170 & P3_ADD_467_U169); 
assign P3_ADD_467_U108 = ~P3_ADD_467_U34; 
assign P3_ADD_467_U167 = ~(P3_ADD_467_U34 & P3_REIP_REG_17__SCAN_IN); 
assign P3_ADD_430_U85 = ~(P3_ADD_430_U170 & P3_ADD_430_U169); 
assign P3_ADD_430_U108 = ~P3_ADD_430_U34; 
assign P3_ADD_430_U167 = ~(P3_ADD_430_U34 & P3_REIP_REG_17__SCAN_IN); 
assign P3_ADD_380_U90 = ~(P3_ADD_380_U179 & P3_ADD_380_U178); 
assign P3_ADD_380_U112 = ~P3_ADD_380_U35; 
assign P3_ADD_380_U176 = ~(P3_ADD_380_U35 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_344_U90 = ~(P3_ADD_344_U179 & P3_ADD_344_U178); 
assign P3_ADD_344_U112 = ~P3_ADD_344_U35; 
assign P3_ADD_344_U176 = ~(P3_ADD_344_U35 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_LT_563_U16 = ~P3_LT_563_U8; 
assign P3_LT_563_U19 = ~(P3_LT_563_U8 & P3_LT_563_U9); 
assign P3_ADD_339_U85 = ~(P3_ADD_339_U170 & P3_ADD_339_U169); 
assign P3_ADD_339_U108 = ~P3_ADD_339_U34; 
assign P3_ADD_339_U167 = ~(P3_ADD_339_U34 & P3_PHYADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_541_U85 = ~(P3_ADD_541_U170 & P3_ADD_541_U169); 
assign P3_ADD_541_U108 = ~P3_ADD_541_U34; 
assign P3_ADD_541_U167 = ~(P3_ADD_541_U34 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_SUB_357_1258_U68 = ~(P3_SUB_357_1258_U290 & P3_SUB_357_1258_U8); 
assign P3_SUB_357_1258_U147 = ~(P3_SUB_357_1258_U100 & P3_SUB_357_1258_U292); 
assign P3_SUB_357_1258_U149 = ~(P3_SUB_357_1258_U288 & P3_SUB_357_1258_U5); 
assign P3_SUB_357_1258_U150 = ~(P3_SUB_357_1258_U286 & P3_SUB_357_1258_U186); 
assign P3_SUB_357_1258_U312 = ~(P3_SUB_357_1258_U177 & P3_SUB_357_1258_U310); 
assign P3_ADD_515_U85 = ~(P3_ADD_515_U170 & P3_ADD_515_U169); 
assign P3_ADD_515_U108 = ~P3_ADD_515_U34; 
assign P3_ADD_515_U167 = ~(P3_ADD_515_U34 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_394_U85 = ~(P3_ADD_394_U174 & P3_ADD_394_U173); 
assign P3_ADD_394_U111 = ~P3_ADD_394_U34; 
assign P3_ADD_394_U171 = ~(P3_ADD_394_U34 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_SUB_414_U16 = P3_SUB_414_U106 & P3_SUB_414_U38; 
assign P3_SUB_414_U103 = ~P3_SUB_414_U38; 
assign P3_SUB_414_U138 = ~(P3_SUB_414_U38 & P3_EBX_REG_30__SCAN_IN); 
assign P3_ADD_441_U85 = ~(P3_ADD_441_U170 & P3_ADD_441_U169); 
assign P3_ADD_441_U108 = ~P3_ADD_441_U34; 
assign P3_ADD_441_U167 = ~(P3_ADD_441_U34 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_349_U90 = ~(P3_ADD_349_U179 & P3_ADD_349_U178); 
assign P3_ADD_349_U112 = ~P3_ADD_349_U35; 
assign P3_ADD_349_U176 = ~(P3_ADD_349_U35 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_405_U85 = ~(P3_ADD_405_U174 & P3_ADD_405_U173); 
assign P3_ADD_405_U111 = ~P3_ADD_405_U34; 
assign P3_ADD_405_U171 = ~(P3_ADD_405_U34 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_553_U90 = ~(P3_ADD_553_U179 & P3_ADD_553_U178); 
assign P3_ADD_553_U112 = ~P3_ADD_553_U35; 
assign P3_ADD_553_U176 = ~(P3_ADD_553_U35 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_558_U90 = ~(P3_ADD_558_U179 & P3_ADD_558_U178); 
assign P3_ADD_558_U112 = ~P3_ADD_558_U35; 
assign P3_ADD_558_U176 = ~(P3_ADD_558_U35 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_385_U90 = ~(P3_ADD_385_U179 & P3_ADD_385_U178); 
assign P3_ADD_385_U112 = ~P3_ADD_385_U35; 
assign P3_ADD_385_U176 = ~(P3_ADD_385_U35 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_547_U90 = ~(P3_ADD_547_U179 & P3_ADD_547_U178); 
assign P3_ADD_547_U112 = ~P3_ADD_547_U35; 
assign P3_ADD_547_U176 = ~(P3_ADD_547_U35 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_371_1212_U108 = ~(P3_ADD_371_1212_U148 & P3_ADD_371_1212_U147); 
assign P3_ADD_371_1212_U212 = ~(P3_ADD_371_1212_U145 & P3_ADD_371_1212_U210); 
assign P3_ADD_494_U85 = ~(P3_ADD_494_U170 & P3_ADD_494_U169); 
assign P3_ADD_494_U108 = ~P3_ADD_494_U34; 
assign P3_ADD_494_U167 = ~(P3_ADD_494_U34 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_536_U85 = ~(P3_ADD_536_U170 & P3_ADD_536_U169); 
assign P3_ADD_536_U108 = ~P3_ADD_536_U34; 
assign P3_ADD_536_U167 = ~(P3_ADD_536_U34 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P2_R2099_U19 = ~(P2_U2741 & P2_R2099_U121); 
assign P2_R2099_U156 = ~(P2_R2099_U121 & P2_R2099_U18); 
assign P2_ADD_391_1196_U21 = ~P2_R2182_U68; 
assign P2_ADD_391_1196_U164 = ~(P2_R2182_U68 & P2_ADD_391_1196_U163); 
assign P2_ADD_391_1196_U421 = ~(P2_R2182_U68 & P2_ADD_391_1196_U22); 
assign P2_ADD_391_1196_U425 = ~(P2_ADD_391_1196_U160 & P2_R2182_U68); 
assign P2_R2182_U128 = ~P2_R2182_U106; 
assign P2_R2182_U130 = ~(P2_R2182_U129 & P2_R2182_U106); 
assign P2_R2182_U190 = ~(P2_R2182_U99 & P2_R2182_U188); 
assign P2_R2182_U210 = ~(P2_U2678 & P2_R2182_U48); 
assign P2_R2182_U212 = ~(P2_U2678 & P2_R2182_U48); 
assign P2_R2182_U217 = ~(P2_U2658 & P2_R2182_U108); 
assign P2_R2182_U219 = ~(P2_U2658 & P2_R2182_U108); 
assign P2_R2167_U37 = ~(P2_R2167_U36 & P2_R2167_U35); 
assign P2_R2027_U90 = ~(P2_R2027_U179 & P2_R2027_U178); 
assign P2_R2027_U112 = ~P2_R2027_U35; 
assign P2_R2027_U176 = ~(P2_R2027_U35 & P2_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P2_R2337_U83 = ~(P2_R2337_U168 & P2_R2337_U167); 
assign P2_R2337_U109 = ~P2_R2337_U35; 
assign P2_R2337_U165 = ~(P2_R2337_U35 & P2_PHYADDRPOINTER_REG_18__SCAN_IN); 
assign P2_R2096_U23 = P2_U2641 & P2_R2096_U99; 
assign P2_R2096_U71 = ~(P2_R2096_U181 & P2_R2096_U180); 
assign P2_R2096_U143 = ~P2_R2096_U99; 
assign P2_R2096_U173 = ~(P2_R2096_U37 & P2_R2096_U99); 
assign P2_R1957_U119 = ~(P2_R1957_U95 & P2_R1957_U77); 
assign P2_R1957_U155 = ~(P2_R1957_U95 & P2_R1957_U77); 
assign P2_ADD_394_U91 = ~(P2_ADD_394_U186 & P2_ADD_394_U185); 
assign P2_ADD_394_U111 = ~P2_ADD_394_U34; 
assign P2_ADD_394_U135 = ~(P2_ADD_394_U34 & P2_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P2_R2267_U18 = P2_R2267_U99 & P2_R2267_U25; 
assign P2_R2267_U27 = ~P2_U3639; 
assign P2_R2267_U96 = ~(P2_R2267_U91 & P2_R2267_U57); 
assign P2_R2267_U138 = ~(P2_R2267_U91 & P2_R2267_U57); 
assign P1_R2027_U61 = ~(P1_R2027_U162 & P1_R2027_U161); 
assign P1_R2027_U62 = ~(P1_R2027_U164 & P1_R2027_U163); 
assign P1_R2027_U128 = ~P1_R2027_U49; 
assign P1_R2027_U157 = ~(P1_R2027_U49 & P1_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P1_R2144_U48 = P1_R2144_U162 & P1_R2144_U109; 
assign P1_R2144_U51 = P1_R2144_U110 & P1_R2144_U109; 
assign P1_R2144_U92 = P1_R2144_U241 & P1_R2144_U240; 
assign P1_R2144_U111 = ~(P1_U2749 & P1_R2144_U199); 
assign P1_R2144_U132 = ~(P1_R2144_U131 & P1_R2144_U93); 
assign P1_R2144_U155 = ~(P1_R2144_U154 & P1_R2144_U114); 
assign P1_R2144_U159 = ~(P1_U2749 & P1_R2144_U106 & P1_R2144_U199); 
assign P1_R2144_U161 = ~(P1_U2749 & P1_R2144_U199); 
assign P1_R2144_U163 = ~(P1_R2144_U116 & P1_R2144_U109); 
assign P1_R2144_U244 = ~(P1_R2144_U243 & P1_R2144_U242); 
assign P1_R2358_U459 = ~(P1_U2352 & P1_R2358_U158); 
assign P1_R2358_U464 = ~(P1_U2352 & P1_R2358_U158); 
assign P1_R2099_U83 = ~(P1_R2099_U340 & P1_R2099_U339); 
assign P1_R2099_U84 = ~(P1_R2099_U342 & P1_R2099_U341); 
assign P1_R2099_U164 = ~P1_R2099_U143; 
assign P1_R2099_U165 = ~P1_R2099_U12; 
assign P1_R2099_U336 = ~(P1_R2099_U58 & P1_R2099_U12); 
assign P1_R2099_U338 = ~(P1_R2099_U61 & P1_R2099_U143); 
assign P1_R2337_U85 = ~(P1_R2337_U170 & P1_R2337_U169); 
assign P1_R2337_U108 = ~P1_R2337_U34; 
assign P1_R2337_U167 = ~(P1_R2337_U34 & P1_PHYADDRPOINTER_REG_17__SCAN_IN); 
assign P1_R2096_U85 = ~(P1_R2096_U170 & P1_R2096_U169); 
assign P1_R2096_U108 = ~P1_R2096_U34; 
assign P1_R2096_U167 = ~(P1_R2096_U34 & P1_REIP_REG_17__SCAN_IN); 
assign P1_ADD_405_U91 = ~(P1_ADD_405_U186 & P1_ADD_405_U185); 
assign P1_ADD_405_U111 = ~P1_ADD_405_U34; 
assign P1_ADD_405_U135 = ~(P1_ADD_405_U34 & P1_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P1_ADD_515_U91 = ~(P1_ADD_515_U182 & P1_ADD_515_U181); 
assign P1_ADD_515_U108 = ~P1_ADD_515_U34; 
assign P1_ADD_515_U131 = ~(P1_ADD_515_U34 & P1_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_U3753 = P3_U3752 & P3_U3751 & P3_U5819; 
assign P3_U3961 = P3_U6466 & P3_U6465 & P3_U6468 & P3_U6467; 
assign P3_U4313 = ~P3_LT_563_1260_U6; 
assign P3_U5798 = ~(P3_U4318 & P3_U5796); 
assign P3_U5824 = ~(P3_ADD_360_1242_U86 & P3_U2395); 
assign P3_U5994 = ~(P3_ADD_558_U90 & P3_U3220); 
assign P3_U5995 = ~(P3_ADD_553_U90 & P3_U4298); 
assign P3_U5996 = ~(P3_ADD_547_U90 & P3_U4299); 
assign P3_U5999 = ~(P3_ADD_531_U90 & P3_U2354); 
assign P3_U6007 = ~(P3_ADD_385_U90 & P3_U2358); 
assign P3_U6008 = ~(P3_ADD_380_U90 & P3_U2359); 
assign P3_U6009 = ~(P3_ADD_349_U90 & P3_U4306); 
assign P3_U6010 = ~(P3_ADD_344_U90 & P3_U2362); 
assign P3_U6021 = ~(P3_ADD_541_U85 & P3_U4300); 
assign P3_U6022 = ~(P3_ADD_536_U85 & P3_U4301); 
assign P3_U6025 = ~(P3_ADD_515_U85 & P3_U4302); 
assign P3_U6026 = ~(P3_ADD_494_U85 & P3_U2356); 
assign P3_U6027 = ~(P3_ADD_476_U85 & P3_U4303); 
assign P3_U6028 = ~(P3_ADD_441_U85 & P3_U4304); 
assign P3_U6029 = ~(P3_ADD_405_U85 & P3_U4305); 
assign P3_U6030 = ~(P3_ADD_394_U85 & P3_U2357); 
assign P3_U6312 = ~(P3_ADD_526_U62 & P3_U2355); 
assign P3_U6336 = ~(P3_ADD_526_U61 & P3_U2355); 
assign P3_U6471 = ~(P3_U2396 & P3_ADD_360_1242_U86); 
assign P3_U6533 = ~(P3_ADD_318_U85 & P3_U2398); 
assign P3_U6538 = ~(P3_ADD_339_U85 & P3_U2388); 
assign P3_U6542 = ~(P3_ADD_315_U81 & P3_U2397); 
assign P3_U6981 = ~(P3_ADD_546_U62 & P3_U2400); 
assign P3_U6986 = ~(P3_ADD_546_U61 & P3_U2400); 
assign P3_U7083 = ~(P3_ADD_552_U62 & P3_U2399); 
assign P3_U7086 = ~(P3_ADD_552_U61 & P3_U2399); 
assign P3_U7238 = ~(P3_ADD_467_U85 & P3_U2601); 
assign P3_U7240 = ~(P3_ADD_430_U85 & P3_U2405); 
assign P3_U7341 = ~(P3_SUB_414_U16 & P3_U2602); 
assign P2_U3351 = ~(P2_R2182_U69 & P2_U3315); 
assign P2_U3893 = P2_U5658 & P2_U5659; 
assign P2_U4277 = P2_U7170 & P2_U7169 & P2_U7168 & P2_U7167; 
assign P2_U4279 = P2_U7178 & P2_U7177 & P2_U7176 & P2_U7175; 
assign P2_U4280 = P2_U7182 & P2_U7181 & P2_U7180 & P2_U7179; 
assign P2_U4281 = P2_U7187 & P2_U7186 & P2_U7185 & P2_U7184; 
assign P2_U4283 = P2_U7195 & P2_U7194 & P2_U7193 & P2_U7192; 
assign P2_U4284 = P2_U7199 & P2_U7198 & P2_U7197 & P2_U7196; 
assign P2_U4289 = P2_U7221 & P2_U7220 & P2_U7219 & P2_U7218; 
assign P2_U4291 = P2_U7229 & P2_U7228 & P2_U7227 & P2_U7226; 
assign P2_U4292 = P2_U7233 & P2_U7232 & P2_U7231 & P2_U7230; 
assign P2_U4297 = P2_U7255 & P2_U7254 & P2_U7253 & P2_U7252; 
assign P2_U4299 = P2_U7263 & P2_U7262 & P2_U7261 & P2_U7260; 
assign P2_U4300 = P2_U7267 & P2_U7266 & P2_U7265 & P2_U7264; 
assign P2_U4305 = P2_U7289 & P2_U7288 & P2_U7287 & P2_U7286; 
assign P2_U4307 = P2_U7297 & P2_U7296 & P2_U7295 & P2_U7294; 
assign P2_U4308 = P2_U7301 & P2_U7300 & P2_U7299 & P2_U7298; 
assign P2_U4313 = P2_U7323 & P2_U7322 & P2_U7321 & P2_U7320; 
assign P2_U4315 = P2_U7331 & P2_U7330 & P2_U7329 & P2_U7328; 
assign P2_U4316 = P2_U7335 & P2_U7334 & P2_U7333 & P2_U7332; 
assign P2_U4321 = P2_U7357 & P2_U7356 & P2_U7355 & P2_U7354; 
assign P2_U4323 = P2_U7365 & P2_U7364 & P2_U7363 & P2_U7362; 
assign P2_U4324 = P2_U7369 & P2_U7368 & P2_U7367 & P2_U7366; 
assign P2_U4329 = P2_U7391 & P2_U7390 & P2_U7389 & P2_U7388; 
assign P2_U4331 = P2_U7399 & P2_U7398 & P2_U7397 & P2_U7396; 
assign P2_U4332 = P2_U7403 & P2_U7402 & P2_U7401 & P2_U7400; 
assign P2_U4633 = ~P2_U3337; 
assign P2_U4637 = ~P2_U3318; 
assign P2_U4661 = ~(P2_U4654 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U4719 = ~(P2_U4714 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U4778 = ~(P2_U4773 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U4835 = ~(P2_U4830 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U4893 = ~(P2_U4888 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U4950 = ~(P2_U4945 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5008 = ~(P2_U5003 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5065 = ~(P2_U5060 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5117 = ~P2_U3430; 
assign P2_U5127 = ~(P2_U3430 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5173 = ~P2_U3441; 
assign P2_U5184 = ~(P2_U3441 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5231 = ~P2_U3453; 
assign P2_U5242 = ~(P2_U3453 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5288 = ~P2_U3464; 
assign P2_U5299 = ~(P2_U3464 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5351 = ~(P2_U5346 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5408 = ~(P2_U5403 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5466 = ~(P2_U5461 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5523 = ~(P2_U5518 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U7171 = ~(P2_U5287 & P2_INSTQUEUE_REG_4__7__SCAN_IN); 
assign P2_U7172 = ~(P2_U5230 & P2_INSTQUEUE_REG_5__7__SCAN_IN); 
assign P2_U7173 = ~(P2_U5172 & P2_INSTQUEUE_REG_6__7__SCAN_IN); 
assign P2_U7174 = ~(P2_U5116 & P2_INSTQUEUE_REG_7__7__SCAN_IN); 
assign P2_U7188 = ~(P2_U5287 & P2_INSTQUEUE_REG_4__6__SCAN_IN); 
assign P2_U7189 = ~(P2_U5230 & P2_INSTQUEUE_REG_5__6__SCAN_IN); 
assign P2_U7190 = ~(P2_U5172 & P2_INSTQUEUE_REG_6__6__SCAN_IN); 
assign P2_U7191 = ~(P2_U5116 & P2_INSTQUEUE_REG_7__6__SCAN_IN); 
assign P2_U7222 = ~(P2_U5287 & P2_INSTQUEUE_REG_4__5__SCAN_IN); 
assign P2_U7223 = ~(P2_U5230 & P2_INSTQUEUE_REG_5__5__SCAN_IN); 
assign P2_U7224 = ~(P2_U5172 & P2_INSTQUEUE_REG_6__5__SCAN_IN); 
assign P2_U7225 = ~(P2_U5116 & P2_INSTQUEUE_REG_7__5__SCAN_IN); 
assign P2_U7256 = ~(P2_U5287 & P2_INSTQUEUE_REG_4__4__SCAN_IN); 
assign P2_U7257 = ~(P2_U5230 & P2_INSTQUEUE_REG_5__4__SCAN_IN); 
assign P2_U7258 = ~(P2_U5172 & P2_INSTQUEUE_REG_6__4__SCAN_IN); 
assign P2_U7259 = ~(P2_U5116 & P2_INSTQUEUE_REG_7__4__SCAN_IN); 
assign P2_U7290 = ~(P2_U5287 & P2_INSTQUEUE_REG_4__3__SCAN_IN); 
assign P2_U7291 = ~(P2_U5230 & P2_INSTQUEUE_REG_5__3__SCAN_IN); 
assign P2_U7292 = ~(P2_U5172 & P2_INSTQUEUE_REG_6__3__SCAN_IN); 
assign P2_U7293 = ~(P2_U5116 & P2_INSTQUEUE_REG_7__3__SCAN_IN); 
assign P2_U7324 = ~(P2_U5287 & P2_INSTQUEUE_REG_4__2__SCAN_IN); 
assign P2_U7325 = ~(P2_U5230 & P2_INSTQUEUE_REG_5__2__SCAN_IN); 
assign P2_U7326 = ~(P2_U5172 & P2_INSTQUEUE_REG_6__2__SCAN_IN); 
assign P2_U7327 = ~(P2_U5116 & P2_INSTQUEUE_REG_7__2__SCAN_IN); 
assign P2_U7358 = ~(P2_U5287 & P2_INSTQUEUE_REG_4__1__SCAN_IN); 
assign P2_U7359 = ~(P2_U5230 & P2_INSTQUEUE_REG_5__1__SCAN_IN); 
assign P2_U7360 = ~(P2_U5172 & P2_INSTQUEUE_REG_6__1__SCAN_IN); 
assign P2_U7361 = ~(P2_U5116 & P2_INSTQUEUE_REG_7__1__SCAN_IN); 
assign P2_U7392 = ~(P2_U5287 & P2_INSTQUEUE_REG_4__0__SCAN_IN); 
assign P2_U7393 = ~(P2_U5230 & P2_INSTQUEUE_REG_5__0__SCAN_IN); 
assign P2_U7394 = ~(P2_U5172 & P2_INSTQUEUE_REG_6__0__SCAN_IN); 
assign P2_U7395 = ~(P2_U5116 & P2_INSTQUEUE_REG_7__0__SCAN_IN); 
assign P2_U8320 = ~(P2_U3242 & P2_R2267_U18); 
assign P2_U8403 = ~(P2_R2337_U83 & P2_U3284); 
assign P1_U2371 = P1_U4222 & P1_U4449; 
assign P1_U2383 = P1_U4222 & P1_U3391; 
assign P1_U2398 = U330 & P1_U2358; 
assign P1_U2399 = U339 & P1_U2358; 
assign P1_U2400 = U329 & P1_U2358; 
assign P1_U2401 = U338 & P1_U2358; 
assign P1_U2402 = U328 & P1_U2358; 
assign P1_U2403 = U337 & P1_U2358; 
assign P1_U2404 = U327 & P1_U2358; 
assign P1_U2405 = U336 & P1_U2358; 
assign P1_U2406 = U326 & P1_U2358; 
assign P1_U2407 = U334 & P1_U2358; 
assign P1_U2408 = U325 & P1_U2358; 
assign P1_U2409 = U333 & P1_U2358; 
assign P1_U2410 = U323 & P1_U2358; 
assign P1_U2411 = U332 & P1_U2358; 
assign P1_U2412 = U322 & P1_U2358; 
assign P1_U2413 = U331 & P1_U2358; 
assign P1_U2414 = P1_U2361 & P1_U3271; 
assign P1_U2415 = P1_U2361 & P1_U3391; 
assign P1_U2416 = P1_U2361 & P1_U3277; 
assign P1_U2417 = P1_U2361 & P1_U3284; 
assign P1_U2418 = P1_U2361 & P1_U3283; 
assign P1_U2419 = P1_U2361 & P1_U3278; 
assign P1_U2420 = P1_U2361 & P1_U4173; 
assign P1_U2421 = P1_U2361 & P1_U4171; 
assign P1_U2424 = P1_U2384 & P1_U3284; 
assign P1_U2800 = ~(P1_U6890 & P1_U6891 & P1_U6889); 
assign P1_U2803 = ~(P1_U6612 & P1_U6611); 
assign P1_U2905 = P1_U6055 & P1_DATAO_REG_31__SCAN_IN; 
assign P1_U2937 = ~(P1_U7540 & P1_U7542); 
assign P1_U2938 = ~(P1_U7539 & P1_U7544); 
assign P1_U2939 = ~(P1_U7538 & P1_U7546); 
assign P1_U2940 = ~(P1_U7537 & P1_U7548); 
assign P1_U2941 = ~(P1_U7536 & P1_U7550); 
assign P1_U2942 = ~(P1_U7535 & P1_U7552); 
assign P1_U2943 = ~(P1_U7534 & P1_U7554); 
assign P1_U2944 = ~(P1_U7533 & P1_U7556); 
assign P1_U2945 = ~(P1_U7532 & P1_U7558); 
assign P1_U2946 = ~(P1_U7531 & P1_U7560); 
assign P1_U2947 = ~(P1_U7530 & P1_U7562); 
assign P1_U2948 = ~(P1_U7529 & P1_U7564); 
assign P1_U2949 = ~(P1_U7528 & P1_U7566); 
assign P1_U2950 = ~(P1_U7527 & P1_U7568); 
assign P1_U2951 = ~(P1_U7526 & P1_U7570); 
assign P1_U2952 = ~(P1_U7525 & P1_U7572); 
assign P1_U2953 = ~(P1_U7524 & P1_U7574); 
assign P1_U2954 = ~(P1_U7523 & P1_U7576); 
assign P1_U2955 = ~(P1_U7522 & P1_U7578); 
assign P1_U2956 = ~(P1_U7521 & P1_U7580); 
assign P1_U2957 = ~(P1_U7520 & P1_U7582); 
assign P1_U2958 = ~(P1_U7519 & P1_U7584); 
assign P1_U2959 = ~(P1_U7518 & P1_U7586); 
assign P1_U2960 = ~(P1_U7517 & P1_U7588); 
assign P1_U2961 = ~(P1_U7516 & P1_U7590); 
assign P1_U2962 = ~(P1_U7515 & P1_U7592); 
assign P1_U2963 = ~(P1_U7514 & P1_U7594); 
assign P1_U2964 = ~(P1_U7513 & P1_U7596); 
assign P1_U2965 = ~(P1_U7512 & P1_U7598); 
assign P1_U2966 = ~(P1_U7511 & P1_U7600); 
assign P1_U2967 = ~(P1_U7510 & P1_U7602); 
assign P1_U3431 = ~(P1_U4228 & P1_U3887); 
assign P1_U3489 = ~(P1_U7775 & P1_U7774); 
assign P1_U3490 = ~(P1_U7777 & P1_U7776); 
assign P1_U3491 = ~(P1_U7779 & P1_U7778); 
assign P1_U3492 = ~(P1_U7781 & P1_U7780); 
assign P1_U3493 = ~(P1_U7783 & P1_U7782); 
assign P1_U4180 = ~(P1_U3967 & P1_U4228); 
assign P1_U4181 = ~(P1_U4228 & P1_U3432); 
assign P1_U4223 = ~P1_U3424; 
assign P1_U5476 = ~P1_U4172; 
assign P1_U5562 = ~(P1_U2368 & P1_U5560); 
assign P1_U5879 = ~(P1_R2337_U85 & P1_U2376); 
assign P1_U6056 = ~(P1_U2385 & P1_LWORD_REG_0__SCAN_IN); 
assign P1_U6057 = ~(P1_U2384 & P1_EAX_REG_0__SCAN_IN); 
assign P1_U6058 = ~(P1_U6055 & P1_DATAO_REG_0__SCAN_IN); 
assign P1_U6059 = ~(P1_U2385 & P1_LWORD_REG_1__SCAN_IN); 
assign P1_U6060 = ~(P1_U2384 & P1_EAX_REG_1__SCAN_IN); 
assign P1_U6061 = ~(P1_U6055 & P1_DATAO_REG_1__SCAN_IN); 
assign P1_U6062 = ~(P1_U2385 & P1_LWORD_REG_2__SCAN_IN); 
assign P1_U6063 = ~(P1_U2384 & P1_EAX_REG_2__SCAN_IN); 
assign P1_U6064 = ~(P1_U6055 & P1_DATAO_REG_2__SCAN_IN); 
assign P1_U6065 = ~(P1_U2385 & P1_LWORD_REG_3__SCAN_IN); 
assign P1_U6066 = ~(P1_U2384 & P1_EAX_REG_3__SCAN_IN); 
assign P1_U6067 = ~(P1_U6055 & P1_DATAO_REG_3__SCAN_IN); 
assign P1_U6068 = ~(P1_U2385 & P1_LWORD_REG_4__SCAN_IN); 
assign P1_U6069 = ~(P1_U2384 & P1_EAX_REG_4__SCAN_IN); 
assign P1_U6070 = ~(P1_U6055 & P1_DATAO_REG_4__SCAN_IN); 
assign P1_U6071 = ~(P1_U2385 & P1_LWORD_REG_5__SCAN_IN); 
assign P1_U6072 = ~(P1_U2384 & P1_EAX_REG_5__SCAN_IN); 
assign P1_U6073 = ~(P1_U6055 & P1_DATAO_REG_5__SCAN_IN); 
assign P1_U6074 = ~(P1_U2385 & P1_LWORD_REG_6__SCAN_IN); 
assign P1_U6075 = ~(P1_U2384 & P1_EAX_REG_6__SCAN_IN); 
assign P1_U6076 = ~(P1_U6055 & P1_DATAO_REG_6__SCAN_IN); 
assign P1_U6077 = ~(P1_U2385 & P1_LWORD_REG_7__SCAN_IN); 
assign P1_U6078 = ~(P1_U2384 & P1_EAX_REG_7__SCAN_IN); 
assign P1_U6079 = ~(P1_U6055 & P1_DATAO_REG_7__SCAN_IN); 
assign P1_U6080 = ~(P1_U2385 & P1_LWORD_REG_8__SCAN_IN); 
assign P1_U6081 = ~(P1_U2384 & P1_EAX_REG_8__SCAN_IN); 
assign P1_U6082 = ~(P1_U6055 & P1_DATAO_REG_8__SCAN_IN); 
assign P1_U6083 = ~(P1_U2385 & P1_LWORD_REG_9__SCAN_IN); 
assign P1_U6084 = ~(P1_U2384 & P1_EAX_REG_9__SCAN_IN); 
assign P1_U6085 = ~(P1_U6055 & P1_DATAO_REG_9__SCAN_IN); 
assign P1_U6086 = ~(P1_U2385 & P1_LWORD_REG_10__SCAN_IN); 
assign P1_U6087 = ~(P1_U2384 & P1_EAX_REG_10__SCAN_IN); 
assign P1_U6088 = ~(P1_U6055 & P1_DATAO_REG_10__SCAN_IN); 
assign P1_U6089 = ~(P1_U2385 & P1_LWORD_REG_11__SCAN_IN); 
assign P1_U6090 = ~(P1_U2384 & P1_EAX_REG_11__SCAN_IN); 
assign P1_U6091 = ~(P1_U6055 & P1_DATAO_REG_11__SCAN_IN); 
assign P1_U6092 = ~(P1_U2385 & P1_LWORD_REG_12__SCAN_IN); 
assign P1_U6093 = ~(P1_U2384 & P1_EAX_REG_12__SCAN_IN); 
assign P1_U6094 = ~(P1_U6055 & P1_DATAO_REG_12__SCAN_IN); 
assign P1_U6095 = ~(P1_U2385 & P1_LWORD_REG_13__SCAN_IN); 
assign P1_U6096 = ~(P1_U2384 & P1_EAX_REG_13__SCAN_IN); 
assign P1_U6097 = ~(P1_U6055 & P1_DATAO_REG_13__SCAN_IN); 
assign P1_U6098 = ~(P1_U2385 & P1_LWORD_REG_14__SCAN_IN); 
assign P1_U6099 = ~(P1_U2384 & P1_EAX_REG_14__SCAN_IN); 
assign P1_U6100 = ~(P1_U6055 & P1_DATAO_REG_14__SCAN_IN); 
assign P1_U6101 = ~(P1_U2385 & P1_LWORD_REG_15__SCAN_IN); 
assign P1_U6102 = ~(P1_U2384 & P1_EAX_REG_15__SCAN_IN); 
assign P1_U6103 = ~(P1_U6055 & P1_DATAO_REG_15__SCAN_IN); 
assign P1_U6105 = ~(P1_U2385 & P1_UWORD_REG_0__SCAN_IN); 
assign P1_U6106 = ~(P1_U6055 & P1_DATAO_REG_16__SCAN_IN); 
assign P1_U6108 = ~(P1_U2385 & P1_UWORD_REG_1__SCAN_IN); 
assign P1_U6109 = ~(P1_U6055 & P1_DATAO_REG_17__SCAN_IN); 
assign P1_U6111 = ~(P1_U2385 & P1_UWORD_REG_2__SCAN_IN); 
assign P1_U6112 = ~(P1_U6055 & P1_DATAO_REG_18__SCAN_IN); 
assign P1_U6114 = ~(P1_U2385 & P1_UWORD_REG_3__SCAN_IN); 
assign P1_U6115 = ~(P1_U6055 & P1_DATAO_REG_19__SCAN_IN); 
assign P1_U6117 = ~(P1_U2385 & P1_UWORD_REG_4__SCAN_IN); 
assign P1_U6118 = ~(P1_U6055 & P1_DATAO_REG_20__SCAN_IN); 
assign P1_U6120 = ~(P1_U2385 & P1_UWORD_REG_5__SCAN_IN); 
assign P1_U6121 = ~(P1_U6055 & P1_DATAO_REG_21__SCAN_IN); 
assign P1_U6123 = ~(P1_U2385 & P1_UWORD_REG_6__SCAN_IN); 
assign P1_U6124 = ~(P1_U6055 & P1_DATAO_REG_22__SCAN_IN); 
assign P1_U6126 = ~(P1_U2385 & P1_UWORD_REG_7__SCAN_IN); 
assign P1_U6127 = ~(P1_U6055 & P1_DATAO_REG_23__SCAN_IN); 
assign P1_U6129 = ~(P1_U2385 & P1_UWORD_REG_8__SCAN_IN); 
assign P1_U6130 = ~(P1_U6055 & P1_DATAO_REG_24__SCAN_IN); 
assign P1_U6132 = ~(P1_U2385 & P1_UWORD_REG_9__SCAN_IN); 
assign P1_U6133 = ~(P1_U6055 & P1_DATAO_REG_25__SCAN_IN); 
assign P1_U6135 = ~(P1_U2385 & P1_UWORD_REG_10__SCAN_IN); 
assign P1_U6136 = ~(P1_U6055 & P1_DATAO_REG_26__SCAN_IN); 
assign P1_U6138 = ~(P1_U2385 & P1_UWORD_REG_11__SCAN_IN); 
assign P1_U6139 = ~(P1_U6055 & P1_DATAO_REG_27__SCAN_IN); 
assign P1_U6141 = ~(P1_U2385 & P1_UWORD_REG_12__SCAN_IN); 
assign P1_U6142 = ~(P1_U6055 & P1_DATAO_REG_28__SCAN_IN); 
assign P1_U6144 = ~(P1_U2385 & P1_UWORD_REG_13__SCAN_IN); 
assign P1_U6145 = ~(P1_U6055 & P1_DATAO_REG_29__SCAN_IN); 
assign P1_U6147 = ~(P1_U2385 & P1_UWORD_REG_14__SCAN_IN); 
assign P1_U6148 = ~(P1_U6055 & P1_DATAO_REG_30__SCAN_IN); 
assign P1_U6156 = ~(P1_U3424 & P1_EAX_REG_0__SCAN_IN); 
assign P1_U6159 = ~(P1_U3424 & P1_EAX_REG_1__SCAN_IN); 
assign P1_U6162 = ~(P1_U3424 & P1_EAX_REG_2__SCAN_IN); 
assign P1_U6165 = ~(P1_U3424 & P1_EAX_REG_3__SCAN_IN); 
assign P1_U6168 = ~(P1_U3424 & P1_EAX_REG_4__SCAN_IN); 
assign P1_U6171 = ~(P1_U3424 & P1_EAX_REG_5__SCAN_IN); 
assign P1_U6174 = ~(P1_U3424 & P1_EAX_REG_6__SCAN_IN); 
assign P1_U6177 = ~(P1_U3424 & P1_EAX_REG_7__SCAN_IN); 
assign P1_U6180 = ~(P1_U3424 & P1_EAX_REG_8__SCAN_IN); 
assign P1_U6183 = ~(P1_U3424 & P1_EAX_REG_9__SCAN_IN); 
assign P1_U6186 = ~(P1_U3424 & P1_EAX_REG_10__SCAN_IN); 
assign P1_U6189 = ~(P1_U3424 & P1_EAX_REG_11__SCAN_IN); 
assign P1_U6192 = ~(P1_U3424 & P1_EAX_REG_12__SCAN_IN); 
assign P1_U6195 = ~(P1_U3424 & P1_EAX_REG_13__SCAN_IN); 
assign P1_U6198 = ~(P1_U3424 & P1_EAX_REG_14__SCAN_IN); 
assign P1_U6201 = ~(P1_U3424 & P1_EAX_REG_15__SCAN_IN); 
assign P1_U6205 = ~(P1_U3424 & P1_EAX_REG_16__SCAN_IN); 
assign P1_U6209 = ~(P1_U3424 & P1_EAX_REG_17__SCAN_IN); 
assign P1_U6213 = ~(P1_U3424 & P1_EAX_REG_18__SCAN_IN); 
assign P1_U6217 = ~(P1_U3424 & P1_EAX_REG_19__SCAN_IN); 
assign P1_U6221 = ~(P1_U3424 & P1_EAX_REG_20__SCAN_IN); 
assign P1_U6225 = ~(P1_U3424 & P1_EAX_REG_21__SCAN_IN); 
assign P1_U6229 = ~(P1_U3424 & P1_EAX_REG_22__SCAN_IN); 
assign P1_U6233 = ~(P1_U3424 & P1_EAX_REG_23__SCAN_IN); 
assign P1_U6237 = ~(P1_U3424 & P1_EAX_REG_24__SCAN_IN); 
assign P1_U6241 = ~(P1_U3424 & P1_EAX_REG_25__SCAN_IN); 
assign P1_U6245 = ~(P1_U3424 & P1_EAX_REG_26__SCAN_IN); 
assign P1_U6249 = ~(P1_U3424 & P1_EAX_REG_27__SCAN_IN); 
assign P1_U6253 = ~(P1_U3424 & P1_EAX_REG_28__SCAN_IN); 
assign P1_U6257 = ~(P1_U3424 & P1_EAX_REG_29__SCAN_IN); 
assign P1_U6261 = ~(P1_U3424 & P1_EAX_REG_30__SCAN_IN); 
assign P1_U6600 = ~P1_U4177; 
assign P1_U6601 = ~(P1_U4177 & P1_FLUSH_REG_SCAN_IN); 
assign P1_U6840 = ~(P1_R2337_U85 & P1_U2352); 
assign P1_U6870 = ~(P1_U3439 & P1_U4460 & P1_U3309); 
assign P1_U7626 = ~(P1_U4502 & P1_U4510); 
assign P1_U7701 = ~(P1_U3467 & P1_U4172); 
assign P1_U7709 = ~(P1_U5509 & P1_U4172); 
assign P1_U7722 = ~(P1_U5518 & P1_U4172); 
assign P1_U7724 = ~(P1_U5529 & P1_U4172); 
assign P1_U7728 = ~(P1_U5535 & P1_U4172); 
assign P1_U7744 = ~(P1_U3424 & P1_EAX_REG_31__SCAN_IN); 
assign P1_U7762 = ~(P1_U4177 & P1_MORE_REG_SCAN_IN); 
assign P3_ADD_526_U99 = ~(P3_ADD_526_U128 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_526_U158 = ~(P3_ADD_526_U128 & P3_ADD_526_U50); 
assign P3_ADD_552_U99 = ~(P3_ADD_552_U128 & P3_EBX_REG_30__SCAN_IN); 
assign P3_ADD_552_U158 = ~(P3_ADD_552_U128 & P3_ADD_552_U50); 
assign P3_ADD_546_U99 = ~(P3_ADD_546_U128 & P3_EAX_REG_30__SCAN_IN); 
assign P3_ADD_546_U158 = ~(P3_ADD_546_U128 & P3_ADD_546_U50); 
assign P3_ADD_476_U36 = ~(P3_ADD_476_U108 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_476_U168 = ~(P3_ADD_476_U108 & P3_ADD_476_U35); 
assign P3_ADD_531_U37 = ~(P3_ADD_531_U112 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_531_U177 = ~(P3_ADD_531_U112 & P3_ADD_531_U36); 
assign P3_SUB_320_U46 = ~P3_ADD_318_U85; 
assign P3_SUB_320_U78 = P3_SUB_320_U155 & P3_SUB_320_U154; 
assign P3_SUB_320_U120 = ~(P3_ADD_318_U85 & P3_SUB_320_U119); 
assign P3_ADD_318_U36 = ~(P3_ADD_318_U108 & P3_PHYADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_318_U168 = ~(P3_ADD_318_U108 & P3_ADD_318_U35); 
assign P3_ADD_315_U36 = ~(P3_ADD_315_U105 & P3_PHYADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_315_U160 = ~(P3_ADD_315_U105 & P3_ADD_315_U35); 
assign P3_ADD_360_1242_U119 = ~P3_ADD_360_1242_U45; 
assign P3_ADD_360_1242_U186 = ~(P3_ADD_360_1242_U42 & P3_ADD_360_1242_U185); 
assign P3_ADD_360_1242_U194 = ~(P3_ADD_360_1242_U148 & P3_ADD_360_1242_U39); 
assign P3_ADD_360_1242_U256 = ~(P3_ADD_360_1242_U45 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_467_U36 = ~(P3_ADD_467_U108 & P3_REIP_REG_17__SCAN_IN); 
assign P3_ADD_467_U168 = ~(P3_ADD_467_U108 & P3_ADD_467_U35); 
assign P3_ADD_430_U36 = ~(P3_ADD_430_U108 & P3_REIP_REG_17__SCAN_IN); 
assign P3_ADD_430_U168 = ~(P3_ADD_430_U108 & P3_ADD_430_U35); 
assign P3_ADD_380_U37 = ~(P3_ADD_380_U112 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_380_U177 = ~(P3_ADD_380_U112 & P3_ADD_380_U36); 
assign P3_ADD_344_U37 = ~(P3_ADD_344_U112 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_344_U177 = ~(P3_ADD_344_U112 & P3_ADD_344_U36); 
assign P3_LT_563_U17 = ~(P3_LT_563_U16 & P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P3_ADD_339_U36 = ~(P3_ADD_339_U108 & P3_PHYADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_339_U168 = ~(P3_ADD_339_U108 & P3_ADD_339_U35); 
assign P3_ADD_541_U36 = ~(P3_ADD_541_U108 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_541_U168 = ~(P3_ADD_541_U108 & P3_ADD_541_U35); 
assign P3_SUB_357_1258_U70 = ~(P3_SUB_357_1258_U312 & P3_SUB_357_1258_U311); 
assign P3_SUB_357_1258_U194 = ~(P3_SUB_357_1258_U193 & P3_SUB_357_1258_U147); 
assign P3_SUB_357_1258_U251 = ~(P3_SUB_357_1258_U250 & P3_SUB_357_1258_U68); 
assign P3_SUB_357_1258_U287 = ~P3_SUB_357_1258_U150; 
assign P3_SUB_357_1258_U289 = ~P3_SUB_357_1258_U149; 
assign P3_SUB_357_1258_U291 = ~P3_SUB_357_1258_U68; 
assign P3_SUB_357_1258_U293 = ~P3_SUB_357_1258_U147; 
assign P3_SUB_357_1258_U462 = ~(P3_SUB_357_1258_U146 & P3_SUB_357_1258_U147); 
assign P3_SUB_357_1258_U469 = ~(P3_SUB_357_1258_U68 & P3_SUB_357_1258_U264); 
assign P3_SUB_357_1258_U476 = ~(P3_SUB_357_1258_U148 & P3_SUB_357_1258_U149); 
assign P3_SUB_357_1258_U481 = ~(P3_SUB_357_1258_U150 & P3_SUB_357_1258_U265); 
assign P3_ADD_515_U36 = ~(P3_ADD_515_U108 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_515_U168 = ~(P3_ADD_515_U108 & P3_ADD_515_U35); 
assign P3_ADD_394_U36 = ~(P3_ADD_394_U111 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_394_U172 = ~(P3_ADD_394_U111 & P3_ADD_394_U35); 
assign P3_SUB_414_U127 = ~(P3_SUB_414_U103 & P3_SUB_414_U61); 
assign P3_SUB_414_U137 = ~(P3_SUB_414_U103 & P3_SUB_414_U61 & P3_EBX_REG_31__SCAN_IN); 
assign P3_SUB_414_U139 = ~(P3_SUB_414_U103 & P3_SUB_414_U61); 
assign P3_ADD_441_U36 = ~(P3_ADD_441_U108 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_441_U168 = ~(P3_ADD_441_U108 & P3_ADD_441_U35); 
assign P3_ADD_349_U37 = ~(P3_ADD_349_U112 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_349_U177 = ~(P3_ADD_349_U112 & P3_ADD_349_U36); 
assign P3_ADD_405_U36 = ~(P3_ADD_405_U111 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_405_U172 = ~(P3_ADD_405_U111 & P3_ADD_405_U35); 
assign P3_ADD_553_U37 = ~(P3_ADD_553_U112 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_553_U177 = ~(P3_ADD_553_U112 & P3_ADD_553_U36); 
assign P3_ADD_558_U37 = ~(P3_ADD_558_U112 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_558_U177 = ~(P3_ADD_558_U112 & P3_ADD_558_U36); 
assign P3_ADD_385_U37 = ~(P3_ADD_385_U112 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_385_U177 = ~(P3_ADD_385_U112 & P3_ADD_385_U36); 
assign P3_ADD_547_U37 = ~(P3_ADD_547_U112 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_547_U177 = ~(P3_ADD_547_U112 & P3_ADD_547_U36); 
assign P3_ADD_371_1212_U48 = ~(P3_ADD_371_1212_U99 & P3_ADD_371_1212_U108); 
assign P3_ADD_371_1212_U88 = ~(P3_ADD_371_1212_U212 & P3_ADD_371_1212_U211); 
assign P3_ADD_371_1212_U149 = ~P3_ADD_371_1212_U108; 
assign P3_ADD_371_1212_U195 = ~(P3_ADD_371_1212_U108 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_371_1212_U204 = ~(P3_ADD_371_1212_U108 & P3_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P3_ADD_494_U36 = ~(P3_ADD_494_U108 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_494_U168 = ~(P3_ADD_494_U108 & P3_ADD_494_U35); 
assign P3_ADD_536_U36 = ~(P3_ADD_536_U108 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_536_U168 = ~(P3_ADD_536_U108 & P3_ADD_536_U35); 
assign P2_R2099_U70 = ~(P2_R2099_U156 & P2_R2099_U155); 
assign P2_R2099_U122 = ~P2_R2099_U19; 
assign P2_R2099_U153 = ~(P2_U2740 & P2_R2099_U19); 
assign P2_ADD_391_1196_U14 = ~P2_R2096_U71; 
assign P2_ADD_391_1196_U123 = ~(P2_ADD_391_1196_U143 & P2_ADD_391_1196_U164); 
assign P2_ADD_391_1196_U422 = ~(P2_ADD_391_1196_U162 & P2_ADD_391_1196_U21); 
assign P2_ADD_391_1196_U424 = ~(P2_R2096_U51 & P2_ADD_391_1196_U22 & P2_ADD_391_1196_U21); 
assign P2_R2182_U40 = P2_R2182_U192 & P2_R2182_U190; 
assign P2_R2182_U97 = P2_R2182_U218 & P2_R2182_U217 & P2_R2182_U181; 
assign P2_R2182_U104 = ~(P2_R2182_U131 & P2_R2182_U130); 
assign P2_R2182_U105 = P2_R2182_U211 & P2_R2182_U210; 
assign P2_R2182_U214 = ~(P2_R2182_U213 & P2_R2182_U212); 
assign P2_R2182_U221 = ~(P2_R2182_U220 & P2_R2182_U219); 
assign P2_R2167_U38 = ~(P2_R2167_U40 & P2_R2167_U39 & P2_R2167_U37); 
assign P2_R2027_U37 = ~(P2_R2027_U112 & P2_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P2_R2027_U177 = ~(P2_R2027_U112 & P2_R2027_U36); 
assign P2_R2337_U37 = ~(P2_R2337_U109 & P2_PHYADDRPOINTER_REG_18__SCAN_IN); 
assign P2_R2337_U166 = ~(P2_R2337_U109 & P2_R2337_U36); 
assign P2_R2096_U4 = P2_U2640 & P2_R2096_U23; 
assign P2_R2096_U144 = ~P2_R2096_U23; 
assign P2_R2096_U171 = ~(P2_R2096_U28 & P2_R2096_U23); 
assign P2_R2096_U174 = ~(P2_R2096_U143 & P2_U2641); 
assign P2_R1957_U45 = ~P2_U3675; 
assign P2_R1957_U78 = P2_R1957_U155 & P2_R1957_U154; 
assign P2_R1957_U120 = ~(P2_U3675 & P2_R1957_U119); 
assign P2_ADD_394_U36 = ~(P2_ADD_394_U111 & P2_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P2_ADD_394_U136 = ~(P2_ADD_394_U111 & P2_ADD_394_U35); 
assign P2_R2267_U26 = ~(P2_R2267_U91 & P2_R2267_U57 & P2_R2267_U27); 
assign P2_R2267_U58 = P2_R2267_U138 & P2_R2267_U137; 
assign P2_R2267_U97 = ~(P2_U3639 & P2_R2267_U96); 
assign P1_R2027_U99 = ~(P1_R2027_U128 & P1_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P1_R2027_U158 = ~(P1_R2027_U128 & P1_R2027_U50); 
assign P1_R2144_U56 = P1_R2144_U159 & P1_R2144_U19; 
assign P1_R2144_U58 = P1_R2144_U19 & P1_R2144_U21 & P1_R2144_U159; 
assign P1_R2144_U62 = P1_R2144_U111 & P1_R2144_U110; 
assign P1_R2144_U91 = ~(P1_R2144_U100 & P1_R2144_U132); 
assign P1_R2144_U117 = ~(P1_R2144_U155 & P1_R2144_U157); 
assign P1_R2144_U137 = ~(P1_R2144_U161 & P1_R2144_U110); 
assign P1_R2144_U245 = ~(P1_R2144_U92 & P1_R2144_U93); 
assign P1_R2144_U246 = ~(P1_R2144_U130 & P1_R2144_U244); 
assign P1_R2358_U157 = ~P1_U2611; 
assign P1_R2358_U458 = ~(P1_U2611 & P1_R2358_U23); 
assign P1_R2358_U466 = ~(P1_R2358_U465 & P1_R2358_U464); 
assign P1_R2358_U473 = ~(P1_U2611 & P1_R2358_U23); 
assign P1_R2099_U13 = ~(P1_R2099_U94 & P1_R2099_U165); 
assign P1_R2099_U142 = ~(P1_R2099_U165 & P1_R2099_U58); 
assign P1_R2099_U335 = ~(P1_R2099_U273 & P1_R2099_U165); 
assign P1_R2099_U337 = ~(P1_R2099_U164 & P1_R2099_U270); 
assign P1_R2337_U36 = ~(P1_R2337_U108 & P1_PHYADDRPOINTER_REG_17__SCAN_IN); 
assign P1_R2337_U168 = ~(P1_R2337_U108 & P1_R2337_U35); 
assign P1_R2096_U36 = ~(P1_R2096_U108 & P1_REIP_REG_17__SCAN_IN); 
assign P1_R2096_U168 = ~(P1_R2096_U108 & P1_R2096_U35); 
assign P1_ADD_405_U36 = ~(P1_ADD_405_U111 & P1_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P1_ADD_405_U136 = ~(P1_ADD_405_U111 & P1_ADD_405_U35); 
assign P1_ADD_515_U36 = ~(P1_ADD_515_U108 & P1_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P1_ADD_515_U132 = ~(P1_ADD_515_U108 & P1_ADD_515_U35); 
assign P3_U2674 = ~(P3_U7087 & P3_U7085 & P3_U7086); 
assign P3_U2675 = ~(P3_U7084 & P3_U7082 & P3_U7083); 
assign P3_U2706 = ~(P3_U6984 & P3_U6983 & P3_U6987 & P3_U6985 & P3_U6986); 
assign P3_U2707 = ~(P3_U6979 & P3_U6978 & P3_U6982 & P3_U6980 & P3_U6981); 
assign P3_U2823 = ~(P3_U6462 & P3_U6461 & P3_U6464 & P3_U6463 & P3_U3961); 
assign P3_U2856 = ~(P3_U5799 & P3_U5797 & P3_U5798); 
assign P3_U3754 = P3_U3755 & P3_U5824; 
assign P3_U3804 = P3_U5996 & P3_U5995; 
assign P3_U3806 = P3_U5998 & P3_U5997 & P3_U5999 & P3_U3805; 
assign P3_U3809 = P3_U6010 & P3_U6009 & P3_U6008 & P3_U6007; 
assign P3_U3814 = P3_U6025 & P3_U6024; 
assign P3_U3816 = P3_U6027 & P3_U6026 & P3_U6028 & P3_U6030 & P3_U6029; 
assign P3_U4087 = P3_U7237 & P3_U4316 & P3_U7238; 
assign P3_U5820 = ~(P3_U3750 & P3_U5802 & P3_U5801 & P3_U3746 & P3_U3753); 
assign P3_U5843 = ~(P3_ADD_371_1212_U88 & P3_U2360); 
assign P3_U5849 = ~(P3_SUB_357_1258_U70 & P3_U2393); 
assign P3_U6475 = ~(P3_U2387 & P3_ADD_371_1212_U88); 
assign P3_U6480 = ~(P3_U2394 & P3_SUB_357_1258_U70); 
assign P2_U3316 = ~P2_R2182_U40; 
assign P2_U3352 = ~(P2_U3337 & P2_U3351); 
assign P2_U3674 = ~(P2_U8404 & P2_U8403); 
assign P2_U4278 = P2_U7174 & P2_U7173 & P2_U7172 & P2_U7171; 
assign P2_U4282 = P2_U7191 & P2_U7190 & P2_U7189 & P2_U7188; 
assign P2_U4290 = P2_U7225 & P2_U7224 & P2_U7223 & P2_U7222; 
assign P2_U4298 = P2_U7259 & P2_U7258 & P2_U7257 & P2_U7256; 
assign P2_U4306 = P2_U7293 & P2_U7292 & P2_U7291 & P2_U7290; 
assign P2_U4314 = P2_U7327 & P2_U7326 & P2_U7325 & P2_U7324; 
assign P2_U4322 = P2_U7361 & P2_U7360 & P2_U7359 & P2_U7358; 
assign P2_U4330 = P2_U7395 & P2_U7394 & P2_U7393 & P2_U7392; 
assign P2_U4634 = ~P2_U3351; 
assign P2_U5121 = ~(P2_U5117 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5178 = ~(P2_U5173 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5236 = ~(P2_U5231 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5293 = ~(P2_U5288 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U5653 = ~(P2_R2182_U40 & P2_U5644); 
assign P2_U8062 = ~(P2_R2182_U40 & P2_U3318); 
assign P2_U8318 = ~(P2_U3242 & P2_R2267_U58); 
assign P1_U2359 = P1_U3431 & P1_STATE2_REG_2__SCAN_IN; 
assign P1_U2373 = P1_U3431 & P1_STATE2_REG_3__SCAN_IN; 
assign P1_U2386 = P1_U4223 & P1_U3423; 
assign P1_U2387 = P1_U3884 & P1_U4223; 
assign P1_U2422 = P1_U4223 & P1_U5461; 
assign P1_U2423 = P1_U4223 & P1_U4231; 
assign P1_U2426 = P1_U3889 & P1_U3431; 
assign P1_U2650 = P1_U6870 & P1_STATE2_REG_2__SCAN_IN; 
assign P1_U2806 = ~(P1_U6601 & P1_U4248); 
assign P1_U2921 = ~(P1_U6102 & P1_U6101 & P1_U6103); 
assign P1_U2922 = ~(P1_U6099 & P1_U6098 & P1_U6100); 
assign P1_U2923 = ~(P1_U6096 & P1_U6095 & P1_U6097); 
assign P1_U2924 = ~(P1_U6093 & P1_U6092 & P1_U6094); 
assign P1_U2925 = ~(P1_U6090 & P1_U6089 & P1_U6091); 
assign P1_U2926 = ~(P1_U6087 & P1_U6086 & P1_U6088); 
assign P1_U2927 = ~(P1_U6084 & P1_U6083 & P1_U6085); 
assign P1_U2928 = ~(P1_U6081 & P1_U6080 & P1_U6082); 
assign P1_U2929 = ~(P1_U6078 & P1_U6077 & P1_U6079); 
assign P1_U2930 = ~(P1_U6075 & P1_U6074 & P1_U6076); 
assign P1_U2931 = ~(P1_U6072 & P1_U6071 & P1_U6073); 
assign P1_U2932 = ~(P1_U6069 & P1_U6068 & P1_U6070); 
assign P1_U2933 = ~(P1_U6066 & P1_U6065 & P1_U6067); 
assign P1_U2934 = ~(P1_U6063 & P1_U6062 & P1_U6064); 
assign P1_U2935 = ~(P1_U6060 & P1_U6059 & P1_U6061); 
assign P1_U2936 = ~(P1_U6057 & P1_U6056 & P1_U6058); 
assign P1_U3414 = ~(P1_U3756 & P1_U5562); 
assign P1_U3868 = P1_U6105 & P1_U6106; 
assign P1_U3869 = P1_U6108 & P1_U6109; 
assign P1_U3870 = P1_U6111 & P1_U6112; 
assign P1_U3871 = P1_U6114 & P1_U6115; 
assign P1_U3872 = P1_U6117 & P1_U6118; 
assign P1_U3873 = P1_U6120 & P1_U6121; 
assign P1_U3874 = P1_U6123 & P1_U6124; 
assign P1_U3875 = P1_U6126 & P1_U6127; 
assign P1_U3876 = P1_U6129 & P1_U6130; 
assign P1_U3877 = P1_U6132 & P1_U6133; 
assign P1_U3878 = P1_U6135 & P1_U6136; 
assign P1_U3879 = P1_U6138 & P1_U6139; 
assign P1_U3880 = P1_U6141 & P1_U6142; 
assign P1_U3881 = P1_U6144 & P1_U6145; 
assign P1_U3882 = P1_U6147 & P1_U6148; 
assign P1_U4025 = P1_U6838 & P1_U6839 & P1_U6840; 
assign P1_U4227 = ~(P1_U4255 & P1_U3431); 
assign P1_U4560 = ~(P1_U2415 & P1_U4534); 
assign P1_U4565 = ~(P1_U2416 & P1_U4534); 
assign P1_U4570 = ~(P1_U2420 & P1_U4534); 
assign P1_U4575 = ~(P1_U2419 & P1_U4534); 
assign P1_U4580 = ~(P1_U2418 & P1_U4534); 
assign P1_U4585 = ~(P1_U2421 & P1_U4534); 
assign P1_U4590 = ~(P1_U2414 & P1_U4534); 
assign P1_U4595 = ~(P1_U2417 & P1_U4534); 
assign P1_U4618 = ~(P1_U4602 & P1_U2415); 
assign P1_U4623 = ~(P1_U4602 & P1_U2416); 
assign P1_U4628 = ~(P1_U4602 & P1_U2420); 
assign P1_U4633 = ~(P1_U4602 & P1_U2419); 
assign P1_U4638 = ~(P1_U4602 & P1_U2418); 
assign P1_U4643 = ~(P1_U4602 & P1_U2421); 
assign P1_U4648 = ~(P1_U4602 & P1_U2414); 
assign P1_U4653 = ~(P1_U4602 & P1_U2417); 
assign P1_U4677 = ~(P1_U4660 & P1_U2415); 
assign P1_U4682 = ~(P1_U4660 & P1_U2416); 
assign P1_U4687 = ~(P1_U4660 & P1_U2420); 
assign P1_U4692 = ~(P1_U4660 & P1_U2419); 
assign P1_U4697 = ~(P1_U4660 & P1_U2418); 
assign P1_U4702 = ~(P1_U4660 & P1_U2421); 
assign P1_U4707 = ~(P1_U4660 & P1_U2414); 
assign P1_U4712 = ~(P1_U4660 & P1_U2417); 
assign P1_U4734 = ~(P1_U4718 & P1_U2415); 
assign P1_U4739 = ~(P1_U4718 & P1_U2416); 
assign P1_U4744 = ~(P1_U4718 & P1_U2420); 
assign P1_U4749 = ~(P1_U4718 & P1_U2419); 
assign P1_U4754 = ~(P1_U4718 & P1_U2418); 
assign P1_U4759 = ~(P1_U4718 & P1_U2421); 
assign P1_U4764 = ~(P1_U4718 & P1_U2414); 
assign P1_U4769 = ~(P1_U4718 & P1_U2417); 
assign P1_U4792 = ~(P1_U4775 & P1_U2415); 
assign P1_U4797 = ~(P1_U4775 & P1_U2416); 
assign P1_U4802 = ~(P1_U4775 & P1_U2420); 
assign P1_U4807 = ~(P1_U4775 & P1_U2419); 
assign P1_U4812 = ~(P1_U4775 & P1_U2418); 
assign P1_U4817 = ~(P1_U4775 & P1_U2421); 
assign P1_U4822 = ~(P1_U4775 & P1_U2414); 
assign P1_U4827 = ~(P1_U4775 & P1_U2417); 
assign P1_U4849 = ~(P1_U4833 & P1_U2415); 
assign P1_U4854 = ~(P1_U4833 & P1_U2416); 
assign P1_U4859 = ~(P1_U4833 & P1_U2420); 
assign P1_U4864 = ~(P1_U4833 & P1_U2419); 
assign P1_U4869 = ~(P1_U4833 & P1_U2418); 
assign P1_U4874 = ~(P1_U4833 & P1_U2421); 
assign P1_U4879 = ~(P1_U4833 & P1_U2414); 
assign P1_U4884 = ~(P1_U4833 & P1_U2417); 
assign P1_U4907 = ~(P1_U4890 & P1_U2415); 
assign P1_U4912 = ~(P1_U4890 & P1_U2416); 
assign P1_U4917 = ~(P1_U4890 & P1_U2420); 
assign P1_U4922 = ~(P1_U4890 & P1_U2419); 
assign P1_U4927 = ~(P1_U4890 & P1_U2418); 
assign P1_U4932 = ~(P1_U4890 & P1_U2421); 
assign P1_U4937 = ~(P1_U4890 & P1_U2414); 
assign P1_U4942 = ~(P1_U4890 & P1_U2417); 
assign P1_U4964 = ~(P1_U4948 & P1_U2415); 
assign P1_U4969 = ~(P1_U4948 & P1_U2416); 
assign P1_U4974 = ~(P1_U4948 & P1_U2420); 
assign P1_U4979 = ~(P1_U4948 & P1_U2419); 
assign P1_U4984 = ~(P1_U4948 & P1_U2418); 
assign P1_U4989 = ~(P1_U4948 & P1_U2421); 
assign P1_U4994 = ~(P1_U4948 & P1_U2414); 
assign P1_U4999 = ~(P1_U4948 & P1_U2417); 
assign P1_U5020 = ~(P1_U4537 & P1_U2415); 
assign P1_U5025 = ~(P1_U4537 & P1_U2416); 
assign P1_U5030 = ~(P1_U4537 & P1_U2420); 
assign P1_U5035 = ~(P1_U4537 & P1_U2419); 
assign P1_U5040 = ~(P1_U4537 & P1_U2418); 
assign P1_U5045 = ~(P1_U4537 & P1_U2421); 
assign P1_U5050 = ~(P1_U4537 & P1_U2414); 
assign P1_U5055 = ~(P1_U4537 & P1_U2417); 
assign P1_U5077 = ~(P1_U5061 & P1_U2415); 
assign P1_U5082 = ~(P1_U5061 & P1_U2416); 
assign P1_U5087 = ~(P1_U5061 & P1_U2420); 
assign P1_U5092 = ~(P1_U5061 & P1_U2419); 
assign P1_U5097 = ~(P1_U5061 & P1_U2418); 
assign P1_U5102 = ~(P1_U5061 & P1_U2421); 
assign P1_U5107 = ~(P1_U5061 & P1_U2414); 
assign P1_U5112 = ~(P1_U5061 & P1_U2417); 
assign P1_U5135 = ~(P1_U5118 & P1_U2415); 
assign P1_U5140 = ~(P1_U5118 & P1_U2416); 
assign P1_U5145 = ~(P1_U5118 & P1_U2420); 
assign P1_U5150 = ~(P1_U5118 & P1_U2419); 
assign P1_U5155 = ~(P1_U5118 & P1_U2418); 
assign P1_U5160 = ~(P1_U5118 & P1_U2421); 
assign P1_U5165 = ~(P1_U5118 & P1_U2414); 
assign P1_U5170 = ~(P1_U5118 & P1_U2417); 
assign P1_U5192 = ~(P1_U5176 & P1_U2415); 
assign P1_U5197 = ~(P1_U5176 & P1_U2416); 
assign P1_U5202 = ~(P1_U5176 & P1_U2420); 
assign P1_U5207 = ~(P1_U5176 & P1_U2419); 
assign P1_U5212 = ~(P1_U5176 & P1_U2418); 
assign P1_U5217 = ~(P1_U5176 & P1_U2421); 
assign P1_U5222 = ~(P1_U5176 & P1_U2414); 
assign P1_U5227 = ~(P1_U5176 & P1_U2417); 
assign P1_U5250 = ~(P1_U5233 & P1_U2415); 
assign P1_U5255 = ~(P1_U5233 & P1_U2416); 
assign P1_U5260 = ~(P1_U5233 & P1_U2420); 
assign P1_U5265 = ~(P1_U5233 & P1_U2419); 
assign P1_U5270 = ~(P1_U5233 & P1_U2418); 
assign P1_U5275 = ~(P1_U5233 & P1_U2421); 
assign P1_U5280 = ~(P1_U5233 & P1_U2414); 
assign P1_U5285 = ~(P1_U5233 & P1_U2417); 
assign P1_U5307 = ~(P1_U5291 & P1_U2415); 
assign P1_U5312 = ~(P1_U5291 & P1_U2416); 
assign P1_U5317 = ~(P1_U5291 & P1_U2420); 
assign P1_U5322 = ~(P1_U5291 & P1_U2419); 
assign P1_U5327 = ~(P1_U5291 & P1_U2418); 
assign P1_U5332 = ~(P1_U5291 & P1_U2421); 
assign P1_U5337 = ~(P1_U5291 & P1_U2414); 
assign P1_U5342 = ~(P1_U5291 & P1_U2417); 
assign P1_U5365 = ~(P1_U5348 & P1_U2415); 
assign P1_U5370 = ~(P1_U5348 & P1_U2416); 
assign P1_U5375 = ~(P1_U5348 & P1_U2420); 
assign P1_U5380 = ~(P1_U5348 & P1_U2419); 
assign P1_U5385 = ~(P1_U5348 & P1_U2418); 
assign P1_U5390 = ~(P1_U5348 & P1_U2421); 
assign P1_U5395 = ~(P1_U5348 & P1_U2414); 
assign P1_U5400 = ~(P1_U5348 & P1_U2417); 
assign P1_U5422 = ~(P1_U5406 & P1_U2415); 
assign P1_U5427 = ~(P1_U5406 & P1_U2416); 
assign P1_U5432 = ~(P1_U5406 & P1_U2420); 
assign P1_U5437 = ~(P1_U5406 & P1_U2419); 
assign P1_U5441 = ~(P1_U5406 & P1_U2418); 
assign P1_U5446 = ~(P1_U5406 & P1_U2421); 
assign P1_U5451 = ~(P1_U5406 & P1_U2414); 
assign P1_U5456 = ~(P1_U5406 & P1_U2417); 
assign P1_U6104 = ~(P1_U2424 & P1_EAX_REG_16__SCAN_IN); 
assign P1_U6107 = ~(P1_U2424 & P1_EAX_REG_17__SCAN_IN); 
assign P1_U6110 = ~(P1_U2424 & P1_EAX_REG_18__SCAN_IN); 
assign P1_U6113 = ~(P1_U2424 & P1_EAX_REG_19__SCAN_IN); 
assign P1_U6116 = ~(P1_U2424 & P1_EAX_REG_20__SCAN_IN); 
assign P1_U6119 = ~(P1_U2424 & P1_EAX_REG_21__SCAN_IN); 
assign P1_U6122 = ~(P1_U2424 & P1_EAX_REG_22__SCAN_IN); 
assign P1_U6125 = ~(P1_U2424 & P1_EAX_REG_23__SCAN_IN); 
assign P1_U6128 = ~(P1_U2424 & P1_EAX_REG_24__SCAN_IN); 
assign P1_U6131 = ~(P1_U2424 & P1_EAX_REG_25__SCAN_IN); 
assign P1_U6134 = ~(P1_U2424 & P1_EAX_REG_26__SCAN_IN); 
assign P1_U6137 = ~(P1_U2424 & P1_EAX_REG_27__SCAN_IN); 
assign P1_U6140 = ~(P1_U2424 & P1_EAX_REG_28__SCAN_IN); 
assign P1_U6143 = ~(P1_U2424 & P1_EAX_REG_29__SCAN_IN); 
assign P1_U6146 = ~(P1_U2424 & P1_EAX_REG_30__SCAN_IN); 
assign P1_U6266 = ~(P1_U2371 & P1_R2099_U86); 
assign P1_U6269 = ~(P1_U2371 & P1_R2099_U87); 
assign P1_U6272 = ~(P1_U2371 & P1_R2099_U138); 
assign P1_U6275 = ~(P1_U2371 & P1_R2099_U42); 
assign P1_U6278 = ~(P1_U2371 & P1_R2099_U41); 
assign P1_U6281 = ~(P1_U2371 & P1_R2099_U40); 
assign P1_U6284 = ~(P1_U2371 & P1_R2099_U39); 
assign P1_U6287 = ~(P1_U2371 & P1_R2099_U38); 
assign P1_U6290 = ~(P1_U2371 & P1_R2099_U37); 
assign P1_U6293 = ~(P1_U2371 & P1_R2099_U36); 
assign P1_U6296 = ~(P1_U2371 & P1_R2099_U85); 
assign P1_U6299 = ~(P1_U2371 & P1_R2099_U84); 
assign P1_U6302 = ~(P1_U2371 & P1_R2099_U83); 
assign P1_U6363 = ~P1_U3431; 
assign P1_U6603 = ~P1_U4180; 
assign P1_U6614 = ~P1_U4181; 
assign P1_U7458 = ~(P1_U3489 & P1_U3262); 
assign P1_U7460 = ~(P1_U3490 & P1_U3262); 
assign P1_U7463 = ~(P1_U3491 & P1_U3262); 
assign P1_U7466 = ~(P1_U3492 & P1_U3262); 
assign P1_U7702 = ~(P1_U5476 & P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P1_U7708 = ~(P1_U5476 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P1_U7721 = ~(P1_U5476 & P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P1_U7723 = ~(P1_U5476 & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P1_U7727 = ~(P1_U5476 & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U7763 = ~(P1_U4237 & P1_U6600); 
assign P1_U7767 = ~(P1_U6609 & P1_U4180); 
assign P1_U7773 = ~(P1_U6615 & P1_U4181); 
assign P1_U7793 = ~(P1_U3493 & P1_U3262); 
assign P3_ADD_526_U59 = ~(P3_ADD_526_U158 & P3_ADD_526_U157); 
assign P3_ADD_526_U129 = ~P3_ADD_526_U99; 
assign P3_ADD_526_U155 = ~(P3_ADD_526_U99 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_552_U59 = ~(P3_ADD_552_U158 & P3_ADD_552_U157); 
assign P3_ADD_552_U129 = ~P3_ADD_552_U99; 
assign P3_ADD_552_U155 = ~(P3_ADD_552_U99 & P3_EBX_REG_31__SCAN_IN); 
assign P3_ADD_546_U59 = ~(P3_ADD_546_U158 & P3_ADD_546_U157); 
assign P3_ADD_546_U129 = ~P3_ADD_546_U99; 
assign P3_ADD_546_U155 = ~(P3_ADD_546_U99 & P3_EAX_REG_31__SCAN_IN); 
assign P3_ADD_476_U84 = ~(P3_ADD_476_U168 & P3_ADD_476_U167); 
assign P3_ADD_476_U109 = ~P3_ADD_476_U36; 
assign P3_ADD_476_U165 = ~(P3_ADD_476_U36 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_531_U89 = ~(P3_ADD_531_U177 & P3_ADD_531_U176); 
assign P3_ADD_531_U113 = ~P3_ADD_531_U37; 
assign P3_ADD_531_U174 = ~(P3_ADD_531_U37 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_SUB_320_U31 = ~(P3_SUB_320_U46 & P3_SUB_320_U77 & P3_SUB_320_U95); 
assign P3_ADD_318_U84 = ~(P3_ADD_318_U168 & P3_ADD_318_U167); 
assign P3_ADD_318_U109 = ~P3_ADD_318_U36; 
assign P3_ADD_318_U165 = ~(P3_ADD_318_U36 & P3_PHYADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_315_U80 = ~(P3_ADD_315_U160 & P3_ADD_315_U159); 
assign P3_ADD_315_U106 = ~P3_ADD_315_U36; 
assign P3_ADD_315_U157 = ~(P3_ADD_315_U36 & P3_PHYADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_360_1242_U4 = P3_ADD_360_1242_U186 & P3_ADD_360_1242_U45; 
assign P3_ADD_360_1242_U46 = ~(P3_ADD_360_1242_U98 & P3_ADD_360_1242_U119); 
assign P3_ADD_360_1242_U106 = P3_ADD_360_1242_U194 & P3_ADD_360_1242_U193; 
assign P3_ADD_360_1242_U183 = ~(P3_ADD_360_1242_U119 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_360_1242_U255 = ~(P3_ADD_360_1242_U119 & P3_ADD_360_1242_U43); 
assign P3_ADD_467_U84 = ~(P3_ADD_467_U168 & P3_ADD_467_U167); 
assign P3_ADD_467_U109 = ~P3_ADD_467_U36; 
assign P3_ADD_467_U165 = ~(P3_ADD_467_U36 & P3_REIP_REG_18__SCAN_IN); 
assign P3_ADD_430_U84 = ~(P3_ADD_430_U168 & P3_ADD_430_U167); 
assign P3_ADD_430_U109 = ~P3_ADD_430_U36; 
assign P3_ADD_430_U165 = ~(P3_ADD_430_U36 & P3_REIP_REG_18__SCAN_IN); 
assign P3_ADD_380_U89 = ~(P3_ADD_380_U177 & P3_ADD_380_U176); 
assign P3_ADD_380_U113 = ~P3_ADD_380_U37; 
assign P3_ADD_380_U174 = ~(P3_ADD_380_U37 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_344_U89 = ~(P3_ADD_344_U177 & P3_ADD_344_U176); 
assign P3_ADD_344_U113 = ~P3_ADD_344_U37; 
assign P3_ADD_344_U174 = ~(P3_ADD_344_U37 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_LT_563_U18 = ~(P3_U3307 & P3_LT_563_U17); 
assign P3_ADD_339_U84 = ~(P3_ADD_339_U168 & P3_ADD_339_U167); 
assign P3_ADD_339_U109 = ~P3_ADD_339_U36; 
assign P3_ADD_339_U165 = ~(P3_ADD_339_U36 & P3_PHYADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_541_U84 = ~(P3_ADD_541_U168 & P3_ADD_541_U167); 
assign P3_ADD_541_U109 = ~P3_ADD_541_U36; 
assign P3_ADD_541_U165 = ~(P3_ADD_541_U36 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_SUB_357_1258_U145 = ~(P3_SUB_357_1258_U195 & P3_SUB_357_1258_U194); 
assign P3_SUB_357_1258_U252 = ~(P3_SUB_357_1258_U113 & P3_SUB_357_1258_U251); 
assign P3_SUB_357_1258_U253 = ~(P3_SUB_357_1258_U291 & P3_SUB_357_1258_U155); 
assign P3_SUB_357_1258_U463 = ~(P3_SUB_357_1258_U293 & P3_SUB_357_1258_U461); 
assign P3_SUB_357_1258_U470 = ~(P3_SUB_357_1258_U468 & P3_SUB_357_1258_U291); 
assign P3_SUB_357_1258_U477 = ~(P3_SUB_357_1258_U289 & P3_SUB_357_1258_U475); 
assign P3_SUB_357_1258_U482 = ~(P3_SUB_357_1258_U287 & P3_SUB_357_1258_U480); 
assign P3_ADD_515_U84 = ~(P3_ADD_515_U168 & P3_ADD_515_U167); 
assign P3_ADD_515_U109 = ~P3_ADD_515_U36; 
assign P3_ADD_515_U165 = ~(P3_ADD_515_U36 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_394_U84 = ~(P3_ADD_394_U172 & P3_ADD_394_U171); 
assign P3_ADD_394_U112 = ~P3_ADD_394_U36; 
assign P3_ADD_394_U169 = ~(P3_ADD_394_U36 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_SUB_414_U62 = P3_SUB_414_U139 & P3_SUB_414_U138; 
assign P3_SUB_414_U136 = ~(P3_SUB_414_U127 & P3_SUB_414_U60); 
assign P3_ADD_441_U84 = ~(P3_ADD_441_U168 & P3_ADD_441_U167); 
assign P3_ADD_441_U109 = ~P3_ADD_441_U36; 
assign P3_ADD_441_U165 = ~(P3_ADD_441_U36 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_349_U89 = ~(P3_ADD_349_U177 & P3_ADD_349_U176); 
assign P3_ADD_349_U113 = ~P3_ADD_349_U37; 
assign P3_ADD_349_U174 = ~(P3_ADD_349_U37 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_405_U84 = ~(P3_ADD_405_U172 & P3_ADD_405_U171); 
assign P3_ADD_405_U112 = ~P3_ADD_405_U36; 
assign P3_ADD_405_U169 = ~(P3_ADD_405_U36 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_553_U89 = ~(P3_ADD_553_U177 & P3_ADD_553_U176); 
assign P3_ADD_553_U113 = ~P3_ADD_553_U37; 
assign P3_ADD_553_U174 = ~(P3_ADD_553_U37 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_558_U89 = ~(P3_ADD_558_U177 & P3_ADD_558_U176); 
assign P3_ADD_558_U113 = ~P3_ADD_558_U37; 
assign P3_ADD_558_U174 = ~(P3_ADD_558_U37 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_385_U89 = ~(P3_ADD_385_U177 & P3_ADD_385_U176); 
assign P3_ADD_385_U113 = ~P3_ADD_385_U37; 
assign P3_ADD_385_U174 = ~(P3_ADD_385_U37 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_547_U89 = ~(P3_ADD_547_U177 & P3_ADD_547_U176); 
assign P3_ADD_547_U113 = ~P3_ADD_547_U37; 
assign P3_ADD_547_U174 = ~(P3_ADD_547_U37 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_371_1212_U117 = ~P3_ADD_371_1212_U48; 
assign P3_ADD_371_1212_U196 = ~(P3_ADD_371_1212_U45 & P3_ADD_371_1212_U195); 
assign P3_ADD_371_1212_U205 = ~(P3_ADD_371_1212_U149 & P3_ADD_371_1212_U42); 
assign P3_ADD_371_1212_U263 = ~(P3_ADD_371_1212_U48 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_494_U84 = ~(P3_ADD_494_U168 & P3_ADD_494_U167); 
assign P3_ADD_494_U109 = ~P3_ADD_494_U36; 
assign P3_ADD_494_U165 = ~(P3_ADD_494_U36 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_536_U84 = ~(P3_ADD_536_U168 & P3_ADD_536_U167); 
assign P3_ADD_536_U109 = ~P3_ADD_536_U36; 
assign P3_ADD_536_U165 = ~(P3_ADD_536_U36 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P2_R2099_U21 = ~(P2_U2740 & P2_R2099_U122); 
assign P2_R2099_U154 = ~(P2_R2099_U122 & P2_R2099_U20); 
assign P2_ADD_391_1196_U24 = ~P2_R2182_U40; 
assign P2_ADD_391_1196_U144 = P2_ADD_391_1196_U425 & P2_ADD_391_1196_U424; 
assign P2_ADD_391_1196_U165 = ~P2_ADD_391_1196_U123; 
assign P2_ADD_391_1196_U166 = P2_R2182_U40 | P2_R2096_U77; 
assign P2_ADD_391_1196_U168 = ~(P2_R2096_U77 & P2_R2182_U40); 
assign P2_ADD_391_1196_U345 = ~(P2_R2182_U40 & P2_ADD_391_1196_U25); 
assign P2_ADD_391_1196_U347 = ~(P2_R2182_U40 & P2_ADD_391_1196_U25); 
assign P2_ADD_391_1196_U423 = ~(P2_ADD_391_1196_U422 & P2_ADD_391_1196_U421); 
assign P2_R2182_U98 = P2_R2182_U185 & P2_R2182_U221; 
assign P2_R2182_U132 = ~P2_R2182_U104; 
assign P2_R2182_U134 = ~(P2_R2182_U133 & P2_R2182_U104); 
assign P2_R2182_U208 = ~(P2_R2182_U103 & P2_R2182_U104); 
assign P2_R2182_U215 = ~(P2_R2182_U105 & P2_R2182_U106); 
assign P2_R2182_U216 = ~(P2_R2182_U128 & P2_R2182_U214); 
assign P2_R2167_U6 = ~(P2_R2167_U42 & P2_R2167_U41 & P2_R2167_U38); 
assign P2_R2027_U89 = ~(P2_R2027_U177 & P2_R2027_U176); 
assign P2_R2027_U113 = ~P2_R2027_U37; 
assign P2_R2027_U174 = ~(P2_R2027_U37 & P2_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P2_R2337_U82 = ~(P2_R2337_U166 & P2_R2337_U165); 
assign P2_R2337_U110 = ~P2_R2337_U37; 
assign P2_R2337_U163 = ~(P2_R2337_U37 & P2_PHYADDRPOINTER_REG_19__SCAN_IN); 
assign P2_R2096_U24 = P2_U2639 & P2_R2096_U4; 
assign P2_R2096_U70 = ~(P2_R2096_U174 & P2_R2096_U173); 
assign P2_R2096_U145 = ~P2_R2096_U4; 
assign P2_R2096_U172 = ~(P2_R2096_U144 & P2_U2640); 
assign P2_R2096_U262 = ~(P2_R2096_U49 & P2_R2096_U4); 
assign P2_R1957_U30 = ~(P2_R1957_U95 & P2_R1957_U77 & P2_R1957_U45); 
assign P2_ADD_394_U67 = ~(P2_ADD_394_U136 & P2_ADD_394_U135); 
assign P2_ADD_394_U112 = ~P2_ADD_394_U36; 
assign P2_ADD_394_U145 = ~(P2_ADD_394_U36 & P2_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P2_R2267_U19 = P2_R2267_U97 & P2_R2267_U26; 
assign P2_R2267_U92 = ~P2_R2267_U26; 
assign P2_R2267_U135 = ~(P2_U2789 & P2_R2267_U26); 
assign P1_R2027_U59 = ~(P1_R2027_U158 & P1_R2027_U157); 
assign P1_R2027_U129 = ~P1_R2027_U99; 
assign P1_R2027_U155 = ~(P1_R2027_U99 & P1_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P1_R2144_U50 = ~(P1_R2144_U246 & P1_R2144_U245); 
assign P1_R2144_U118 = ~(P1_R2144_U51 & P1_R2144_U117); 
assign P1_R2144_U133 = ~P1_R2144_U91; 
assign P1_R2144_U134 = ~(P1_R2144_U91 & P1_R2144_U109); 
assign P1_R2144_U158 = ~(P1_R2144_U117 & P1_R2144_U110 & P1_R2144_U55); 
assign P1_R2144_U238 = ~(P1_R2144_U163 & P1_R2144_U91); 
assign P1_R2278_U29 = ~P1_U2800; 
assign P1_R2278_U32 = ~(P1_U2800 & P1_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P1_R2278_U610 = ~(P1_U2800 & P1_R2278_U30); 
assign P1_R2358_U457 = ~(P1_U2352 & P1_R2358_U157); 
assign P1_R2358_U472 = ~(P1_U2352 & P1_R2358_U157); 
assign P1_R2099_U81 = ~(P1_R2099_U336 & P1_R2099_U335); 
assign P1_R2099_U82 = ~(P1_R2099_U338 & P1_R2099_U337); 
assign P1_R2099_U166 = ~P1_R2099_U142; 
assign P1_R2099_U167 = ~P1_R2099_U13; 
assign P1_R2099_U332 = ~(P1_R2099_U56 & P1_R2099_U13); 
assign P1_R2099_U334 = ~(P1_R2099_U59 & P1_R2099_U142); 
assign P1_R2337_U84 = ~(P1_R2337_U168 & P1_R2337_U167); 
assign P1_R2337_U109 = ~P1_R2337_U36; 
assign P1_R2337_U165 = ~(P1_R2337_U36 & P1_PHYADDRPOINTER_REG_18__SCAN_IN); 
assign P1_R2096_U84 = ~(P1_R2096_U168 & P1_R2096_U167); 
assign P1_R2096_U109 = ~P1_R2096_U36; 
assign P1_R2096_U165 = ~(P1_R2096_U36 & P1_REIP_REG_18__SCAN_IN); 
assign P1_LT_563_U8 = ~P1_U3491; 
assign P1_LT_563_U9 = ~P1_U3490; 
assign P1_LT_563_U12 = ~P1_U3489; 
assign P1_LT_563_U15 = ~P1_U3492; 
assign P1_LT_563_U16 = ~P1_U3493; 
assign P1_LT_563_U21 = ~(P1_U3491 & P1_LT_563_U7); 
assign P1_LT_563_U22 = ~(P1_U3490 & P1_LT_563_U10); 
assign P1_LT_563_U27 = ~(P1_U3489 & P1_LT_563_U11); 
assign P1_ADD_405_U67 = ~(P1_ADD_405_U136 & P1_ADD_405_U135); 
assign P1_ADD_405_U112 = ~P1_ADD_405_U36; 
assign P1_ADD_405_U145 = ~(P1_ADD_405_U36 & P1_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P1_ADD_515_U66 = ~(P1_ADD_515_U132 & P1_ADD_515_U131); 
assign P1_ADD_515_U109 = ~P1_ADD_515_U36; 
assign P1_ADD_515_U143 = ~(P1_ADD_515_U36 & P1_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_U3760 = P3_U3759 & P3_U3758 & P3_U5843; 
assign P3_U3962 = P3_U6474 & P3_U6473 & P3_U6476 & P3_U6475; 
assign P3_U5822 = ~(P3_U4318 & P3_U5820); 
assign P3_U5848 = ~(P3_ADD_360_1242_U106 & P3_U2395); 
assign P3_U5872 = ~(P3_ADD_360_1242_U4 & P3_U2395); 
assign P3_U6018 = ~(P3_ADD_558_U89 & P3_U3220); 
assign P3_U6019 = ~(P3_ADD_553_U89 & P3_U4298); 
assign P3_U6020 = ~(P3_ADD_547_U89 & P3_U4299); 
assign P3_U6023 = ~(P3_ADD_531_U89 & P3_U2354); 
assign P3_U6031 = ~(P3_ADD_385_U89 & P3_U2358); 
assign P3_U6032 = ~(P3_ADD_380_U89 & P3_U2359); 
assign P3_U6033 = ~(P3_ADD_349_U89 & P3_U4306); 
assign P3_U6034 = ~(P3_ADD_344_U89 & P3_U2362); 
assign P3_U6045 = ~(P3_ADD_541_U84 & P3_U4300); 
assign P3_U6046 = ~(P3_ADD_536_U84 & P3_U4301); 
assign P3_U6049 = ~(P3_ADD_515_U84 & P3_U4302); 
assign P3_U6050 = ~(P3_ADD_494_U84 & P3_U2356); 
assign P3_U6051 = ~(P3_ADD_476_U84 & P3_U4303); 
assign P3_U6052 = ~(P3_ADD_441_U84 & P3_U4304); 
assign P3_U6053 = ~(P3_ADD_405_U84 & P3_U4305); 
assign P3_U6054 = ~(P3_ADD_394_U84 & P3_U2357); 
assign P3_U6360 = ~(P3_ADD_526_U59 & P3_U2355); 
assign P3_U6479 = ~(P3_U2396 & P3_ADD_360_1242_U106); 
assign P3_U6487 = ~(P3_U2396 & P3_ADD_360_1242_U4); 
assign P3_U6541 = ~(P3_ADD_318_U84 & P3_U2398); 
assign P3_U6546 = ~(P3_ADD_339_U84 & P3_U2388); 
assign P3_U6550 = ~(P3_ADD_315_U80 & P3_U2397); 
assign P3_U6991 = ~(P3_ADD_546_U59 & P3_U2400); 
assign P3_U7089 = ~(P3_ADD_552_U59 & P3_U2399); 
assign P3_U7246 = ~(P3_ADD_467_U84 & P3_U2601); 
assign P3_U7248 = ~(P3_ADD_430_U84 & P3_U2405); 
assign P3_U7349 = ~(P3_SUB_414_U62 & P3_U2602); 
assign P2_U3297 = ~P2_R2167_U6; 
assign P2_U3305 = ~(P2_R2167_U6 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U3319 = ~(P2_U3352 & P2_U3314); 
assign P2_U3338 = ~(P2_R2182_U69 & P2_U3352); 
assign P2_U3892 = P2_U5653 & P2_U5654; 
assign P2_U4635 = ~P2_U3352; 
assign P2_U5580 = ~(P2_U4436 & P2_R2167_U6); 
assign P2_U6227 = ~(P2_U4057 & P2_U4421 & P2_R2167_U6); 
assign P2_U6567 = ~(P2_U4433 & P2_R2167_U6); 
assign P2_U7183 = ~(P2_U4280 & P2_U4279 & P2_U4278 & P2_U4277); 
assign P2_U7200 = ~(P2_U4284 & P2_U4283 & P2_U4282 & P2_U4281); 
assign P2_U7234 = ~(P2_U4292 & P2_U4291 & P2_U4290 & P2_U4289); 
assign P2_U7268 = ~(P2_U4300 & P2_U4299 & P2_U4298 & P2_U4297); 
assign P2_U7302 = ~(P2_U4308 & P2_U4307 & P2_U4306 & P2_U4305); 
assign P2_U7336 = ~(P2_U4316 & P2_U4315 & P2_U4314 & P2_U4313); 
assign P2_U7370 = ~(P2_U4324 & P2_U4323 & P2_U4322 & P2_U4321); 
assign P2_U7404 = ~(P2_U4332 & P2_U4331 & P2_U4330 & P2_U4329); 
assign P2_U8050 = ~(P2_R2167_U6 & P2_U4435); 
assign P2_U8063 = ~(P2_U4637 & P2_U3316); 
assign P2_U8071 = ~(P2_U4433 & P2_U2359 & P2_R2167_U6); 
assign P2_U8120 = ~(P2_U8118 & P2_R2167_U6); 
assign P2_U8316 = ~(P2_U3242 & P2_R2267_U19); 
assign P2_U8401 = ~(P2_R2337_U82 & P2_U3284); 
assign P1_U2360 = P1_U3414 & P1_STATE2_REG_2__SCAN_IN; 
assign P1_U2362 = P1_U2359 & P1_U4208; 
assign P1_U2363 = P1_U2359 & P1_U4210; 
assign P1_U2370 = P1_U3414 & P1_U3263; 
assign P1_U2377 = P1_U3762 & P1_U3414; 
assign P1_U2486 = ~(P1_R2144_U43 | P1_R2144_U50); 
assign P1_U2649 = P1_R2144_U50 & P1_U6746; 
assign P1_U2666 = ~(P1_U6837 & P1_U4025); 
assign P1_U2673 = ~(P1_U7458 & P1_U7457); 
assign P1_U2674 = ~(P1_U7460 & P1_U7459); 
assign P1_U2675 = ~(P1_U4168 & P1_U7463); 
assign P1_U2676 = ~(P1_U4169 & P1_U7466); 
assign P1_U2677 = ~(P1_U7794 & P1_U7793 & P1_U7467); 
assign P1_U2906 = ~(P1_U3882 & P1_U6146); 
assign P1_U2907 = ~(P1_U3881 & P1_U6143); 
assign P1_U2908 = ~(P1_U3880 & P1_U6140); 
assign P1_U2909 = ~(P1_U3879 & P1_U6137); 
assign P1_U2910 = ~(P1_U3878 & P1_U6134); 
assign P1_U2911 = ~(P1_U3877 & P1_U6131); 
assign P1_U2912 = ~(P1_U3876 & P1_U6128); 
assign P1_U2913 = ~(P1_U3875 & P1_U6125); 
assign P1_U2914 = ~(P1_U3874 & P1_U6122); 
assign P1_U2915 = ~(P1_U3873 & P1_U6119); 
assign P1_U2916 = ~(P1_U3872 & P1_U6116); 
assign P1_U2917 = ~(P1_U3871 & P1_U6113); 
assign P1_U2918 = ~(P1_U3870 & P1_U6110); 
assign P1_U2919 = ~(P1_U3869 & P1_U6107); 
assign P1_U2920 = ~(P1_U3868 & P1_U6104); 
assign P1_U3310 = ~P1_R2144_U50; 
assign P1_U3313 = ~(P1_R2144_U50 & P1_R2144_U43); 
assign P1_U3325 = ~(P1_R2144_U50 & P1_U3309); 
assign P1_U3468 = ~(P1_U7702 & P1_U7701); 
assign P1_U3469 = ~(P1_U7709 & P1_U7708); 
assign P1_U3472 = ~(P1_U7722 & P1_U7721); 
assign P1_U3473 = ~(P1_U7724 & P1_U7723); 
assign P1_U3474 = ~(P1_U7728 & P1_U7727); 
assign P1_U3484 = ~(P1_U7763 & P1_U7762); 
assign P1_U5553 = ~(P1_U4226 & P1_R2144_U50); 
assign P1_U5564 = ~P1_U3414; 
assign P1_U5884 = ~(P1_R2337_U84 & P1_U2376); 
assign P1_U6154 = ~(P1_U2422 & U346); 
assign P1_U6157 = ~(P1_U2422 & U335); 
assign P1_U6160 = ~(P1_U2422 & U324); 
assign P1_U6163 = ~(P1_U2422 & U321); 
assign P1_U6166 = ~(P1_U2422 & U320); 
assign P1_U6169 = ~(P1_U2422 & U319); 
assign P1_U6172 = ~(P1_U2422 & U318); 
assign P1_U6175 = ~(P1_U2422 & U317); 
assign P1_U6178 = ~(P1_U2422 & U316); 
assign P1_U6181 = ~(P1_U2422 & U315); 
assign P1_U6184 = ~(P1_U2422 & U345); 
assign P1_U6187 = ~(P1_U2422 & U344); 
assign P1_U6190 = ~(P1_U2422 & U343); 
assign P1_U6193 = ~(P1_U2422 & U342); 
assign P1_U6196 = ~(P1_U2422 & U341); 
assign P1_U6199 = ~(P1_U2422 & U340); 
assign P1_U6202 = ~(P1_U2423 & U339); 
assign P1_U6203 = ~(P1_U2387 & U346); 
assign P1_U6206 = ~(P1_U2423 & U338); 
assign P1_U6207 = ~(P1_U2387 & U335); 
assign P1_U6210 = ~(P1_U2423 & U337); 
assign P1_U6211 = ~(P1_U2387 & U324); 
assign P1_U6214 = ~(P1_U2423 & U336); 
assign P1_U6215 = ~(P1_U2387 & U321); 
assign P1_U6218 = ~(P1_U2423 & U334); 
assign P1_U6219 = ~(P1_U2387 & U320); 
assign P1_U6222 = ~(P1_U2423 & U333); 
assign P1_U6223 = ~(P1_U2387 & U319); 
assign P1_U6226 = ~(P1_U2423 & U332); 
assign P1_U6227 = ~(P1_U2387 & U318); 
assign P1_U6230 = ~(P1_U2423 & U331); 
assign P1_U6231 = ~(P1_U2387 & U317); 
assign P1_U6234 = ~(P1_U2423 & U330); 
assign P1_U6235 = ~(P1_U2387 & U316); 
assign P1_U6238 = ~(P1_U2423 & U329); 
assign P1_U6239 = ~(P1_U2387 & U315); 
assign P1_U6242 = ~(P1_U2423 & U328); 
assign P1_U6243 = ~(P1_U2387 & U345); 
assign P1_U6246 = ~(P1_U2423 & U327); 
assign P1_U6247 = ~(P1_U2387 & U344); 
assign P1_U6250 = ~(P1_U2423 & U326); 
assign P1_U6251 = ~(P1_U2387 & U343); 
assign P1_U6254 = ~(P1_U2423 & U325); 
assign P1_U6255 = ~(P1_U2387 & U342); 
assign P1_U6258 = ~(P1_U2423 & U323); 
assign P1_U6259 = ~(P1_U2387 & U341); 
assign P1_U6262 = ~(P1_U2423 & U322); 
assign P1_U6305 = ~(P1_U2371 & P1_R2099_U82); 
assign P1_U6308 = ~(P1_U2371 & P1_R2099_U81); 
assign P1_U6372 = ~(P1_U2426 & P1_R2182_U34); 
assign P1_U6373 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_0__SCAN_IN); 
assign P1_U6375 = ~(P1_U6363 & P1_REIP_REG_0__SCAN_IN); 
assign P1_U6380 = ~(P1_U2426 & P1_R2182_U33); 
assign P1_U6381 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_1__SCAN_IN); 
assign P1_U6383 = ~(P1_U6363 & P1_REIP_REG_1__SCAN_IN); 
assign P1_U6388 = ~(P1_U2426 & P1_R2182_U42); 
assign P1_U6389 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_2__SCAN_IN); 
assign P1_U6391 = ~(P1_U6363 & P1_REIP_REG_2__SCAN_IN); 
assign P1_U6396 = ~(P1_U2426 & P1_R2182_U25); 
assign P1_U6397 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_3__SCAN_IN); 
assign P1_U6399 = ~(P1_U6363 & P1_REIP_REG_3__SCAN_IN); 
assign P1_U6404 = ~(P1_U2426 & P1_R2182_U24); 
assign P1_U6405 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_4__SCAN_IN); 
assign P1_U6407 = ~(P1_U6363 & P1_REIP_REG_4__SCAN_IN); 
assign P1_U6412 = ~(P1_R2182_U5 & P1_U2426); 
assign P1_U6413 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_5__SCAN_IN); 
assign P1_U6415 = ~(P1_U6363 & P1_REIP_REG_5__SCAN_IN); 
assign P1_U6419 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_6__SCAN_IN); 
assign P1_U6422 = ~(P1_U6363 & P1_REIP_REG_6__SCAN_IN); 
assign P1_U6426 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_7__SCAN_IN); 
assign P1_U6429 = ~(P1_U6363 & P1_REIP_REG_7__SCAN_IN); 
assign P1_U6433 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_8__SCAN_IN); 
assign P1_U6436 = ~(P1_U6363 & P1_REIP_REG_8__SCAN_IN); 
assign P1_U6440 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_9__SCAN_IN); 
assign P1_U6443 = ~(P1_U6363 & P1_REIP_REG_9__SCAN_IN); 
assign P1_U6447 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_10__SCAN_IN); 
assign P1_U6450 = ~(P1_U6363 & P1_REIP_REG_10__SCAN_IN); 
assign P1_U6454 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_11__SCAN_IN); 
assign P1_U6457 = ~(P1_U6363 & P1_REIP_REG_11__SCAN_IN); 
assign P1_U6461 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_12__SCAN_IN); 
assign P1_U6464 = ~(P1_U6363 & P1_REIP_REG_12__SCAN_IN); 
assign P1_U6468 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_13__SCAN_IN); 
assign P1_U6471 = ~(P1_U6363 & P1_REIP_REG_13__SCAN_IN); 
assign P1_U6475 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_14__SCAN_IN); 
assign P1_U6478 = ~(P1_U6363 & P1_REIP_REG_14__SCAN_IN); 
assign P1_U6482 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_15__SCAN_IN); 
assign P1_U6485 = ~(P1_U6363 & P1_REIP_REG_15__SCAN_IN); 
assign P1_U6489 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_16__SCAN_IN); 
assign P1_U6492 = ~(P1_U6363 & P1_REIP_REG_16__SCAN_IN); 
assign P1_U6496 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_17__SCAN_IN); 
assign P1_U6499 = ~(P1_U6363 & P1_REIP_REG_17__SCAN_IN); 
assign P1_U6503 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_18__SCAN_IN); 
assign P1_U6506 = ~(P1_U6363 & P1_REIP_REG_18__SCAN_IN); 
assign P1_U6510 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_19__SCAN_IN); 
assign P1_U6513 = ~(P1_U6363 & P1_REIP_REG_19__SCAN_IN); 
assign P1_U6517 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_20__SCAN_IN); 
assign P1_U6520 = ~(P1_U6363 & P1_REIP_REG_20__SCAN_IN); 
assign P1_U6524 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_21__SCAN_IN); 
assign P1_U6527 = ~(P1_U6363 & P1_REIP_REG_21__SCAN_IN); 
assign P1_U6531 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_22__SCAN_IN); 
assign P1_U6534 = ~(P1_U6363 & P1_REIP_REG_22__SCAN_IN); 
assign P1_U6538 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_23__SCAN_IN); 
assign P1_U6541 = ~(P1_U6363 & P1_REIP_REG_23__SCAN_IN); 
assign P1_U6545 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_24__SCAN_IN); 
assign P1_U6548 = ~(P1_U6363 & P1_REIP_REG_24__SCAN_IN); 
assign P1_U6552 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_25__SCAN_IN); 
assign P1_U6555 = ~(P1_U6363 & P1_REIP_REG_25__SCAN_IN); 
assign P1_U6559 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_26__SCAN_IN); 
assign P1_U6562 = ~(P1_U6363 & P1_REIP_REG_26__SCAN_IN); 
assign P1_U6566 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_27__SCAN_IN); 
assign P1_U6569 = ~(P1_U6363 & P1_REIP_REG_27__SCAN_IN); 
assign P1_U6573 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_28__SCAN_IN); 
assign P1_U6576 = ~(P1_U6363 & P1_REIP_REG_28__SCAN_IN); 
assign P1_U6580 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_29__SCAN_IN); 
assign P1_U6583 = ~(P1_U6363 & P1_REIP_REG_29__SCAN_IN); 
assign P1_U6587 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_30__SCAN_IN); 
assign P1_U6590 = ~(P1_U6363 & P1_REIP_REG_30__SCAN_IN); 
assign P1_U6594 = ~(P1_U2373 & P1_PHYADDRPOINTER_REG_31__SCAN_IN); 
assign P1_U6597 = ~(P1_U6363 & P1_REIP_REG_31__SCAN_IN); 
assign P1_U6836 = ~(P1_R2337_U84 & P1_U2352); 
assign P1_U6886 = ~(P1_U4159 & P1_R2144_U50); 
assign P1_U7766 = ~(P1_U6603 & P1_REQUESTPENDING_REG_SCAN_IN); 
assign P1_U7772 = ~(P1_U6614 & P1_READREQUEST_REG_SCAN_IN); 
assign P3_ADD_526_U156 = ~(P3_ADD_526_U129 & P3_ADD_526_U98); 
assign P3_ADD_552_U156 = ~(P3_ADD_552_U129 & P3_ADD_552_U98); 
assign P3_ADD_546_U156 = ~(P3_ADD_546_U129 & P3_ADD_546_U98); 
assign P3_ADD_476_U38 = ~(P3_ADD_476_U109 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_476_U166 = ~(P3_ADD_476_U109 & P3_ADD_476_U37); 
assign P3_ADD_531_U39 = ~(P3_ADD_531_U113 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_531_U175 = ~(P3_ADD_531_U113 & P3_ADD_531_U38); 
assign P3_SUB_320_U9 = P3_SUB_320_U120 & P3_SUB_320_U31; 
assign P3_SUB_320_U75 = ~P3_ADD_318_U84; 
assign P3_SUB_320_U96 = ~P3_SUB_320_U31; 
assign P3_SUB_320_U152 = ~(P3_ADD_318_U84 & P3_SUB_320_U31); 
assign P3_ADD_318_U38 = ~(P3_ADD_318_U109 & P3_PHYADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_318_U166 = ~(P3_ADD_318_U109 & P3_ADD_318_U37); 
assign P3_ADD_315_U38 = ~(P3_ADD_315_U106 & P3_PHYADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_315_U158 = ~(P3_ADD_315_U106 & P3_ADD_315_U37); 
assign P3_ADD_360_1242_U84 = ~(P3_ADD_360_1242_U256 & P3_ADD_360_1242_U255); 
assign P3_ADD_360_1242_U154 = ~P3_ADD_360_1242_U46; 
assign P3_ADD_360_1242_U182 = ~(P3_ADD_360_1242_U47 & P3_ADD_360_1242_U46); 
assign P3_ADD_360_1242_U184 = ~(P3_ADD_360_1242_U44 & P3_ADD_360_1242_U183); 
assign P3_ADD_467_U38 = ~(P3_ADD_467_U109 & P3_REIP_REG_18__SCAN_IN); 
assign P3_ADD_467_U166 = ~(P3_ADD_467_U109 & P3_ADD_467_U37); 
assign P3_ADD_430_U38 = ~(P3_ADD_430_U109 & P3_REIP_REG_18__SCAN_IN); 
assign P3_ADD_430_U166 = ~(P3_ADD_430_U109 & P3_ADD_430_U37); 
assign P3_ADD_380_U39 = ~(P3_ADD_380_U113 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_380_U175 = ~(P3_ADD_380_U113 & P3_ADD_380_U38); 
assign P3_ADD_344_U39 = ~(P3_ADD_344_U113 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_344_U175 = ~(P3_ADD_344_U113 & P3_ADD_344_U38); 
assign P3_LT_563_U21 = ~(P3_LT_563_U19 & P3_LT_563_U20 & P3_LT_563_U18); 
assign P3_ADD_339_U38 = ~(P3_ADD_339_U109 & P3_PHYADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_339_U166 = ~(P3_ADD_339_U109 & P3_ADD_339_U37); 
assign P3_ADD_541_U38 = ~(P3_ADD_541_U109 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_541_U166 = ~(P3_ADD_541_U109 & P3_ADD_541_U37); 
assign P3_SUB_357_1258_U90 = ~(P3_SUB_357_1258_U463 & P3_SUB_357_1258_U462); 
assign P3_SUB_357_1258_U91 = ~(P3_SUB_357_1258_U470 & P3_SUB_357_1258_U469); 
assign P3_SUB_357_1258_U92 = ~(P3_SUB_357_1258_U477 & P3_SUB_357_1258_U476); 
assign P3_SUB_357_1258_U93 = ~(P3_SUB_357_1258_U482 & P3_SUB_357_1258_U481); 
assign P3_SUB_357_1258_U196 = ~P3_SUB_357_1258_U145; 
assign P3_SUB_357_1258_U198 = ~(P3_SUB_357_1258_U197 & P3_SUB_357_1258_U145); 
assign P3_SUB_357_1258_U255 = ~(P3_SUB_357_1258_U114 & P3_SUB_357_1258_U253); 
assign P3_SUB_357_1258_U455 = ~(P3_SUB_357_1258_U144 & P3_SUB_357_1258_U145); 
assign P3_ADD_515_U38 = ~(P3_ADD_515_U109 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_515_U166 = ~(P3_ADD_515_U109 & P3_ADD_515_U37); 
assign P3_ADD_394_U38 = ~(P3_ADD_394_U112 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_394_U170 = ~(P3_ADD_394_U112 & P3_ADD_394_U37); 
assign P3_SUB_414_U51 = ~(P3_SUB_414_U137 & P3_SUB_414_U136); 
assign P3_ADD_441_U38 = ~(P3_ADD_441_U109 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_441_U166 = ~(P3_ADD_441_U109 & P3_ADD_441_U37); 
assign P3_ADD_349_U39 = ~(P3_ADD_349_U113 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_349_U175 = ~(P3_ADD_349_U113 & P3_ADD_349_U38); 
assign P3_ADD_405_U38 = ~(P3_ADD_405_U112 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_405_U170 = ~(P3_ADD_405_U112 & P3_ADD_405_U37); 
assign P3_ADD_553_U39 = ~(P3_ADD_553_U113 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_553_U175 = ~(P3_ADD_553_U113 & P3_ADD_553_U38); 
assign P3_ADD_558_U39 = ~(P3_ADD_558_U113 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_558_U175 = ~(P3_ADD_558_U113 & P3_ADD_558_U38); 
assign P3_ADD_385_U39 = ~(P3_ADD_385_U113 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_385_U175 = ~(P3_ADD_385_U113 & P3_ADD_385_U38); 
assign P3_ADD_547_U39 = ~(P3_ADD_547_U113 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_ADD_547_U175 = ~(P3_ADD_547_U113 & P3_ADD_547_U38); 
assign P3_ADD_371_1212_U5 = P3_ADD_371_1212_U196 & P3_ADD_371_1212_U48; 
assign P3_ADD_371_1212_U49 = ~(P3_ADD_371_1212_U100 & P3_ADD_371_1212_U117); 
assign P3_ADD_371_1212_U109 = P3_ADD_371_1212_U205 & P3_ADD_371_1212_U204; 
assign P3_ADD_371_1212_U193 = ~(P3_ADD_371_1212_U117 & P3_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P3_ADD_371_1212_U262 = ~(P3_ADD_371_1212_U117 & P3_ADD_371_1212_U46); 
assign P3_ADD_494_U38 = ~(P3_ADD_494_U109 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_494_U166 = ~(P3_ADD_494_U109 & P3_ADD_494_U37); 
assign P3_ADD_536_U38 = ~(P3_ADD_536_U109 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_536_U166 = ~(P3_ADD_536_U109 & P3_ADD_536_U37); 
assign P2_R2099_U69 = ~(P2_R2099_U154 & P2_R2099_U153); 
assign P2_R2099_U123 = ~P2_R2099_U21; 
assign P2_R2099_U151 = ~(P2_U2739 & P2_R2099_U21); 
assign P2_ADD_391_1196_U32 = ~P2_R2096_U70; 
assign P2_ADD_391_1196_U167 = ~(P2_ADD_391_1196_U166 & P2_ADD_391_1196_U123); 
assign P2_ADD_391_1196_U306 = ~(P2_ADD_391_1196_U423 & P2_ADD_391_1196_U23); 
assign P2_ADD_391_1196_U344 = ~(P2_R2096_U77 & P2_ADD_391_1196_U24); 
assign P2_ADD_391_1196_U346 = ~(P2_R2096_U77 & P2_ADD_391_1196_U24); 
assign P2_R2182_U76 = ~(P2_R2182_U216 & P2_R2182_U215); 
assign P2_R2182_U102 = ~(P2_R2182_U135 & P2_R2182_U134); 
assign P2_R2182_U209 = ~(P2_R2182_U132 & P2_R2182_U207); 
assign P2_R2027_U39 = ~(P2_R2027_U113 & P2_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P2_R2027_U175 = ~(P2_R2027_U113 & P2_R2027_U38); 
assign P2_R2337_U39 = ~(P2_R2337_U110 & P2_PHYADDRPOINTER_REG_19__SCAN_IN); 
assign P2_R2337_U164 = ~(P2_R2337_U110 & P2_R2337_U38); 
assign P2_R2096_U19 = P2_U2638 & P2_R2096_U24; 
assign P2_R2096_U69 = ~(P2_R2096_U172 & P2_R2096_U171); 
assign P2_R2096_U146 = ~P2_R2096_U24; 
assign P2_R2096_U260 = ~(P2_R2096_U27 & P2_R2096_U24); 
assign P2_R2096_U263 = ~(P2_R2096_U145 & P2_U2639); 
assign P2_R1957_U9 = P2_R1957_U120 & P2_R1957_U30; 
assign P2_R1957_U75 = ~P2_U3674; 
assign P2_R1957_U96 = ~P2_R1957_U30; 
assign P2_R1957_U152 = ~(P2_U3674 & P2_R1957_U30); 
assign P2_ADD_394_U38 = ~(P2_ADD_394_U112 & P2_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P2_ADD_394_U146 = ~(P2_ADD_394_U112 & P2_ADD_394_U37); 
assign P2_R2267_U30 = ~(P2_R2267_U44 & P2_R2267_U92); 
assign P2_R2267_U94 = ~(P2_R2267_U92 & P2_R2267_U55); 
assign P2_R2267_U136 = ~(P2_R2267_U92 & P2_R2267_U55); 
assign P1_R2027_U156 = ~(P1_R2027_U129 & P1_R2027_U98); 
assign P1_R2144_U83 = ~(P1_R2144_U56 & P1_R2144_U158); 
assign P1_R2144_U84 = ~(P1_R2144_U111 & P1_R2144_U118); 
assign P1_R2144_U135 = ~(P1_R2144_U134 & P1_R2144_U116); 
assign P1_R2144_U138 = ~(P1_R2144_U134 & P1_R2144_U116 & P1_R2144_U137); 
assign P1_R2144_U160 = ~(P1_R2144_U58 & P1_R2144_U158); 
assign P1_R2144_U239 = ~(P1_R2144_U48 & P1_R2144_U133); 
assign P1_R2278_U232 = ~P1_R2278_U32; 
assign P1_R2278_U555 = ~(P1_R2278_U32 & P1_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P1_R2278_U609 = ~(P1_R2278_U29 & P1_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P1_R2358_U11 = P1_R2358_U458 & P1_R2358_U457; 
assign P1_R2358_U31 = ~P1_U2650; 
assign P1_R2358_U209 = ~(P1_U2650 & P1_R2358_U430); 
assign P1_R2358_U474 = ~(P1_R2358_U473 & P1_R2358_U472); 
assign P1_R2099_U14 = ~(P1_R2099_U95 & P1_R2099_U167); 
assign P1_R2099_U141 = ~(P1_R2099_U167 & P1_R2099_U56); 
assign P1_R2099_U331 = ~(P1_R2099_U279 & P1_R2099_U167); 
assign P1_R2099_U333 = ~(P1_R2099_U166 & P1_R2099_U276); 
assign P1_R2337_U38 = ~(P1_R2337_U109 & P1_PHYADDRPOINTER_REG_18__SCAN_IN); 
assign P1_R2337_U166 = ~(P1_R2337_U109 & P1_R2337_U37); 
assign P1_R2096_U38 = ~(P1_R2096_U109 & P1_REIP_REG_18__SCAN_IN); 
assign P1_R2096_U166 = ~(P1_R2096_U109 & P1_R2096_U37); 
assign P1_LT_563_U13 = P1_LT_563_U21 & P1_LT_563_U22; 
assign P1_LT_563_U17 = ~(P1_LT_563_U16 & P1_LT_563_U15 & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P1_LT_563_U18 = ~(P1_LT_563_U15 & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P1_LT_563_U19 = ~(P1_LT_563_U8 & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P1_LT_563_U24 = ~(P1_LT_563_U9 & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P1_LT_563_U25 = ~(P1_LT_563_U12 & P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P1_LT_563_U28 = ~(P1_LT_563_U16 & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P1_ADD_405_U38 = ~(P1_ADD_405_U112 & P1_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P1_ADD_405_U146 = ~(P1_ADD_405_U112 & P1_ADD_405_U37); 
assign P1_ADD_515_U38 = ~(P1_ADD_515_U109 & P1_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P1_ADD_515_U144 = ~(P1_ADD_515_U109 & P1_ADD_515_U37); 
assign P3_U2673 = ~(P3_U7090 & P3_U7088 & P3_U7089); 
assign P3_U2705 = ~(P3_U6989 & P3_U6988 & P3_U6992 & P3_U6990 & P3_U6991); 
assign P3_U2822 = ~(P3_U6470 & P3_U6469 & P3_U6472 & P3_U6471 & P3_U3962); 
assign P3_U2855 = ~(P3_U5823 & P3_U5821 & P3_U5822); 
assign P3_U3761 = P3_U3762 & P3_U5848; 
assign P3_U3813 = P3_U6020 & P3_U6019; 
assign P3_U3815 = P3_U6022 & P3_U6021 & P3_U6023 & P3_U3814; 
assign P3_U3817 = P3_U6034 & P3_U6033 & P3_U6032 & P3_U6031; 
assign P3_U3821 = P3_U6049 & P3_U6048; 
assign P3_U3822 = P3_U6051 & P3_U6050 & P3_U6052 & P3_U6054 & P3_U6053; 
assign P3_U4090 = P3_U7245 & P3_U4316 & P3_U7246; 
assign P3_U5844 = ~(P3_U3757 & P3_U5826 & P3_U5825 & P3_U3754 & P3_U3760); 
assign P3_U5867 = ~(P3_ADD_371_1212_U109 & P3_U2360); 
assign P3_U5873 = ~(P3_SUB_357_1258_U93 & P3_U2393); 
assign P3_U5891 = ~(P3_ADD_371_1212_U5 & P3_U2360); 
assign P3_U5896 = ~(P3_ADD_360_1242_U84 & P3_U2395); 
assign P3_U5897 = ~(P3_SUB_357_1258_U92 & P3_U2393); 
assign P3_U5921 = ~(P3_SUB_357_1258_U91 & P3_U2393); 
assign P3_U5969 = ~(P3_SUB_357_1258_U90 & P3_U2393); 
assign P3_U6483 = ~(P3_U2387 & P3_ADD_371_1212_U109); 
assign P3_U6488 = ~(P3_U2394 & P3_SUB_357_1258_U93); 
assign P3_U6491 = ~(P3_U2387 & P3_ADD_371_1212_U5); 
assign P3_U6495 = ~(P3_U2396 & P3_ADD_360_1242_U84); 
assign P3_U6496 = ~(P3_U2394 & P3_SUB_357_1258_U92); 
assign P3_U6504 = ~(P3_U2394 & P3_SUB_357_1258_U91); 
assign P3_U6520 = ~(P3_U2394 & P3_SUB_357_1258_U90); 
assign P3_U7358 = ~(P3_SUB_414_U51 & P3_U2602); 
assign P2_U2462 = P2_R2182_U76 & P2_R2182_U40; 
assign P2_U2475 = P2_U4635 & P2_R2182_U69; 
assign P2_U2501 = ~(P2_R2182_U40 | P2_R2182_U76); 
assign P2_U2513 = P2_U5580 & P2_U5579; 
assign P2_U3317 = ~P2_R2182_U76; 
assign P2_U3353 = ~(P2_U4635 & P2_U3314); 
assign P2_U3378 = ~(P2_R2182_U76 & P2_U3316); 
assign P2_U3579 = ~(P2_U8063 & P2_U8062); 
assign P2_U3673 = ~(P2_U8402 & P2_U8401); 
assign P2_U4469 = ~P2_U3305; 
assign P2_U4636 = ~P2_U3319; 
assign P2_U4639 = ~(P2_R2182_U76 & P2_U3318); 
assign P2_U4656 = ~(P2_U4655 & P2_U3304 & P2_U3305); 
assign P2_U4709 = ~P2_U3338; 
assign P2_U5649 = ~(P2_R2182_U76 & P2_U5644); 
assign P2_U6229 = ~(P2_U6228 & P2_U6227); 
assign P2_U6469 = ~(P2_U4435 & P2_U3297); 
assign P2_U6568 = ~(P2_U6567 & P2_U6566); 
assign P2_U8051 = ~(P2_U4604 & P2_U3297); 
assign P2_U8054 = ~(P2_U4427 & P2_U3297); 
assign P2_U8070 = ~(P2_U4435 & P2_U3297); 
assign P2_U8119 = ~(P2_U3253 & P2_U3278 & P2_U3297); 
assign P2_U8146 = ~(P2_U2616 & P2_U3297); 
assign P2_U8298 = ~(P2_U2616 & P2_U7183); 
assign P2_U8300 = ~(P2_U2616 & P2_U7200); 
assign P2_U8302 = ~(P2_U2616 & P2_U7234); 
assign P2_U8304 = ~(P2_U2616 & P2_U7268); 
assign P2_U8306 = ~(P2_U2616 & P2_U7302); 
assign P2_U8308 = ~(P2_U2616 & P2_U7336); 
assign P2_U8310 = ~(P2_U2616 & P2_U7370); 
assign P2_U8312 = ~(P2_U2616 & P2_U7404); 
assign P1_U2369 = P1_U2362 & P1_U4497; 
assign P1_U2374 = P1_U2360 & P1_U4214; 
assign P1_U2375 = P1_U2360 & P1_U4216; 
assign P1_U2378 = P1_U2360 & P1_U5569; 
assign P1_U2379 = P1_U2363 & P1_U3280; 
assign P1_U2380 = P1_U2360 & P1_U7608; 
assign P1_U2799 = ~(P1_U4028 & P1_U6887 & P1_U6886); 
assign P1_U3331 = ~(P1_R2144_U43 & P1_U3310); 
assign P1_U3485 = ~(P1_U7767 & P1_U7766); 
assign P1_U3487 = ~(P1_U7773 & P1_U7772); 
assign P1_U3753 = P1_U5552 & P1_U5553; 
assign P1_U4024 = P1_U6834 & P1_U6835 & P1_U6836; 
assign P1_U4229 = ~(P1_U2362 & P1_U3272); 
assign P1_U4230 = ~(P1_U2363 & P1_U4377); 
assign P1_U4524 = ~P1_U3325; 
assign P1_U4528 = ~P1_U3313; 
assign P1_U5575 = ~(P1_U2370 & P1_REIP_REG_0__SCAN_IN); 
assign P1_U5576 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P1_U5582 = ~(P1_U2370 & P1_REIP_REG_1__SCAN_IN); 
assign P1_U5583 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P1_U5589 = ~(P1_U2370 & P1_REIP_REG_2__SCAN_IN); 
assign P1_U5590 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P1_U5596 = ~(P1_U2370 & P1_REIP_REG_3__SCAN_IN); 
assign P1_U5597 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P1_U5603 = ~(P1_U2370 & P1_REIP_REG_4__SCAN_IN); 
assign P1_U5604 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P1_U5610 = ~(P1_U2370 & P1_REIP_REG_5__SCAN_IN); 
assign P1_U5611 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P1_U5617 = ~(P1_U2370 & P1_REIP_REG_6__SCAN_IN); 
assign P1_U5618 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P1_U5624 = ~(P1_U2370 & P1_REIP_REG_7__SCAN_IN); 
assign P1_U5625 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P1_U5631 = ~(P1_U2370 & P1_REIP_REG_8__SCAN_IN); 
assign P1_U5632 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P1_U5638 = ~(P1_U2370 & P1_REIP_REG_9__SCAN_IN); 
assign P1_U5639 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P1_U5645 = ~(P1_U2370 & P1_REIP_REG_10__SCAN_IN); 
assign P1_U5646 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P1_U5652 = ~(P1_U2370 & P1_REIP_REG_11__SCAN_IN); 
assign P1_U5653 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P1_U5659 = ~(P1_U2370 & P1_REIP_REG_12__SCAN_IN); 
assign P1_U5660 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P1_U5666 = ~(P1_U2370 & P1_REIP_REG_13__SCAN_IN); 
assign P1_U5667 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P1_U5673 = ~(P1_U2370 & P1_REIP_REG_14__SCAN_IN); 
assign P1_U5674 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P1_U5680 = ~(P1_U2370 & P1_REIP_REG_15__SCAN_IN); 
assign P1_U5681 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P1_U5687 = ~(P1_U2370 & P1_REIP_REG_16__SCAN_IN); 
assign P1_U5688 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P1_U5694 = ~(P1_U2370 & P1_REIP_REG_17__SCAN_IN); 
assign P1_U5695 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P1_U5701 = ~(P1_U2370 & P1_REIP_REG_18__SCAN_IN); 
assign P1_U5702 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P1_U5708 = ~(P1_U2370 & P1_REIP_REG_19__SCAN_IN); 
assign P1_U5709 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P1_U5715 = ~(P1_U2370 & P1_REIP_REG_20__SCAN_IN); 
assign P1_U5716 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P1_U5722 = ~(P1_U2370 & P1_REIP_REG_21__SCAN_IN); 
assign P1_U5723 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P1_U5729 = ~(P1_U2370 & P1_REIP_REG_22__SCAN_IN); 
assign P1_U5730 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P1_U5736 = ~(P1_U2370 & P1_REIP_REG_23__SCAN_IN); 
assign P1_U5737 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P1_U5743 = ~(P1_U2370 & P1_REIP_REG_24__SCAN_IN); 
assign P1_U5744 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P1_U5750 = ~(P1_U2370 & P1_REIP_REG_25__SCAN_IN); 
assign P1_U5751 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P1_U5757 = ~(P1_U2370 & P1_REIP_REG_26__SCAN_IN); 
assign P1_U5758 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P1_U5764 = ~(P1_U2370 & P1_REIP_REG_27__SCAN_IN); 
assign P1_U5765 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P1_U5771 = ~(P1_U2370 & P1_REIP_REG_28__SCAN_IN); 
assign P1_U5772 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P1_U5778 = ~(P1_U2370 & P1_REIP_REG_29__SCAN_IN); 
assign P1_U5779 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P1_U5785 = ~(P1_U2370 & P1_REIP_REG_30__SCAN_IN); 
assign P1_U5786 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P1_U5792 = ~(P1_U2370 & P1_REIP_REG_31__SCAN_IN); 
assign P1_U5793 = ~(P1_U5564 & P1_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_526_U58 = ~(P3_ADD_526_U156 & P3_ADD_526_U155); 
assign P3_ADD_552_U58 = ~(P3_ADD_552_U156 & P3_ADD_552_U155); 
assign P3_ADD_546_U58 = ~(P3_ADD_546_U156 & P3_ADD_546_U155); 
assign P3_ADD_476_U83 = ~(P3_ADD_476_U166 & P3_ADD_476_U165); 
assign P3_ADD_476_U110 = ~P3_ADD_476_U38; 
assign P3_ADD_476_U163 = ~(P3_ADD_476_U38 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_531_U88 = ~(P3_ADD_531_U175 & P3_ADD_531_U174); 
assign P3_ADD_531_U114 = ~P3_ADD_531_U39; 
assign P3_ADD_531_U172 = ~(P3_ADD_531_U39 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_SUB_320_U117 = ~(P3_SUB_320_U96 & P3_SUB_320_U75); 
assign P3_SUB_320_U153 = ~(P3_SUB_320_U96 & P3_SUB_320_U75); 
assign P3_ADD_318_U83 = ~(P3_ADD_318_U166 & P3_ADD_318_U165); 
assign P3_ADD_318_U110 = ~P3_ADD_318_U38; 
assign P3_ADD_318_U163 = ~(P3_ADD_318_U38 & P3_PHYADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_315_U79 = ~(P3_ADD_315_U158 & P3_ADD_315_U157); 
assign P3_ADD_315_U107 = ~P3_ADD_315_U38; 
assign P3_ADD_315_U155 = ~(P3_ADD_315_U38 & P3_PHYADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_360_1242_U5 = P3_ADD_360_1242_U184 & P3_ADD_360_1242_U46; 
assign P3_ADD_360_1242_U50 = ~(P3_ADD_360_1242_U154 & P3_ADD_360_1242_U99); 
assign P3_ADD_360_1242_U76 = ~(P3_ADD_360_1242_U154 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_467_U83 = ~(P3_ADD_467_U166 & P3_ADD_467_U165); 
assign P3_ADD_467_U110 = ~P3_ADD_467_U38; 
assign P3_ADD_467_U163 = ~(P3_ADD_467_U38 & P3_REIP_REG_19__SCAN_IN); 
assign P3_ADD_430_U83 = ~(P3_ADD_430_U166 & P3_ADD_430_U165); 
assign P3_ADD_430_U110 = ~P3_ADD_430_U38; 
assign P3_ADD_430_U163 = ~(P3_ADD_430_U38 & P3_REIP_REG_19__SCAN_IN); 
assign P3_ADD_380_U88 = ~(P3_ADD_380_U175 & P3_ADD_380_U174); 
assign P3_ADD_380_U114 = ~P3_ADD_380_U39; 
assign P3_ADD_380_U172 = ~(P3_ADD_380_U39 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_344_U88 = ~(P3_ADD_344_U175 & P3_ADD_344_U174); 
assign P3_ADD_344_U114 = ~P3_ADD_344_U39; 
assign P3_ADD_344_U172 = ~(P3_ADD_344_U39 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_LT_563_U24 = ~(P3_LT_563_U22 & P3_LT_563_U23 & P3_LT_563_U21); 
assign P3_ADD_339_U83 = ~(P3_ADD_339_U166 & P3_ADD_339_U165); 
assign P3_ADD_339_U110 = ~P3_ADD_339_U38; 
assign P3_ADD_339_U163 = ~(P3_ADD_339_U38 & P3_PHYADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_541_U83 = ~(P3_ADD_541_U166 & P3_ADD_541_U165); 
assign P3_ADD_541_U110 = ~P3_ADD_541_U38; 
assign P3_ADD_541_U163 = ~(P3_ADD_541_U38 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_SUB_357_1258_U15 = P3_SUB_357_1258_U255 & P3_SUB_357_1258_U252; 
assign P3_SUB_357_1258_U67 = ~(P3_SUB_357_1258_U102 & P3_SUB_357_1258_U198); 
assign P3_SUB_357_1258_U143 = ~(P3_SUB_357_1258_U199 & P3_SUB_357_1258_U198); 
assign P3_SUB_357_1258_U456 = ~(P3_SUB_357_1258_U196 & P3_SUB_357_1258_U454); 
assign P3_ADD_515_U83 = ~(P3_ADD_515_U166 & P3_ADD_515_U165); 
assign P3_ADD_515_U110 = ~P3_ADD_515_U38; 
assign P3_ADD_515_U163 = ~(P3_ADD_515_U38 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_394_U83 = ~(P3_ADD_394_U170 & P3_ADD_394_U169); 
assign P3_ADD_394_U113 = ~P3_ADD_394_U38; 
assign P3_ADD_394_U167 = ~(P3_ADD_394_U38 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_441_U83 = ~(P3_ADD_441_U166 & P3_ADD_441_U165); 
assign P3_ADD_441_U110 = ~P3_ADD_441_U38; 
assign P3_ADD_441_U163 = ~(P3_ADD_441_U38 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_349_U88 = ~(P3_ADD_349_U175 & P3_ADD_349_U174); 
assign P3_ADD_349_U114 = ~P3_ADD_349_U39; 
assign P3_ADD_349_U172 = ~(P3_ADD_349_U39 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_405_U83 = ~(P3_ADD_405_U170 & P3_ADD_405_U169); 
assign P3_ADD_405_U113 = ~P3_ADD_405_U38; 
assign P3_ADD_405_U167 = ~(P3_ADD_405_U38 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_553_U88 = ~(P3_ADD_553_U175 & P3_ADD_553_U174); 
assign P3_ADD_553_U114 = ~P3_ADD_553_U39; 
assign P3_ADD_553_U172 = ~(P3_ADD_553_U39 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_558_U88 = ~(P3_ADD_558_U175 & P3_ADD_558_U174); 
assign P3_ADD_558_U114 = ~P3_ADD_558_U39; 
assign P3_ADD_558_U172 = ~(P3_ADD_558_U39 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_385_U88 = ~(P3_ADD_385_U175 & P3_ADD_385_U174); 
assign P3_ADD_385_U114 = ~P3_ADD_385_U39; 
assign P3_ADD_385_U172 = ~(P3_ADD_385_U39 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_547_U88 = ~(P3_ADD_547_U175 & P3_ADD_547_U174); 
assign P3_ADD_547_U114 = ~P3_ADD_547_U39; 
assign P3_ADD_547_U172 = ~(P3_ADD_547_U39 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_371_1212_U86 = ~(P3_ADD_371_1212_U263 & P3_ADD_371_1212_U262); 
assign P3_ADD_371_1212_U163 = ~P3_ADD_371_1212_U49; 
assign P3_ADD_371_1212_U192 = ~(P3_ADD_371_1212_U50 & P3_ADD_371_1212_U49); 
assign P3_ADD_371_1212_U194 = ~(P3_ADD_371_1212_U47 & P3_ADD_371_1212_U193); 
assign P3_ADD_494_U83 = ~(P3_ADD_494_U166 & P3_ADD_494_U165); 
assign P3_ADD_494_U110 = ~P3_ADD_494_U38; 
assign P3_ADD_494_U163 = ~(P3_ADD_494_U38 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_536_U83 = ~(P3_ADD_536_U166 & P3_ADD_536_U165); 
assign P3_ADD_536_U110 = ~P3_ADD_536_U38; 
assign P3_ADD_536_U163 = ~(P3_ADD_536_U38 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P2_R2099_U24 = ~(P2_U2739 & P2_R2099_U123); 
assign P2_R2099_U152 = ~(P2_R2099_U123 & P2_R2099_U22); 
assign P2_ADD_391_1196_U12 = ~(P2_ADD_391_1196_U144 & P2_ADD_391_1196_U306); 
assign P2_ADD_391_1196_U26 = ~P2_R2182_U76; 
assign P2_ADD_391_1196_U33 = ~P2_R2096_U69; 
assign P2_ADD_391_1196_U118 = ~(P2_ADD_391_1196_U168 & P2_ADD_391_1196_U167); 
assign P2_ADD_391_1196_U122 = P2_ADD_391_1196_U345 & P2_ADD_391_1196_U344; 
assign P2_ADD_391_1196_U170 = P2_R2182_U76 | P2_R2096_U75; 
assign P2_ADD_391_1196_U172 = ~(P2_R2096_U75 & P2_R2182_U76); 
assign P2_ADD_391_1196_U333 = ~(P2_R2182_U76 & P2_ADD_391_1196_U27); 
assign P2_ADD_391_1196_U335 = ~(P2_R2182_U76 & P2_ADD_391_1196_U27); 
assign P2_ADD_391_1196_U348 = ~(P2_ADD_391_1196_U347 & P2_ADD_391_1196_U346); 
assign P2_R2182_U21 = P2_U2676 & P2_R2182_U102; 
assign P2_R2182_U75 = ~(P2_R2182_U209 & P2_R2182_U208); 
assign P2_R2182_U136 = ~P2_R2182_U102; 
assign P2_R2182_U201 = ~(P2_R2182_U24 & P2_R2182_U102); 
assign P2_R2027_U88 = ~(P2_R2027_U175 & P2_R2027_U174); 
assign P2_R2027_U114 = ~P2_R2027_U39; 
assign P2_R2027_U172 = ~(P2_R2027_U39 & P2_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P2_R2337_U81 = ~(P2_R2337_U164 & P2_R2337_U163); 
assign P2_R2337_U111 = ~P2_R2337_U39; 
assign P2_R2337_U161 = ~(P2_R2337_U39 & P2_PHYADDRPOINTER_REG_20__SCAN_IN); 
assign P2_R2096_U20 = P2_U2637 & P2_R2096_U19; 
assign P2_R2096_U97 = ~(P2_R2096_U263 & P2_R2096_U262); 
assign P2_R2096_U147 = ~P2_R2096_U19; 
assign P2_R2096_U258 = ~(P2_R2096_U33 & P2_R2096_U19); 
assign P2_R2096_U261 = ~(P2_R2096_U146 & P2_U2638); 
assign P2_R1957_U117 = ~(P2_R1957_U96 & P2_R1957_U75); 
assign P2_R1957_U153 = ~(P2_R1957_U96 & P2_R1957_U75); 
assign P2_ADD_394_U72 = ~(P2_ADD_394_U146 & P2_ADD_394_U145); 
assign P2_ADD_394_U113 = ~P2_ADD_394_U38; 
assign P2_ADD_394_U165 = ~(P2_ADD_394_U38 & P2_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P2_R2267_U56 = P2_R2267_U136 & P2_R2267_U135; 
assign P2_R2267_U93 = ~P2_R2267_U30; 
assign P2_R2267_U95 = ~(P2_U2788 & P2_R2267_U94); 
assign P2_R2267_U165 = ~(P2_U2787 & P2_R2267_U30); 
assign P1_R2027_U58 = ~(P1_R2027_U156 & P1_R2027_U155); 
assign P1_R2144_U49 = ~(P1_R2144_U239 & P1_R2144_U238); 
assign P1_R2144_U99 = ~(P1_R2144_U53 & P1_R2144_U84); 
assign P1_R2144_U119 = ~P1_R2144_U84; 
assign P1_R2144_U123 = ~P1_R2144_U83; 
assign P1_R2144_U124 = ~(P1_R2144_U83 & P1_R2144_U105); 
assign P1_R2144_U136 = ~(P1_R2144_U62 & P1_R2144_U135); 
assign P1_R2144_U215 = ~(P1_R2144_U59 & P1_R2144_U160 & P1_R2144_U81); 
assign P1_R2144_U216 = ~(P1_R2144_U149 & P1_R2144_U83); 
assign P1_R2144_U218 = ~(P1_R2144_U150 & P1_R2144_U84); 
assign P1_R2278_U99 = ~(P1_R2278_U610 & P1_R2278_U609); 
assign P1_R2278_U556 = ~(P1_R2278_U232 & P1_R2278_U31); 
assign P1_R2358_U29 = ~P1_U2649; 
assign P1_R2358_U163 = ~P1_U2666; 
assign P1_R2358_U206 = ~(P1_U2649 & P1_R2358_U427); 
assign P1_R2358_U208 = ~(P1_R2358_U434 & P1_R2358_U433 & P1_R2358_U31); 
assign P1_R2358_U210 = ~(P1_R2358_U209 & P1_R2358_U23); 
assign P1_R2358_U488 = ~(P1_U2666 & P1_R2358_U23); 
assign P1_R2358_U500 = ~(P1_U2666 & P1_R2358_U23); 
assign P1_R584_U6 = ~P1_U2676; 
assign P1_R584_U7 = ~P1_U2677; 
assign P1_R584_U8 = ~P1_U2674; 
assign P1_R584_U9 = ~P1_U2675; 
assign P1_R2099_U79 = ~(P1_R2099_U332 & P1_R2099_U331); 
assign P1_R2099_U80 = ~(P1_R2099_U334 & P1_R2099_U333); 
assign P1_R2099_U168 = ~P1_R2099_U141; 
assign P1_R2099_U169 = ~P1_R2099_U14; 
assign P1_R2099_U328 = ~(P1_R2099_U55 & P1_R2099_U14); 
assign P1_R2099_U330 = ~(P1_R2099_U57 & P1_R2099_U141); 
assign P1_R2337_U83 = ~(P1_R2337_U166 & P1_R2337_U165); 
assign P1_R2337_U110 = ~P1_R2337_U38; 
assign P1_R2337_U163 = ~(P1_R2337_U38 & P1_PHYADDRPOINTER_REG_19__SCAN_IN); 
assign P1_LT_563_1260_U7 = ~P1_U2673; 
assign P1_R2096_U83 = ~(P1_R2096_U166 & P1_R2096_U165); 
assign P1_R2096_U110 = ~P1_R2096_U38; 
assign P1_R2096_U163 = ~(P1_R2096_U38 & P1_REIP_REG_19__SCAN_IN); 
assign P1_LT_563_U14 = P1_LT_563_U24 & P1_LT_563_U25; 
assign P1_LT_563_U20 = ~(P1_LT_563_U28 & P1_LT_563_U19 & P1_LT_563_U18 & P1_LT_563_U17); 
assign P1_ADD_405_U72 = ~(P1_ADD_405_U146 & P1_ADD_405_U145); 
assign P1_ADD_405_U113 = ~P1_ADD_405_U38; 
assign P1_ADD_405_U165 = ~(P1_ADD_405_U38 & P1_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P1_ADD_515_U72 = ~(P1_ADD_515_U144 & P1_ADD_515_U143); 
assign P1_ADD_515_U110 = ~P1_ADD_515_U38; 
assign P1_ADD_515_U163 = ~(P1_ADD_515_U38 & P1_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_U3767 = P3_U3766 & P3_U3765 & P3_U5867; 
assign P3_U3768 = P3_U3769 & P3_U5873; 
assign P3_U3774 = P3_U3773 & P3_U3772 & P3_U5891; 
assign P3_U3775 = P3_U3776 & P3_U5897; 
assign P3_U3963 = P3_U6482 & P3_U6481 & P3_U6484 & P3_U6483; 
assign P3_U3964 = P3_U6490 & P3_U6489 & P3_U6492 & P3_U6491; 
assign P3_U5846 = ~(P3_U4318 & P3_U5844); 
assign P3_U5915 = ~(P3_ADD_371_1212_U86 & P3_U2360); 
assign P3_U5920 = ~(P3_ADD_360_1242_U5 & P3_U2395); 
assign P3_U5945 = ~(P3_SUB_357_1258_U15 & P3_U2393); 
assign P3_U6042 = ~(P3_ADD_558_U88 & P3_U3220); 
assign P3_U6043 = ~(P3_ADD_553_U88 & P3_U4298); 
assign P3_U6044 = ~(P3_ADD_547_U88 & P3_U4299); 
assign P3_U6047 = ~(P3_ADD_531_U88 & P3_U2354); 
assign P3_U6055 = ~(P3_ADD_385_U88 & P3_U2358); 
assign P3_U6056 = ~(P3_ADD_380_U88 & P3_U2359); 
assign P3_U6057 = ~(P3_ADD_349_U88 & P3_U4306); 
assign P3_U6058 = ~(P3_ADD_344_U88 & P3_U2362); 
assign P3_U6069 = ~(P3_ADD_541_U83 & P3_U4300); 
assign P3_U6070 = ~(P3_ADD_536_U83 & P3_U4301); 
assign P3_U6073 = ~(P3_ADD_515_U83 & P3_U4302); 
assign P3_U6074 = ~(P3_ADD_494_U83 & P3_U2356); 
assign P3_U6075 = ~(P3_ADD_476_U83 & P3_U4303); 
assign P3_U6076 = ~(P3_ADD_441_U83 & P3_U4304); 
assign P3_U6077 = ~(P3_ADD_405_U83 & P3_U4305); 
assign P3_U6078 = ~(P3_ADD_394_U83 & P3_U2357); 
assign P3_U6384 = ~(P3_ADD_526_U58 & P3_U2355); 
assign P3_U6499 = ~(P3_U2387 & P3_ADD_371_1212_U86); 
assign P3_U6503 = ~(P3_U2396 & P3_ADD_360_1242_U5); 
assign P3_U6512 = ~(P3_U2394 & P3_SUB_357_1258_U15); 
assign P3_U6549 = ~(P3_ADD_318_U83 & P3_U2398); 
assign P3_U6554 = ~(P3_ADD_339_U83 & P3_U2388); 
assign P3_U6558 = ~(P3_ADD_315_U79 & P3_U2397); 
assign P3_U6994 = ~(P3_ADD_546_U58 & P3_U2400); 
assign P3_U7091 = ~(P3_ADD_552_U58 & P3_U2399); 
assign P3_U7254 = ~(P3_ADD_467_U83 & P3_U2601); 
assign P3_U7256 = ~(P3_ADD_430_U83 & P3_U2405); 
assign P2_U2460 = P2_R2182_U40 & P2_U3317; 
assign P2_U2463 = P2_U4637 & P2_U2462; 
assign P2_U2469 = P2_U4633 & P2_U2462; 
assign P2_U2472 = P2_U4634 & P2_U2462; 
assign P2_U2477 = P2_U2476 & P2_U2462; 
assign P2_U2502 = P2_U2501 & P2_U4637; 
assign P2_U2506 = P2_U2501 & P2_U4633; 
assign P2_U2508 = P2_U2501 & P2_U4634; 
assign P2_U2510 = P2_U2501 & P2_U2476; 
assign P2_U3306 = ~(P2_U4656 & P2_U3284); 
assign P2_U3622 = ~(P2_U8298 & P2_U8297); 
assign P2_U3623 = ~(P2_U8300 & P2_U8299); 
assign P2_U3624 = ~(P2_U8302 & P2_U8301); 
assign P2_U3625 = ~(P2_U8304 & P2_U8303); 
assign P2_U3626 = ~(P2_U8306 & P2_U8305); 
assign P2_U3627 = ~(P2_U8308 & P2_U8307); 
assign P2_U3628 = ~(P2_U8310 & P2_U8309); 
assign P2_U3629 = ~(P2_U8312 & P2_U8311); 
assign P2_U3871 = P2_U8071 & P2_U8070 & P2_U3870 & P2_U2512; 
assign P2_U3891 = P2_U5649 & P2_U5650; 
assign P2_U4393 = P2_U8055 & P2_U8054; 
assign P2_U4397 = P2_U8120 & P2_U8119; 
assign P2_U4404 = P2_U8146 & P2_U8145; 
assign P2_U4462 = ~(P2_U2374 & P2_U6568); 
assign P2_U4630 = ~(P2_U3719 & P2_U4469); 
assign P2_U4638 = ~P2_U3378; 
assign P2_U4657 = ~(P2_U4637 & P2_U2462); 
assign P2_U4715 = ~(P2_U4633 & P2_U2462); 
assign P2_U4767 = ~P2_U3353; 
assign P2_U4774 = ~(P2_U4634 & P2_U2462); 
assign P2_U4831 = ~(P2_U2476 & P2_U2462); 
assign P2_U5347 = ~(P2_U2501 & P2_U4637); 
assign P2_U5404 = ~(P2_U2501 & P2_U4633); 
assign P2_U5462 = ~(P2_U2501 & P2_U4634); 
assign P2_U5519 = ~(P2_U2501 & P2_U2476); 
assign P2_U5612 = ~(P2_R2182_U76 & P2_U4469); 
assign P2_U5621 = ~(P2_R2182_U40 & P2_U4469); 
assign P2_U5631 = ~(P2_R2182_U68 & P2_U4469); 
assign P2_U5638 = ~(P2_R2182_U69 & P2_U4469); 
assign P2_U5645 = ~(P2_U4636 & P2_U3579); 
assign P2_U5656 = ~(P2_U3338 & P2_U3353); 
assign P2_U6230 = ~(P2_U4411 & P2_U6229); 
assign P2_U6326 = ~(P2_U2513 & P2_U3254); 
assign P2_U6470 = ~(P2_U3578 & P2_U6469); 
assign P2_U8064 = ~P2_U3579; 
assign P2_U8108 = ~(P2_U3579 & P2_U3319); 
assign P2_U8314 = ~(P2_U3242 & P2_R2267_U56); 
assign P2_U8399 = ~(P2_R2337_U81 & P2_U3284); 
assign P1_U2604 = P1_U2379 & P1_EBX_REG_31__SCAN_IN; 
assign P1_U2665 = ~(P1_U6833 & P1_U4024); 
assign P1_U3311 = ~P1_R2144_U49; 
assign P1_U3332 = ~(P1_U3325 & P1_U3331); 
assign P1_U3765 = P1_U5575 & P1_U5576; 
assign P1_U3769 = P1_U5582 & P1_U5583; 
assign P1_U3773 = P1_U5589 & P1_U5590; 
assign P1_U3777 = P1_U5596 & P1_U5597; 
assign P1_U3779 = P1_U5603 & P1_U5604; 
assign P1_U3782 = P1_U5610 & P1_U5611; 
assign P1_U3785 = P1_U5617 & P1_U5618; 
assign P1_U3788 = P1_U5624 & P1_U5625; 
assign P1_U3791 = P1_U5631 & P1_U5632; 
assign P1_U3794 = P1_U5638 & P1_U5639; 
assign P1_U3797 = P1_U5645 & P1_U5646; 
assign P1_U3800 = P1_U5652 & P1_U5653; 
assign P1_U3803 = P1_U5659 & P1_U5660; 
assign P1_U3806 = P1_U5666 & P1_U5667; 
assign P1_U3809 = P1_U5673 & P1_U5674; 
assign P1_U3812 = P1_U5680 & P1_U5681; 
assign P1_U3815 = P1_U5687 & P1_U5688; 
assign P1_U3818 = P1_U5694 & P1_U5695; 
assign P1_U3821 = P1_U5701 & P1_U5702; 
assign P1_U3824 = P1_U5708 & P1_U5709; 
assign P1_U3827 = P1_U5715 & P1_U5716; 
assign P1_U3830 = P1_U5722 & P1_U5723; 
assign P1_U3833 = P1_U5729 & P1_U5730; 
assign P1_U3836 = P1_U5736 & P1_U5737; 
assign P1_U3839 = P1_U5743 & P1_U5744; 
assign P1_U3842 = P1_U5750 & P1_U5751; 
assign P1_U3845 = P1_U5757 & P1_U5758; 
assign P1_U3848 = P1_U5764 & P1_U5765; 
assign P1_U3851 = P1_U5771 & P1_U5772; 
assign P1_U3854 = P1_U5778 & P1_U5779; 
assign P1_U3857 = P1_U5785 & P1_U5786; 
assign P1_U3860 = P1_U5792 & P1_U5793; 
assign P1_U4525 = ~P1_U3331; 
assign P1_U5548 = ~(P1_U4226 & P1_R2144_U49); 
assign P1_U5570 = ~(P1_R2099_U86 & P1_U2380); 
assign P1_U5571 = ~(P1_R2027_U5 & P1_U2378); 
assign P1_U5572 = ~(P1_R2278_U99 & P1_U2377); 
assign P1_U5573 = ~(P1_ADD_405_U4 & P1_U2375); 
assign P1_U5574 = ~(P1_U2374 & P1_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P1_U5577 = ~(P1_R2099_U87 & P1_U2380); 
assign P1_U5578 = ~(P1_R2027_U71 & P1_U2378); 
assign P1_U5580 = ~(P1_ADD_405_U85 & P1_U2375); 
assign P1_U5581 = ~(P1_ADD_515_U4 & P1_U2374); 
assign P1_U5584 = ~(P1_R2099_U138 & P1_U2380); 
assign P1_U5585 = ~(P1_R2027_U60 & P1_U2378); 
assign P1_U5587 = ~(P1_ADD_405_U5 & P1_U2375); 
assign P1_U5588 = ~(P1_ADD_515_U67 & P1_U2374); 
assign P1_U5591 = ~(P1_R2099_U42 & P1_U2380); 
assign P1_U5592 = ~(P1_R2027_U57 & P1_U2378); 
assign P1_U5594 = ~(P1_ADD_405_U95 & P1_U2375); 
assign P1_U5595 = ~(P1_ADD_515_U85 & P1_U2374); 
assign P1_U5598 = ~(P1_R2099_U41 & P1_U2380); 
assign P1_U5599 = ~(P1_R2027_U56 & P1_U2378); 
assign P1_U5601 = ~(P1_ADD_405_U76 & P1_U2375); 
assign P1_U5602 = ~(P1_ADD_515_U76 & P1_U2374); 
assign P1_U5605 = ~(P1_R2099_U40 & P1_U2380); 
assign P1_U5606 = ~(P1_R2027_U55 & P1_U2378); 
assign P1_U5608 = ~(P1_ADD_405_U79 & P1_U2375); 
assign P1_U5609 = ~(P1_ADD_515_U79 & P1_U2374); 
assign P1_U5612 = ~(P1_R2099_U39 & P1_U2380); 
assign P1_U5613 = ~(P1_R2027_U54 & P1_U2378); 
assign P1_U5615 = ~(P1_ADD_405_U63 & P1_U2375); 
assign P1_U5616 = ~(P1_ADD_515_U62 & P1_U2374); 
assign P1_U5619 = ~(P1_R2099_U38 & P1_U2380); 
assign P1_U5620 = ~(P1_R2027_U53 & P1_U2378); 
assign P1_U5622 = ~(P1_ADD_405_U89 & P1_U2375); 
assign P1_U5623 = ~(P1_ADD_515_U89 & P1_U2374); 
assign P1_U5626 = ~(P1_R2099_U37 & P1_U2380); 
assign P1_U5627 = ~(P1_R2027_U52 & P1_U2378); 
assign P1_U5629 = ~(P1_ADD_405_U80 & P1_U2375); 
assign P1_U5630 = ~(P1_ADD_515_U80 & P1_U2374); 
assign P1_U5633 = ~(P1_R2099_U36 & P1_U2380); 
assign P1_U5634 = ~(P1_R2027_U51 & P1_U2378); 
assign P1_U5636 = ~(P1_ADD_405_U70 & P1_U2375); 
assign P1_U5637 = ~(P1_ADD_515_U70 & P1_U2374); 
assign P1_U5640 = ~(P1_R2099_U85 & P1_U2380); 
assign P1_U5641 = ~(P1_R2027_U81 & P1_U2378); 
assign P1_U5643 = ~(P1_ADD_405_U83 & P1_U2375); 
assign P1_U5644 = ~(P1_ADD_515_U83 & P1_U2374); 
assign P1_U5647 = ~(P1_R2099_U84 & P1_U2380); 
assign P1_U5648 = ~(P1_R2027_U80 & P1_U2378); 
assign P1_U5650 = ~(P1_ADD_405_U73 & P1_U2375); 
assign P1_U5651 = ~(P1_ADD_515_U73 & P1_U2374); 
assign P1_U5654 = ~(P1_R2099_U83 & P1_U2380); 
assign P1_U5655 = ~(P1_R2027_U79 & P1_U2378); 
assign P1_U5657 = ~(P1_ADD_405_U88 & P1_U2375); 
assign P1_U5658 = ~(P1_ADD_515_U88 & P1_U2374); 
assign P1_U5661 = ~(P1_R2099_U82 & P1_U2380); 
assign P1_U5662 = ~(P1_R2027_U78 & P1_U2378); 
assign P1_U5664 = ~(P1_ADD_405_U69 & P1_U2375); 
assign P1_U5665 = ~(P1_ADD_515_U69 & P1_U2374); 
assign P1_U5668 = ~(P1_R2099_U81 & P1_U2380); 
assign P1_U5669 = ~(P1_R2027_U77 & P1_U2378); 
assign P1_U5671 = ~(P1_ADD_405_U78 & P1_U2375); 
assign P1_U5672 = ~(P1_ADD_515_U78 & P1_U2374); 
assign P1_U5675 = ~(P1_R2099_U80 & P1_U2380); 
assign P1_U5676 = ~(P1_R2027_U76 & P1_U2378); 
assign P1_U5678 = ~(P1_ADD_405_U75 & P1_U2375); 
assign P1_U5679 = ~(P1_ADD_515_U75 & P1_U2374); 
assign P1_U5682 = ~(P1_R2099_U79 & P1_U2380); 
assign P1_U5683 = ~(P1_R2027_U75 & P1_U2378); 
assign P1_U5685 = ~(P1_ADD_405_U91 & P1_U2375); 
assign P1_U5686 = ~(P1_ADD_515_U91 & P1_U2374); 
assign P1_U5690 = ~(P1_R2027_U74 & P1_U2378); 
assign P1_U5692 = ~(P1_ADD_405_U67 & P1_U2375); 
assign P1_U5693 = ~(P1_ADD_515_U66 & P1_U2374); 
assign P1_U5697 = ~(P1_R2027_U73 & P1_U2378); 
assign P1_U5699 = ~(P1_ADD_405_U72 & P1_U2375); 
assign P1_U5700 = ~(P1_ADD_515_U72 & P1_U2374); 
assign P1_U5704 = ~(P1_R2027_U72 & P1_U2378); 
assign P1_U5711 = ~(P1_R2027_U70 & P1_U2378); 
assign P1_U5718 = ~(P1_R2027_U69 & P1_U2378); 
assign P1_U5725 = ~(P1_R2027_U68 & P1_U2378); 
assign P1_U5732 = ~(P1_R2027_U67 & P1_U2378); 
assign P1_U5739 = ~(P1_R2027_U66 & P1_U2378); 
assign P1_U5746 = ~(P1_R2027_U65 & P1_U2378); 
assign P1_U5753 = ~(P1_R2027_U64 & P1_U2378); 
assign P1_U5760 = ~(P1_R2027_U63 & P1_U2378); 
assign P1_U5767 = ~(P1_R2027_U62 & P1_U2378); 
assign P1_U5774 = ~(P1_R2027_U61 & P1_U2378); 
assign P1_U5781 = ~(P1_R2027_U59 & P1_U2378); 
assign P1_U5788 = ~(P1_R2027_U58 & P1_U2378); 
assign P1_U5800 = ~(P1_U2372 & P1_R2278_U99); 
assign P1_U5889 = ~(P1_R2337_U83 & P1_U2376); 
assign P1_U6311 = ~(P1_U2371 & P1_R2099_U80); 
assign P1_U6314 = ~(P1_U2371 & P1_R2099_U79); 
assign P1_U6832 = ~(P1_R2337_U83 & P1_U2352); 
assign P1_U6869 = ~(P1_R2144_U49 & P1_U6746); 
assign P1_U6883 = ~(P1_U4159 & P1_R2144_U49); 
assign P1_U7481 = ~(P1_U2379 & P1_U3429); 
assign P1_U7482 = ~(P1_U2369 & P1_U6367); 
assign P1_U7483 = ~(P1_U3888 & P1_U2369); 
assign P1_U7691 = ~(P1_R2144_U49 & P1_U3313); 
assign P3_ADD_476_U40 = ~(P3_ADD_476_U110 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_476_U164 = ~(P3_ADD_476_U110 & P3_ADD_476_U39); 
assign P3_ADD_531_U41 = ~(P3_ADD_531_U114 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_531_U173 = ~(P3_ADD_531_U114 & P3_ADD_531_U40); 
assign P3_SUB_320_U45 = ~P3_ADD_318_U83; 
assign P3_SUB_320_U76 = P3_SUB_320_U153 & P3_SUB_320_U152; 
assign P3_SUB_320_U118 = ~(P3_ADD_318_U83 & P3_SUB_320_U117); 
assign P3_ADD_318_U40 = ~(P3_ADD_318_U110 & P3_PHYADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_318_U164 = ~(P3_ADD_318_U110 & P3_ADD_318_U39); 
assign P3_ADD_315_U40 = ~(P3_ADD_315_U107 & P3_PHYADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_315_U156 = ~(P3_ADD_315_U107 & P3_ADD_315_U39); 
assign P3_ADD_360_1242_U6 = P3_ADD_360_1242_U182 & P3_ADD_360_1242_U76; 
assign P3_ADD_360_1242_U155 = ~P3_ADD_360_1242_U76; 
assign P3_ADD_360_1242_U156 = ~P3_ADD_360_1242_U50; 
assign P3_ADD_360_1242_U251 = ~(P3_ADD_360_1242_U50 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_360_1242_U253 = ~(P3_ADD_360_1242_U76 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_467_U40 = ~(P3_ADD_467_U110 & P3_REIP_REG_19__SCAN_IN); 
assign P3_ADD_467_U164 = ~(P3_ADD_467_U110 & P3_ADD_467_U39); 
assign P3_ADD_430_U40 = ~(P3_ADD_430_U110 & P3_REIP_REG_19__SCAN_IN); 
assign P3_ADD_430_U164 = ~(P3_ADD_430_U110 & P3_ADD_430_U39); 
assign P3_ADD_380_U41 = ~(P3_ADD_380_U114 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_380_U173 = ~(P3_ADD_380_U114 & P3_ADD_380_U40); 
assign P3_ADD_344_U41 = ~(P3_ADD_344_U114 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_344_U173 = ~(P3_ADD_344_U114 & P3_ADD_344_U40); 
assign P3_LT_563_U27 = ~(P3_LT_563_U25 & P3_LT_563_U26 & P3_LT_563_U24); 
assign P3_ADD_339_U40 = ~(P3_ADD_339_U110 & P3_PHYADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_339_U164 = ~(P3_ADD_339_U110 & P3_ADD_339_U39); 
assign P3_ADD_541_U40 = ~(P3_ADD_541_U110 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_541_U164 = ~(P3_ADD_541_U110 & P3_ADD_541_U39); 
assign P3_SUB_357_1258_U89 = ~(P3_SUB_357_1258_U456 & P3_SUB_357_1258_U455); 
assign P3_SUB_357_1258_U200 = ~P3_SUB_357_1258_U143; 
assign P3_SUB_357_1258_U201 = ~(P3_SUB_357_1258_U101 & P3_SUB_357_1258_U143); 
assign P3_SUB_357_1258_U202 = ~P3_SUB_357_1258_U67; 
assign P3_SUB_357_1258_U247 = ~(P3_SUB_357_1258_U143 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_SUB_357_1258_U272 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U67); 
assign P3_SUB_357_1258_U448 = ~(P3_SUB_357_1258_U142 & P3_SUB_357_1258_U143); 
assign P3_ADD_515_U40 = ~(P3_ADD_515_U110 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_515_U164 = ~(P3_ADD_515_U110 & P3_ADD_515_U39); 
assign P3_ADD_394_U40 = ~(P3_ADD_394_U113 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_394_U168 = ~(P3_ADD_394_U113 & P3_ADD_394_U39); 
assign P3_ADD_441_U40 = ~(P3_ADD_441_U110 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_441_U164 = ~(P3_ADD_441_U110 & P3_ADD_441_U39); 
assign P3_ADD_349_U41 = ~(P3_ADD_349_U114 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_349_U173 = ~(P3_ADD_349_U114 & P3_ADD_349_U40); 
assign P3_ADD_405_U40 = ~(P3_ADD_405_U113 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_405_U168 = ~(P3_ADD_405_U113 & P3_ADD_405_U39); 
assign P3_ADD_553_U41 = ~(P3_ADD_553_U114 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_553_U173 = ~(P3_ADD_553_U114 & P3_ADD_553_U40); 
assign P3_ADD_558_U41 = ~(P3_ADD_558_U114 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_558_U173 = ~(P3_ADD_558_U114 & P3_ADD_558_U40); 
assign P3_ADD_385_U41 = ~(P3_ADD_385_U114 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_385_U173 = ~(P3_ADD_385_U114 & P3_ADD_385_U40); 
assign P3_ADD_547_U41 = ~(P3_ADD_547_U114 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_547_U173 = ~(P3_ADD_547_U114 & P3_ADD_547_U40); 
assign P3_ADD_371_1212_U6 = P3_ADD_371_1212_U194 & P3_ADD_371_1212_U49; 
assign P3_ADD_371_1212_U53 = ~(P3_ADD_371_1212_U163 & P3_ADD_371_1212_U101); 
assign P3_ADD_371_1212_U78 = ~(P3_ADD_371_1212_U163 & P3_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P3_ADD_494_U40 = ~(P3_ADD_494_U110 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_494_U164 = ~(P3_ADD_494_U110 & P3_ADD_494_U39); 
assign P3_ADD_536_U40 = ~(P3_ADD_536_U110 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_536_U164 = ~(P3_ADD_536_U110 & P3_ADD_536_U39); 
assign P2_R2099_U68 = ~(P2_R2099_U152 & P2_R2099_U151); 
assign P2_R2099_U124 = ~P2_R2099_U24; 
assign P2_R2099_U149 = ~(P2_U2738 & P2_R2099_U24); 
assign P2_ADD_391_1196_U28 = ~P2_R2182_U75; 
assign P2_ADD_391_1196_U49 = ~P2_R2096_U97; 
assign P2_ADD_391_1196_U169 = ~P2_ADD_391_1196_U118; 
assign P2_ADD_391_1196_U171 = ~(P2_ADD_391_1196_U170 & P2_ADD_391_1196_U118); 
assign P2_ADD_391_1196_U174 = P2_R2182_U75 | P2_R2096_U74; 
assign P2_ADD_391_1196_U176 = ~(P2_R2096_U74 & P2_R2182_U75); 
assign P2_ADD_391_1196_U326 = ~(P2_R2182_U75 & P2_ADD_391_1196_U29); 
assign P2_ADD_391_1196_U328 = ~(P2_R2182_U75 & P2_ADD_391_1196_U29); 
assign P2_ADD_391_1196_U332 = ~(P2_R2096_U75 & P2_ADD_391_1196_U26); 
assign P2_ADD_391_1196_U334 = ~(P2_R2096_U75 & P2_ADD_391_1196_U26); 
assign P2_ADD_391_1196_U349 = ~(P2_ADD_391_1196_U122 & P2_ADD_391_1196_U123); 
assign P2_ADD_391_1196_U350 = ~(P2_ADD_391_1196_U165 & P2_ADD_391_1196_U348); 
assign P2_R2182_U9 = P2_U2675 & P2_R2182_U21; 
assign P2_R2182_U137 = ~P2_R2182_U21; 
assign P2_R2182_U199 = ~(P2_R2182_U22 & P2_R2182_U21); 
assign P2_R2182_U202 = ~(P2_R2182_U136 & P2_U2676); 
assign P2_R2027_U41 = ~(P2_R2027_U114 & P2_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P2_R2027_U173 = ~(P2_R2027_U114 & P2_R2027_U40); 
assign P2_R2337_U41 = ~(P2_R2337_U111 & P2_PHYADDRPOINTER_REG_20__SCAN_IN); 
assign P2_R2337_U162 = ~(P2_R2337_U111 & P2_R2337_U40); 
assign P2_R2096_U21 = P2_U2636 & P2_R2096_U20; 
assign P2_R2096_U96 = ~(P2_R2096_U261 & P2_R2096_U260); 
assign P2_R2096_U148 = ~P2_R2096_U20; 
assign P2_R2096_U256 = ~(P2_R2096_U32 & P2_R2096_U20); 
assign P2_R2096_U259 = ~(P2_R2096_U147 & P2_U2637); 
assign P2_R1957_U44 = ~P2_U3673; 
assign P2_R1957_U76 = P2_R1957_U153 & P2_R1957_U152; 
assign P2_R1957_U118 = ~(P2_U3673 & P2_R1957_U117); 
assign P2_ADD_394_U40 = ~(P2_ADD_394_U113 & P2_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P2_ADD_394_U166 = ~(P2_ADD_394_U113 & P2_ADD_394_U39); 
assign P2_R2267_U20 = P2_R2267_U95 & P2_R2267_U30; 
assign P2_R2267_U31 = ~(P2_R2267_U45 & P2_R2267_U93); 
assign P2_R2267_U132 = ~(P2_R2267_U93 & P2_R2267_U86); 
assign P2_R2267_U166 = ~(P2_R2267_U93 & P2_R2267_U86); 
assign P1_R2144_U8 = P1_R2144_U138 & P1_R2144_U136; 
assign P1_R2144_U79 = ~(P1_R2144_U99 & P1_R2144_U54); 
assign P1_R2144_U82 = P1_R2144_U215 & P1_R2144_U214; 
assign P1_R2144_U125 = ~(P1_R2144_U21 & P1_R2144_U124); 
assign P1_R2144_U127 = ~(P1_R2144_U60 & P1_R2144_U124); 
assign P1_R2144_U212 = ~(P1_R2144_U57 & P1_R2144_U124 & P1_R2144_U23); 
assign P1_R2144_U217 = ~(P1_R2144_U44 & P1_R2144_U123); 
assign P1_R2144_U219 = ~(P1_R2144_U46 & P1_R2144_U119); 
assign P1_R2278_U33 = ~P1_U2799; 
assign P1_R2278_U213 = ~(P1_U2799 & P1_R2278_U232); 
assign P1_R2278_U557 = ~(P1_R2278_U556 & P1_R2278_U555); 
assign P1_R2278_U558 = ~(P1_U2799 & P1_R2278_U32 & P1_R2278_U31); 
assign P1_R2358_U200 = ~(P1_R2358_U209 & P1_R2358_U208); 
assign P1_R2358_U205 = ~(P1_R2358_U432 & P1_R2358_U431 & P1_R2358_U29); 
assign P1_R2358_U246 = ~(P1_U2352 & P1_R2358_U208); 
assign P1_R2358_U487 = ~(P1_U2352 & P1_R2358_U163); 
assign P1_R2358_U499 = ~(P1_U2352 & P1_R2358_U163); 
assign P1_LT_589_U7 = P1_R584_U7 & P1_R584_U6; 
assign P1_R2099_U15 = ~(P1_R2099_U169 & P1_R2099_U55); 
assign P1_R2099_U327 = ~(P1_R2099_U258 & P1_R2099_U169); 
assign P1_R2099_U329 = ~(P1_R2099_U168 & P1_R2099_U282); 
assign P1_R2337_U40 = ~(P1_R2337_U110 & P1_PHYADDRPOINTER_REG_19__SCAN_IN); 
assign P1_R2337_U164 = ~(P1_R2337_U110 & P1_R2337_U39); 
assign P1_LT_563_1260_U8 = ~(P1_R584_U8 & P1_LT_563_1260_U7); 
assign P1_LT_563_1260_U9 = ~(P1_R584_U9 & P1_LT_563_1260_U7); 
assign P1_R2096_U40 = ~(P1_R2096_U110 & P1_REIP_REG_19__SCAN_IN); 
assign P1_R2096_U164 = ~(P1_R2096_U110 & P1_R2096_U39); 
assign P1_LT_563_U23 = ~(P1_LT_563_U13 & P1_LT_563_U20); 
assign P1_ADD_405_U40 = ~(P1_ADD_405_U113 & P1_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P1_ADD_405_U166 = ~(P1_ADD_405_U113 & P1_ADD_405_U39); 
assign P1_ADD_515_U40 = ~(P1_ADD_515_U110 & P1_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P1_ADD_515_U164 = ~(P1_ADD_515_U110 & P1_ADD_515_U39); 
assign P3_U2672 = ~(P3_U7092 & P3_U7091); 
assign P3_U2704 = ~(P3_U6995 & P3_U6993 & P3_U6994); 
assign P3_U2820 = ~(P3_U6486 & P3_U6485 & P3_U6487 & P3_U6488 & P3_U3964); 
assign P3_U2821 = ~(P3_U6478 & P3_U6477 & P3_U6480 & P3_U6479 & P3_U3963); 
assign P3_U2854 = ~(P3_U5847 & P3_U5845 & P3_U5846); 
assign P3_U3781 = P3_U3780 & P3_U3779 & P3_U5915; 
assign P3_U3782 = P3_U3783 & P3_U5920; 
assign P3_U3819 = P3_U6044 & P3_U6043; 
assign P3_U3823 = P3_U6058 & P3_U6057 & P3_U6056 & P3_U6055; 
assign P3_U3827 = P3_U6073 & P3_U6072; 
assign P3_U3829 = P3_U6075 & P3_U6074 & P3_U6076 & P3_U6078 & P3_U6077; 
assign P3_U3965 = P3_U6498 & P3_U6497 & P3_U6500 & P3_U6499; 
assign P3_U4093 = P3_U7253 & P3_U4316 & P3_U7254; 
assign P3_U5868 = ~(P3_U3764 & P3_U5850 & P3_U5849 & P3_U3761 & P3_U3767); 
assign P3_U5892 = ~(P3_U5874 & P3_U3771 & P3_U5872 & P3_U3774 & P3_U3768); 
assign P3_U5939 = ~(P3_ADD_371_1212_U6 & P3_U2360); 
assign P3_U5944 = ~(P3_ADD_360_1242_U6 & P3_U2395); 
assign P3_U5993 = ~(P3_SUB_357_1258_U89 & P3_U2393); 
assign P3_U6507 = ~(P3_U2387 & P3_ADD_371_1212_U6); 
assign P3_U6511 = ~(P3_U2396 & P3_ADD_360_1242_U6); 
assign P3_U6528 = ~(P3_U2394 & P3_SUB_357_1258_U89); 
assign P2_U2459 = P2_U8053 & P2_U8052 & P2_U4393; 
assign P2_U2482 = P2_U4638 & P2_U4637; 
assign P2_U2485 = P2_U4638 & P2_U4633; 
assign P2_U2487 = P2_U4638 & P2_U4634; 
assign P2_U2489 = P2_U4638 & P2_U2476; 
assign P2_U2494 = P2_U4633 & P2_U2460; 
assign P2_U2496 = P2_U4634 & P2_U2460; 
assign P2_U2498 = P2_U2476 & P2_U2460; 
assign P2_U2812 = P2_U3242 & P2_R2267_U20; 
assign P2_U3425 = ~(P2_U2460 & P2_U4637); 
assign P2_U3541 = ~(P2_U6231 & P2_U6230); 
assign P2_U3542 = ~(P2_U2374 & P2_U6326); 
assign P2_U3543 = ~(P2_U2374 & P2_U6470); 
assign P2_U3546 = ~(P2_U4069 & P2_U4462); 
assign P2_U3672 = ~(P2_U8400 & P2_U8399); 
assign P2_U4402 = ~(P2_U4462 & P2_U4188); 
assign P2_U4403 = ~(P2_U3534 & P2_U4462); 
assign P2_U4406 = ~(P2_U2513 & P2_U3871); 
assign P2_U4443 = ~P2_U3306; 
assign P2_U4889 = ~(P2_U4638 & P2_U4637); 
assign P2_U4946 = ~(P2_U4638 & P2_U4633); 
assign P2_U5004 = ~(P2_U4638 & P2_U4634); 
assign P2_U5061 = ~(P2_U4638 & P2_U2476); 
assign P2_U5174 = ~(P2_U4633 & P2_U2460); 
assign P2_U5232 = ~(P2_U4634 & P2_U2460); 
assign P2_U5289 = ~(P2_U2476 & P2_U2460); 
assign P2_U5614 = ~(P2_U5613 & P2_U5612); 
assign P2_U5657 = ~(P2_U2398 & P2_U5656); 
assign P2_U6859 = ~(P2_U4421 & P2_U4468 & P2_U4404); 
assign P2_U8107 = ~(P2_U8064 & P2_U4636); 
assign P1_U2476 = P1_R2144_U8 & P1_R2144_U49; 
assign P1_U2508 = ~(P1_R2144_U49 | P1_R2144_U8); 
assign P1_U2647 = P1_R2144_U8 & P1_U6746; 
assign P1_U2648 = ~(P1_U3440 & P1_U6869); 
assign P1_U2798 = ~(P1_U6884 & P1_U6885 & P1_U6883); 
assign P1_U3312 = ~P1_R2144_U8; 
assign P1_U3314 = ~(P1_U3332 & P1_U3309); 
assign P1_U3326 = ~(P1_R2144_U43 & P1_U3332); 
assign P1_U3342 = ~(P1_R2144_U8 & P1_U3311); 
assign P1_U3752 = P1_U5547 & P1_U5548; 
assign P1_U3763 = P1_U5571 & P1_U5570; 
assign P1_U3764 = P1_U5573 & P1_U5572; 
assign P1_U3766 = P1_U3765 & P1_U5574; 
assign P1_U3767 = P1_U5578 & P1_U5577; 
assign P1_U3770 = P1_U3769 & P1_U5581; 
assign P1_U3771 = P1_U5585 & P1_U5584; 
assign P1_U3774 = P1_U3773 & P1_U5588; 
assign P1_U3775 = P1_U5592 & P1_U5591 & P1_U5594; 
assign P1_U3778 = P1_U5599 & P1_U5598 & P1_U5601; 
assign P1_U3780 = P1_U3779 & P1_U5602; 
assign P1_U3781 = P1_U5606 & P1_U5605 & P1_U5608; 
assign P1_U3783 = P1_U3782 & P1_U5609; 
assign P1_U3784 = P1_U5613 & P1_U5612 & P1_U5615; 
assign P1_U3786 = P1_U3785 & P1_U5616; 
assign P1_U3787 = P1_U5620 & P1_U5619 & P1_U5622; 
assign P1_U3789 = P1_U3788 & P1_U5623; 
assign P1_U3790 = P1_U5627 & P1_U5626 & P1_U5629; 
assign P1_U3792 = P1_U3791 & P1_U5630; 
assign P1_U3793 = P1_U5634 & P1_U5633 & P1_U5636; 
assign P1_U3795 = P1_U3794 & P1_U5637; 
assign P1_U3796 = P1_U5641 & P1_U5640 & P1_U5643; 
assign P1_U3798 = P1_U3797 & P1_U5644; 
assign P1_U3799 = P1_U5648 & P1_U5647 & P1_U5650; 
assign P1_U3801 = P1_U3800 & P1_U5651; 
assign P1_U3802 = P1_U5655 & P1_U5654 & P1_U5657; 
assign P1_U3804 = P1_U3803 & P1_U5658; 
assign P1_U3805 = P1_U5662 & P1_U5664; 
assign P1_U3807 = P1_U3806 & P1_U5665; 
assign P1_U3808 = P1_U5669 & P1_U5671; 
assign P1_U3810 = P1_U3809 & P1_U5672; 
assign P1_U3811 = P1_U5676 & P1_U5678; 
assign P1_U3813 = P1_U3812 & P1_U5679; 
assign P1_U3814 = P1_U5683 & P1_U5685; 
assign P1_U3816 = P1_U3815 & P1_U5686; 
assign P1_U3817 = P1_U5690 & P1_U5692; 
assign P1_U3819 = P1_U3818 & P1_U5693; 
assign P1_U3820 = P1_U5697 & P1_U5699; 
assign P1_U3822 = P1_U3821 & P1_U5700; 
assign P1_U4023 = P1_U6830 & P1_U6831 & P1_U6832; 
assign P1_U4526 = ~P1_U3332; 
assign P1_U4530 = ~(P1_R2144_U8 & P1_U3313); 
assign P1_U5544 = ~(P1_U4226 & P1_R2144_U8); 
assign P1_U6368 = ~(P1_U2604 & P1_R2099_U86); 
assign P1_U6376 = ~(P1_U2604 & P1_R2099_U87); 
assign P1_U6384 = ~(P1_U2604 & P1_R2099_U138); 
assign P1_U6392 = ~(P1_U2604 & P1_R2099_U42); 
assign P1_U6400 = ~(P1_U2604 & P1_R2099_U41); 
assign P1_U6408 = ~(P1_U2604 & P1_R2099_U40); 
assign P1_U6416 = ~(P1_U2604 & P1_R2099_U39); 
assign P1_U6423 = ~(P1_U2604 & P1_R2099_U38); 
assign P1_U6430 = ~(P1_U2604 & P1_R2099_U37); 
assign P1_U6437 = ~(P1_U2604 & P1_R2099_U36); 
assign P1_U6444 = ~(P1_U2604 & P1_R2099_U85); 
assign P1_U6451 = ~(P1_U2604 & P1_R2099_U84); 
assign P1_U6458 = ~(P1_U2604 & P1_R2099_U83); 
assign P1_U6465 = ~(P1_U2604 & P1_R2099_U82); 
assign P1_U6472 = ~(P1_U2604 & P1_R2099_U81); 
assign P1_U6479 = ~(P1_U2604 & P1_R2099_U80); 
assign P1_U6486 = ~(P1_U2604 & P1_R2099_U79); 
assign P1_U6881 = ~(P1_U4159 & P1_R2144_U8); 
assign P1_U7484 = ~(P1_U7481 & P1_U4229 & P1_U7482); 
assign P1_U7485 = ~(P1_U7483 & P1_U4230); 
assign P1_U7692 = ~(P1_U4528 & P1_U3311); 
assign P3_ADD_476_U82 = ~(P3_ADD_476_U164 & P3_ADD_476_U163); 
assign P3_ADD_476_U111 = ~P3_ADD_476_U40; 
assign P3_ADD_476_U161 = ~(P3_ADD_476_U40 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_531_U87 = ~(P3_ADD_531_U173 & P3_ADD_531_U172); 
assign P3_ADD_531_U115 = ~P3_ADD_531_U41; 
assign P3_ADD_531_U170 = ~(P3_ADD_531_U41 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_SUB_320_U32 = ~(P3_SUB_320_U45 & P3_SUB_320_U75 & P3_SUB_320_U96); 
assign P3_ADD_318_U82 = ~(P3_ADD_318_U164 & P3_ADD_318_U163); 
assign P3_ADD_318_U111 = ~P3_ADD_318_U40; 
assign P3_ADD_318_U161 = ~(P3_ADD_318_U40 & P3_PHYADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_315_U78 = ~(P3_ADD_315_U156 & P3_ADD_315_U155); 
assign P3_ADD_315_U108 = ~P3_ADD_315_U40; 
assign P3_ADD_315_U153 = ~(P3_ADD_315_U40 & P3_PHYADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_360_1242_U53 = ~(P3_ADD_360_1242_U100 & P3_ADD_360_1242_U156); 
assign P3_ADD_360_1242_U178 = ~(P3_ADD_360_1242_U156 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_360_1242_U180 = ~(P3_ADD_360_1242_U155 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_360_1242_U252 = ~(P3_ADD_360_1242_U156 & P3_ADD_360_1242_U52); 
assign P3_ADD_360_1242_U254 = ~(P3_ADD_360_1242_U155 & P3_ADD_360_1242_U49); 
assign P3_ADD_467_U82 = ~(P3_ADD_467_U164 & P3_ADD_467_U163); 
assign P3_ADD_467_U111 = ~P3_ADD_467_U40; 
assign P3_ADD_467_U161 = ~(P3_ADD_467_U40 & P3_REIP_REG_20__SCAN_IN); 
assign P3_ADD_430_U82 = ~(P3_ADD_430_U164 & P3_ADD_430_U163); 
assign P3_ADD_430_U111 = ~P3_ADD_430_U40; 
assign P3_ADD_430_U161 = ~(P3_ADD_430_U40 & P3_REIP_REG_20__SCAN_IN); 
assign P3_ADD_380_U87 = ~(P3_ADD_380_U173 & P3_ADD_380_U172); 
assign P3_ADD_380_U115 = ~P3_ADD_380_U41; 
assign P3_ADD_380_U170 = ~(P3_ADD_380_U41 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_344_U87 = ~(P3_ADD_344_U173 & P3_ADD_344_U172); 
assign P3_ADD_344_U115 = ~P3_ADD_344_U41; 
assign P3_ADD_344_U170 = ~(P3_ADD_344_U41 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_LT_563_U6 = ~(P3_LT_563_U27 & P3_LT_563_U28); 
assign P3_ADD_339_U82 = ~(P3_ADD_339_U164 & P3_ADD_339_U163); 
assign P3_ADD_339_U111 = ~P3_ADD_339_U40; 
assign P3_ADD_339_U161 = ~(P3_ADD_339_U40 & P3_PHYADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_541_U82 = ~(P3_ADD_541_U164 & P3_ADD_541_U163); 
assign P3_ADD_541_U111 = ~P3_ADD_541_U40; 
assign P3_ADD_541_U161 = ~(P3_ADD_541_U40 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_SUB_357_1258_U141 = ~(P3_SUB_357_1258_U272 & P3_SUB_357_1258_U201 & P3_SUB_357_1258_U273); 
assign P3_SUB_357_1258_U246 = ~(P3_SUB_357_1258_U202 & P3_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P3_SUB_357_1258_U442 = ~(P3_SUB_357_1258_U201 & P3_SUB_357_1258_U39); 
assign P3_SUB_357_1258_U449 = ~(P3_SUB_357_1258_U200 & P3_SUB_357_1258_U447); 
assign P3_ADD_515_U82 = ~(P3_ADD_515_U164 & P3_ADD_515_U163); 
assign P3_ADD_515_U111 = ~P3_ADD_515_U40; 
assign P3_ADD_515_U161 = ~(P3_ADD_515_U40 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_394_U82 = ~(P3_ADD_394_U168 & P3_ADD_394_U167); 
assign P3_ADD_394_U114 = ~P3_ADD_394_U40; 
assign P3_ADD_394_U163 = ~(P3_ADD_394_U40 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_441_U82 = ~(P3_ADD_441_U164 & P3_ADD_441_U163); 
assign P3_ADD_441_U111 = ~P3_ADD_441_U40; 
assign P3_ADD_441_U161 = ~(P3_ADD_441_U40 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_349_U87 = ~(P3_ADD_349_U173 & P3_ADD_349_U172); 
assign P3_ADD_349_U115 = ~P3_ADD_349_U41; 
assign P3_ADD_349_U170 = ~(P3_ADD_349_U41 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_405_U82 = ~(P3_ADD_405_U168 & P3_ADD_405_U167); 
assign P3_ADD_405_U114 = ~P3_ADD_405_U40; 
assign P3_ADD_405_U163 = ~(P3_ADD_405_U40 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_553_U87 = ~(P3_ADD_553_U173 & P3_ADD_553_U172); 
assign P3_ADD_553_U115 = ~P3_ADD_553_U41; 
assign P3_ADD_553_U170 = ~(P3_ADD_553_U41 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_558_U87 = ~(P3_ADD_558_U173 & P3_ADD_558_U172); 
assign P3_ADD_558_U115 = ~P3_ADD_558_U41; 
assign P3_ADD_558_U170 = ~(P3_ADD_558_U41 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_385_U87 = ~(P3_ADD_385_U173 & P3_ADD_385_U172); 
assign P3_ADD_385_U115 = ~P3_ADD_385_U41; 
assign P3_ADD_385_U170 = ~(P3_ADD_385_U41 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_547_U87 = ~(P3_ADD_547_U173 & P3_ADD_547_U172); 
assign P3_ADD_547_U115 = ~P3_ADD_547_U41; 
assign P3_ADD_547_U170 = ~(P3_ADD_547_U41 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_371_1212_U7 = P3_ADD_371_1212_U192 & P3_ADD_371_1212_U78; 
assign P3_ADD_371_1212_U164 = ~P3_ADD_371_1212_U78; 
assign P3_ADD_371_1212_U165 = ~P3_ADD_371_1212_U53; 
assign P3_ADD_371_1212_U258 = ~(P3_ADD_371_1212_U53 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_371_1212_U260 = ~(P3_ADD_371_1212_U78 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_494_U82 = ~(P3_ADD_494_U164 & P3_ADD_494_U163); 
assign P3_ADD_494_U111 = ~P3_ADD_494_U40; 
assign P3_ADD_494_U161 = ~(P3_ADD_494_U40 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_536_U82 = ~(P3_ADD_536_U164 & P3_ADD_536_U163); 
assign P3_ADD_536_U111 = ~P3_ADD_536_U40; 
assign P3_ADD_536_U161 = ~(P3_ADD_536_U40 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P2_R2099_U25 = ~(P2_R2099_U124 & P2_U2738); 
assign P2_R2099_U150 = ~(P2_R2099_U124 & P2_R2099_U23); 
assign P2_ADD_391_1196_U47 = ~P2_R2096_U96; 
assign P2_ADD_391_1196_U92 = ~(P2_ADD_391_1196_U350 & P2_ADD_391_1196_U349); 
assign P2_ADD_391_1196_U116 = ~(P2_ADD_391_1196_U172 & P2_ADD_391_1196_U171); 
assign P2_ADD_391_1196_U117 = P2_ADD_391_1196_U333 & P2_ADD_391_1196_U332; 
assign P2_ADD_391_1196_U325 = ~(P2_R2096_U74 & P2_ADD_391_1196_U28); 
assign P2_ADD_391_1196_U327 = ~(P2_R2096_U74 & P2_ADD_391_1196_U28); 
assign P2_ADD_391_1196_U336 = ~(P2_ADD_391_1196_U335 & P2_ADD_391_1196_U334); 
assign P2_R2182_U10 = P2_U2674 & P2_R2182_U9; 
assign P2_R2182_U74 = ~(P2_R2182_U202 & P2_R2182_U201); 
assign P2_R2182_U138 = ~P2_R2182_U9; 
assign P2_R2182_U197 = ~(P2_R2182_U35 & P2_R2182_U9); 
assign P2_R2182_U200 = ~(P2_R2182_U137 & P2_U2675); 
assign P2_R2027_U87 = ~(P2_R2027_U173 & P2_R2027_U172); 
assign P2_R2027_U115 = ~P2_R2027_U41; 
assign P2_R2027_U170 = ~(P2_R2027_U41 & P2_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P2_R2337_U80 = ~(P2_R2337_U162 & P2_R2337_U161); 
assign P2_R2337_U112 = ~P2_R2337_U41; 
assign P2_R2337_U159 = ~(P2_R2337_U41 & P2_PHYADDRPOINTER_REG_21__SCAN_IN); 
assign P2_R2096_U17 = P2_U2635 & P2_R2096_U21; 
assign P2_R2096_U95 = ~(P2_R2096_U259 & P2_R2096_U258); 
assign P2_R2096_U149 = ~P2_R2096_U21; 
assign P2_R2096_U254 = ~(P2_R2096_U31 & P2_R2096_U21); 
assign P2_R2096_U257 = ~(P2_R2096_U148 & P2_U2636); 
assign P2_R2256_U6 = ~P2_U3629; 
assign P2_R2256_U7 = ~P2_U3628; 
assign P2_R2256_U8 = ~P2_U3627; 
assign P2_R2256_U9 = ~P2_U3626; 
assign P2_R2256_U11 = ~P2_U3625; 
assign P2_R2256_U13 = ~P2_U3624; 
assign P2_R2256_U15 = ~P2_U3622; 
assign P2_R2256_U16 = ~P2_U3623; 
assign P2_R2256_U23 = P2_U3622 & P2_U3623; 
assign P2_R2256_U29 = ~(P2_U7873 & P2_U3629); 
assign P2_R2256_U30 = ~(P2_U7873 & P2_U3629 & P2_U3628); 
assign P2_R2256_U33 = ~(P2_U7873 & P2_U3629); 
assign P2_R2256_U37 = P2_U3627 | P2_U7873; 
assign P2_R2256_U39 = ~(P2_U7873 & P2_U3627); 
assign P2_R2256_U58 = ~(P2_U3627 & P2_U2616); 
assign P2_R2256_U60 = ~(P2_U3627 & P2_U2616); 
assign P2_R2256_U70 = ~(P2_U3629 & P2_U2616); 
assign P2_R1957_U31 = ~(P2_R1957_U96 & P2_R1957_U75 & P2_R1957_U44); 
assign P2_ADD_394_U82 = ~(P2_ADD_394_U166 & P2_ADD_394_U165); 
assign P2_ADD_394_U114 = ~P2_ADD_394_U40; 
assign P2_ADD_394_U137 = ~(P2_ADD_394_U40 & P2_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P2_R2267_U87 = P2_R2267_U166 & P2_R2267_U165; 
assign P2_R2267_U102 = ~P2_R2267_U31; 
assign P2_R2267_U133 = ~(P2_U2786 & P2_R2267_U132); 
assign P2_R2267_U163 = ~(P2_U2785 & P2_R2267_U31); 
assign P1_R2144_U10 = P1_R2144_U213 & P1_R2144_U212 & P1_R2144_U82; 
assign P1_R2144_U24 = ~(P1_R2144_U79 & P1_R2144_U63); 
assign P1_R2144_U25 = ~(P1_R2144_U6 & P1_R2144_U79); 
assign P1_R2144_U45 = ~(P1_R2144_U217 & P1_R2144_U216); 
assign P1_R2144_U47 = ~(P1_R2144_U219 & P1_R2144_U218); 
assign P1_R2144_U78 = ~(P1_R2144_U29 & P1_R2144_U79); 
assign P1_R2144_U96 = ~(P1_R2144_U79 & P1_R2144_U66); 
assign P1_R2144_U97 = ~(P1_R2144_U67 & P1_R2144_U79); 
assign P1_R2144_U121 = ~P1_R2144_U79; 
assign P1_R2144_U128 = ~(P1_R2144_U61 & P1_R2144_U125); 
assign P1_R2144_U211 = ~(P1_R2144_U29 & P1_R2144_U79); 
assign P1_R2278_U230 = ~P1_R2278_U213; 
assign P1_R2278_U233 = ~(P1_R2278_U33 & P1_R2278_U32); 
assign P1_R2278_U429 = ~(P1_R2278_U557 & P1_R2278_U33); 
assign P1_R2358_U106 = P1_R2358_U206 & P1_R2358_U205; 
assign P1_R2358_U120 = P1_R2358_U208 & P1_R2358_U205; 
assign P1_R2358_U164 = ~P1_U2665; 
assign P1_R2358_U193 = ~(P1_R2358_U209 & P1_R2358_U246); 
assign P1_R2358_U331 = ~P1_R2358_U200; 
assign P1_R2358_U346 = ~(P1_R2358_U206 & P1_R2358_U205); 
assign P1_R2358_U490 = ~(P1_U2665 & P1_R2358_U23); 
assign P1_R2358_U497 = ~(P1_U2665 & P1_R2358_U23); 
assign P1_R2358_U501 = ~(P1_R2358_U500 & P1_R2358_U499); 
assign P1_R2358_U610 = ~(P1_U2352 & P1_R2358_U200); 
assign P1_LT_589_U8 = ~(P1_LT_589_U7 | P1_R584_U9 | P1_R584_U8); 
assign P1_R2099_U77 = ~(P1_R2099_U328 & P1_R2099_U327); 
assign P1_R2099_U78 = ~(P1_R2099_U330 & P1_R2099_U329); 
assign P1_R2099_U170 = ~P1_R2099_U15; 
assign P1_R2099_U326 = ~(P1_R2099_U54 & P1_R2099_U15); 
assign P1_R2337_U82 = ~(P1_R2337_U164 & P1_R2337_U163); 
assign P1_R2337_U111 = ~P1_R2337_U40; 
assign P1_R2337_U161 = ~(P1_R2337_U40 & P1_PHYADDRPOINTER_REG_20__SCAN_IN); 
assign P1_LT_563_1260_U6 = P1_LT_563_1260_U9 & P1_LT_563_1260_U8; 
assign P1_R2096_U82 = ~(P1_R2096_U164 & P1_R2096_U163); 
assign P1_R2096_U111 = ~P1_R2096_U40; 
assign P1_R2096_U161 = ~(P1_R2096_U40 & P1_REIP_REG_20__SCAN_IN); 
assign P1_LT_563_U26 = ~(P1_LT_563_U14 & P1_LT_563_U23); 
assign P1_ADD_405_U82 = ~(P1_ADD_405_U166 & P1_ADD_405_U165); 
assign P1_ADD_405_U114 = ~P1_ADD_405_U40; 
assign P1_ADD_405_U137 = ~(P1_ADD_405_U40 & P1_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P1_ADD_515_U82 = ~(P1_ADD_515_U164 & P1_ADD_515_U163); 
assign P1_ADD_515_U111 = ~P1_ADD_515_U40; 
assign P1_ADD_515_U135 = ~(P1_ADD_515_U40 & P1_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_U2819 = ~(P3_U6494 & P3_U6493 & P3_U6495 & P3_U6496 & P3_U3965); 
assign P3_U3120 = ~(P3_U7949 & P3_U7948 & P3_U3262 & P3_U4313 & P3_LT_563_U6); 
assign P3_U3788 = P3_U3787 & P3_U3786 & P3_U5939; 
assign P3_U3789 = P3_U3790 & P3_U5944; 
assign P3_U3966 = P3_U6508 & P3_U6505 & P3_U6506 & P3_U6507; 
assign P3_U5870 = ~(P3_U4318 & P3_U5868); 
assign P3_U5894 = ~(P3_U4318 & P3_U5892); 
assign P3_U5916 = ~(P3_U5898 & P3_U3778 & P3_U5896 & P3_U3775 & P3_U3781); 
assign P3_U5963 = ~(P3_ADD_371_1212_U7 & P3_U2360); 
assign P3_U6066 = ~(P3_ADD_558_U87 & P3_U3220); 
assign P3_U6067 = ~(P3_ADD_553_U87 & P3_U4298); 
assign P3_U6068 = ~(P3_ADD_547_U87 & P3_U4299); 
assign P3_U6071 = ~(P3_ADD_531_U87 & P3_U2354); 
assign P3_U6079 = ~(P3_ADD_385_U87 & P3_U2358); 
assign P3_U6080 = ~(P3_ADD_380_U87 & P3_U2359); 
assign P3_U6081 = ~(P3_ADD_349_U87 & P3_U4306); 
assign P3_U6082 = ~(P3_ADD_344_U87 & P3_U2362); 
assign P3_U6093 = ~(P3_ADD_541_U82 & P3_U4300); 
assign P3_U6094 = ~(P3_ADD_536_U82 & P3_U4301); 
assign P3_U6097 = ~(P3_ADD_515_U82 & P3_U4302); 
assign P3_U6098 = ~(P3_ADD_494_U82 & P3_U2356); 
assign P3_U6099 = ~(P3_ADD_476_U82 & P3_U4303); 
assign P3_U6100 = ~(P3_ADD_441_U82 & P3_U4304); 
assign P3_U6101 = ~(P3_ADD_405_U82 & P3_U4305); 
assign P3_U6102 = ~(P3_ADD_394_U82 & P3_U2357); 
assign P3_U6515 = ~(P3_U2387 & P3_ADD_371_1212_U7); 
assign P3_U6557 = ~(P3_ADD_318_U82 & P3_U2398); 
assign P3_U6562 = ~(P3_ADD_339_U82 & P3_U2388); 
assign P3_U6566 = ~(P3_ADD_315_U78 & P3_U2397); 
assign P3_U7262 = ~(P3_ADD_467_U82 & P3_U2601); 
assign P3_U7264 = ~(P3_ADD_430_U82 & P3_U2405); 
assign P2_U2362 = P2_U2398 & P2_U4443; 
assign P2_U2364 = P2_U3546 & P2_STATE2_REG_2__SCAN_IN; 
assign P2_U2365 = P2_U4443 & P2_STATE2_REG_3__SCAN_IN; 
assign P2_U2366 = P2_U3546 & P2_STATE2_REG_1__SCAN_IN; 
assign P2_U2378 = P2_U3546 & P2_STATE2_REG_3__SCAN_IN; 
assign P2_U2396 = P2_U3541 & P2_U3284; 
assign P2_U2399 = U314 & P2_U4443; 
assign P2_U2400 = U303 & P2_U4443; 
assign P2_U2401 = U292 & P2_U4443; 
assign P2_U2402 = U289 & P2_U4443; 
assign P2_U2403 = U288 & P2_U4443; 
assign P2_U2404 = U287 & P2_U4443; 
assign P2_U2405 = U286 & P2_U4443; 
assign P2_U2406 = U285 & P2_U4443; 
assign P2_U2430 = P2_U3541 & P2_STATE2_REG_0__SCAN_IN; 
assign P2_U2435 = P2_U2356 & P2_U3541; 
assign P2_U2811 = P2_U3242 & P2_R2267_U87; 
assign P2_U3291 = ~(P2_U3713 & P2_U2459); 
assign P2_U3426 = ~(P2_U3378 & P2_U4639 & P2_U3425); 
assign P2_U3722 = P2_U4661 & P2_U4662 & P2_U4443; 
assign P2_U3731 = P2_U4719 & P2_U4720 & P2_U4443; 
assign P2_U3740 = P2_U4778 & P2_U4779 & P2_U4443; 
assign P2_U3749 = P2_U4835 & P2_U4836 & P2_U4443; 
assign P2_U3758 = P2_U4893 & P2_U4894 & P2_U4443; 
assign P2_U3767 = P2_U4950 & P2_U4951 & P2_U4443; 
assign P2_U3776 = P2_U5008 & P2_U5009 & P2_U4443; 
assign P2_U3785 = P2_U5065 & P2_U5066 & P2_U4443; 
assign P2_U3794 = P2_U5121 & P2_U5122 & P2_U4443; 
assign P2_U3803 = P2_U5178 & P2_U5179 & P2_U4443; 
assign P2_U3812 = P2_U5236 & P2_U5237 & P2_U4443; 
assign P2_U3821 = P2_U5293 & P2_U5294 & P2_U4443; 
assign P2_U3830 = P2_U5351 & P2_U5352 & P2_U4443; 
assign P2_U3839 = P2_U5408 & P2_U5409 & P2_U4443; 
assign P2_U3848 = P2_U5466 & P2_U5467 & P2_U4443; 
assign P2_U3857 = P2_U5523 & P2_U5524 & P2_U4443; 
assign P2_U4440 = ~P2_U3543; 
assign P2_U4441 = ~P2_U3542; 
assign P2_U4446 = ~(P2_U4461 & P2_U3546); 
assign P2_U4451 = ~P2_U3425; 
assign P2_U5581 = ~P2_U4406; 
assign P2_U5582 = ~(P2_U2374 & P2_U4406); 
assign P2_U5660 = ~(P2_U3893 & P2_U5657); 
assign P2_U6232 = ~P2_U3541; 
assign P2_U6330 = ~(P2_U3542 & P2_EAX_REG_0__SCAN_IN); 
assign P2_U6334 = ~(P2_U3542 & P2_EAX_REG_1__SCAN_IN); 
assign P2_U6338 = ~(P2_U3542 & P2_EAX_REG_2__SCAN_IN); 
assign P2_U6342 = ~(P2_U3542 & P2_EAX_REG_3__SCAN_IN); 
assign P2_U6346 = ~(P2_U3542 & P2_EAX_REG_4__SCAN_IN); 
assign P2_U6350 = ~(P2_U3542 & P2_EAX_REG_5__SCAN_IN); 
assign P2_U6354 = ~(P2_U3542 & P2_EAX_REG_6__SCAN_IN); 
assign P2_U6358 = ~(P2_U3542 & P2_EAX_REG_7__SCAN_IN); 
assign P2_U6362 = ~(P2_U3542 & P2_EAX_REG_8__SCAN_IN); 
assign P2_U6366 = ~(P2_U3542 & P2_EAX_REG_9__SCAN_IN); 
assign P2_U6370 = ~(P2_U3542 & P2_EAX_REG_10__SCAN_IN); 
assign P2_U6374 = ~(P2_U3542 & P2_EAX_REG_11__SCAN_IN); 
assign P2_U6378 = ~(P2_U3542 & P2_EAX_REG_12__SCAN_IN); 
assign P2_U6382 = ~(P2_U3542 & P2_EAX_REG_13__SCAN_IN); 
assign P2_U6386 = ~(P2_U3542 & P2_EAX_REG_14__SCAN_IN); 
assign P2_U6390 = ~(P2_U3542 & P2_EAX_REG_15__SCAN_IN); 
assign P2_U6395 = ~(P2_U3542 & P2_EAX_REG_16__SCAN_IN); 
assign P2_U6400 = ~(P2_U3542 & P2_EAX_REG_17__SCAN_IN); 
assign P2_U6405 = ~(P2_U3542 & P2_EAX_REG_18__SCAN_IN); 
assign P2_U6410 = ~(P2_U3542 & P2_EAX_REG_19__SCAN_IN); 
assign P2_U6415 = ~(P2_U3542 & P2_EAX_REG_20__SCAN_IN); 
assign P2_U6420 = ~(P2_U3542 & P2_EAX_REG_21__SCAN_IN); 
assign P2_U6425 = ~(P2_U3542 & P2_EAX_REG_22__SCAN_IN); 
assign P2_U6430 = ~(P2_U3542 & P2_EAX_REG_23__SCAN_IN); 
assign P2_U6435 = ~(P2_U3542 & P2_EAX_REG_24__SCAN_IN); 
assign P2_U6440 = ~(P2_U3542 & P2_EAX_REG_25__SCAN_IN); 
assign P2_U6445 = ~(P2_U3542 & P2_EAX_REG_26__SCAN_IN); 
assign P2_U6450 = ~(P2_U3542 & P2_EAX_REG_27__SCAN_IN); 
assign P2_U6455 = ~(P2_U3542 & P2_EAX_REG_28__SCAN_IN); 
assign P2_U6460 = ~(P2_U3542 & P2_EAX_REG_29__SCAN_IN); 
assign P2_U6465 = ~(P2_U3542 & P2_EAX_REG_30__SCAN_IN); 
assign P2_U6468 = ~(P2_U3542 & P2_EAX_REG_31__SCAN_IN); 
assign P2_U6473 = ~(P2_U3543 & P2_EBX_REG_0__SCAN_IN); 
assign P2_U6476 = ~(P2_U3543 & P2_EBX_REG_1__SCAN_IN); 
assign P2_U6479 = ~(P2_U3543 & P2_EBX_REG_2__SCAN_IN); 
assign P2_U6482 = ~(P2_U3543 & P2_EBX_REG_3__SCAN_IN); 
assign P2_U6485 = ~(P2_U3543 & P2_EBX_REG_4__SCAN_IN); 
assign P2_U6488 = ~(P2_U3543 & P2_EBX_REG_5__SCAN_IN); 
assign P2_U6491 = ~(P2_U3543 & P2_EBX_REG_6__SCAN_IN); 
assign P2_U6494 = ~(P2_U3543 & P2_EBX_REG_7__SCAN_IN); 
assign P2_U6497 = ~(P2_U3543 & P2_EBX_REG_8__SCAN_IN); 
assign P2_U6500 = ~(P2_U3543 & P2_EBX_REG_9__SCAN_IN); 
assign P2_U6503 = ~(P2_U3543 & P2_EBX_REG_10__SCAN_IN); 
assign P2_U6506 = ~(P2_U3543 & P2_EBX_REG_11__SCAN_IN); 
assign P2_U6509 = ~(P2_U3543 & P2_EBX_REG_12__SCAN_IN); 
assign P2_U6512 = ~(P2_U3543 & P2_EBX_REG_13__SCAN_IN); 
assign P2_U6515 = ~(P2_U3543 & P2_EBX_REG_14__SCAN_IN); 
assign P2_U6518 = ~(P2_U3543 & P2_EBX_REG_15__SCAN_IN); 
assign P2_U6521 = ~(P2_U3543 & P2_EBX_REG_16__SCAN_IN); 
assign P2_U6524 = ~(P2_U3543 & P2_EBX_REG_17__SCAN_IN); 
assign P2_U6527 = ~(P2_U3543 & P2_EBX_REG_18__SCAN_IN); 
assign P2_U6530 = ~(P2_U3543 & P2_EBX_REG_19__SCAN_IN); 
assign P2_U6533 = ~(P2_U3543 & P2_EBX_REG_20__SCAN_IN); 
assign P2_U6536 = ~(P2_U3543 & P2_EBX_REG_21__SCAN_IN); 
assign P2_U6539 = ~(P2_U3543 & P2_EBX_REG_22__SCAN_IN); 
assign P2_U6542 = ~(P2_U3543 & P2_EBX_REG_23__SCAN_IN); 
assign P2_U6545 = ~(P2_U3543 & P2_EBX_REG_24__SCAN_IN); 
assign P2_U6548 = ~(P2_U3543 & P2_EBX_REG_25__SCAN_IN); 
assign P2_U6551 = ~(P2_U3543 & P2_EBX_REG_26__SCAN_IN); 
assign P2_U6554 = ~(P2_U3543 & P2_EBX_REG_27__SCAN_IN); 
assign P2_U6557 = ~(P2_U3543 & P2_EBX_REG_28__SCAN_IN); 
assign P2_U6560 = ~(P2_U3543 & P2_EBX_REG_29__SCAN_IN); 
assign P2_U6563 = ~(P2_U3543 & P2_EBX_REG_30__SCAN_IN); 
assign P2_U6565 = ~(P2_U3543 & P2_EBX_REG_31__SCAN_IN); 
assign P2_U6570 = ~P2_U3546; 
assign P2_U6843 = ~P2_U4402; 
assign P2_U6853 = ~(P2_U2374 & P2_U2459); 
assign P2_U6857 = ~P2_U4403; 
assign P2_U6861 = ~(P2_U6859 & P2_MEMORYFETCH_REG_SCAN_IN); 
assign P2_U8109 = ~(P2_U8108 & P2_U8107); 
assign P2_U8138 = ~(P2_U6852 & P2_U4402); 
assign P2_U8144 = ~(P2_U6858 & P2_U4403); 
assign P2_U8287 = ~(P2_U3616 & P2_U4406); 
assign P2_U8290 = ~(P2_U5611 & P2_U4406); 
assign P2_U8292 = ~(P2_U5619 & P2_U4406); 
assign P2_U8294 = ~(P2_U5629 & P2_U4406); 
assign P2_U8296 = ~(P2_U5637 & P2_U4406); 
assign P2_U8395 = ~(P2_R2337_U80 & P2_U3284); 
assign P1_U2474 = P1_R2144_U49 & P1_U3312; 
assign P1_U2477 = P1_U4528 & P1_U2476; 
assign P1_U2481 = P1_U4524 & P1_U2476; 
assign P1_U2483 = P1_U4525 & P1_U2476; 
assign P1_U2485 = P1_U4526 & P1_R2144_U43; 
assign P1_U2487 = P1_U2486 & P1_U2476; 
assign P1_U2509 = P1_U2508 & P1_U4528; 
assign P1_U2512 = P1_U2508 & P1_U4524; 
assign P1_U2514 = P1_U2508 & P1_U4525; 
assign P1_U2516 = P1_U2508 & P1_U2486; 
assign P1_U2643 = P1_R2144_U10 & P1_U6746; 
assign P1_U2645 = P1_R2144_U45 & P1_U6746; 
assign P1_U2646 = P1_R2144_U47 & P1_U6746; 
assign P1_U2664 = ~(P1_U6829 & P1_U4023); 
assign P1_U2797 = ~(P1_U6882 & P1_U6881); 
assign P1_U3031 = ~(P1_U3764 & P1_U3763 & P1_U3766); 
assign P1_U3333 = ~(P1_U4526 & P1_U3309); 
assign P1_U3454 = ~(P1_U7692 & P1_U7691); 
assign P1_U3751 = P1_U5543 & P1_U5544; 
assign P1_U3894 = P1_U6400 & P1_U4227; 
assign P1_U3896 = P1_U6408 & P1_U4227; 
assign P1_U3898 = P1_U6416 & P1_U4227; 
assign P1_U3900 = P1_U6423 & P1_U4227; 
assign P1_U3902 = P1_U6430 & P1_U4227; 
assign P1_U3904 = P1_U6437 & P1_U4227; 
assign P1_U3906 = P1_U6444 & P1_U4227; 
assign P1_U3908 = P1_U6451 & P1_U4227; 
assign P1_U3910 = P1_U6458 & P1_U4227; 
assign P1_U3912 = P1_U6465 & P1_U4227; 
assign P1_U3914 = P1_U6472 & P1_U4227; 
assign P1_U3916 = P1_U6479 & P1_U4227; 
assign P1_U3918 = P1_U6486 & P1_U4227; 
assign P1_U4225 = ~P1_LT_563_1260_U6; 
assign P1_U4527 = ~P1_U3314; 
assign P1_U4529 = ~P1_U3342; 
assign P1_U4548 = ~(P1_U4528 & P1_U2476); 
assign P1_U4600 = ~P1_U3326; 
assign P1_U4606 = ~(P1_U4524 & P1_U2476); 
assign P1_U4665 = ~(P1_U4525 & P1_U2476); 
assign P1_U4722 = ~(P1_U2486 & P1_U2476); 
assign P1_U5238 = ~(P1_U2508 & P1_U4528); 
assign P1_U5295 = ~(P1_U2508 & P1_U4524); 
assign P1_U5353 = ~(P1_U2508 & P1_U4525); 
assign P1_U5410 = ~(P1_U2508 & P1_U2486); 
assign P1_U5689 = ~(P1_R2099_U78 & P1_U2380); 
assign P1_U5696 = ~(P1_R2099_U77 & P1_U2380); 
assign P1_U5706 = ~(P1_ADD_405_U82 & P1_U2375); 
assign P1_U5707 = ~(P1_ADD_515_U82 & P1_U2374); 
assign P1_U5894 = ~(P1_R2337_U82 & P1_U2376); 
assign P1_U6317 = ~(P1_U2371 & P1_R2099_U78); 
assign P1_U6320 = ~(P1_U2371 & P1_R2099_U77); 
assign P1_U6369 = ~(P1_U7485 & P1_REIP_REG_0__SCAN_IN); 
assign P1_U6370 = ~(P1_U7484 & P1_EBX_REG_0__SCAN_IN); 
assign P1_U6377 = ~(P1_R2096_U4 & P1_U7485); 
assign P1_U6378 = ~(P1_U7484 & P1_EBX_REG_1__SCAN_IN); 
assign P1_U6385 = ~(P1_R2096_U71 & P1_U7485); 
assign P1_U6386 = ~(P1_U7484 & P1_EBX_REG_2__SCAN_IN); 
assign P1_U6393 = ~(P1_R2096_U68 & P1_U7485); 
assign P1_U6394 = ~(P1_U7484 & P1_EBX_REG_3__SCAN_IN); 
assign P1_U6401 = ~(P1_R2096_U67 & P1_U7485); 
assign P1_U6402 = ~(P1_U7484 & P1_EBX_REG_4__SCAN_IN); 
assign P1_U6409 = ~(P1_R2096_U66 & P1_U7485); 
assign P1_U6410 = ~(P1_U7484 & P1_EBX_REG_5__SCAN_IN); 
assign P1_U6417 = ~(P1_R2096_U65 & P1_U7485); 
assign P1_U6418 = ~(P1_U7484 & P1_EBX_REG_6__SCAN_IN); 
assign P1_U6424 = ~(P1_R2096_U64 & P1_U7485); 
assign P1_U6425 = ~(P1_U7484 & P1_EBX_REG_7__SCAN_IN); 
assign P1_U6431 = ~(P1_R2096_U63 & P1_U7485); 
assign P1_U6432 = ~(P1_U7484 & P1_EBX_REG_8__SCAN_IN); 
assign P1_U6438 = ~(P1_R2096_U62 & P1_U7485); 
assign P1_U6439 = ~(P1_U7484 & P1_EBX_REG_9__SCAN_IN); 
assign P1_U6445 = ~(P1_R2096_U91 & P1_U7485); 
assign P1_U6446 = ~(P1_U7484 & P1_EBX_REG_10__SCAN_IN); 
assign P1_U6452 = ~(P1_R2096_U90 & P1_U7485); 
assign P1_U6453 = ~(P1_U7484 & P1_EBX_REG_11__SCAN_IN); 
assign P1_U6459 = ~(P1_R2096_U89 & P1_U7485); 
assign P1_U6460 = ~(P1_U7484 & P1_EBX_REG_12__SCAN_IN); 
assign P1_U6466 = ~(P1_R2096_U88 & P1_U7485); 
assign P1_U6467 = ~(P1_U7484 & P1_EBX_REG_13__SCAN_IN); 
assign P1_U6473 = ~(P1_R2096_U87 & P1_U7485); 
assign P1_U6474 = ~(P1_U7484 & P1_EBX_REG_14__SCAN_IN); 
assign P1_U6480 = ~(P1_R2096_U86 & P1_U7485); 
assign P1_U6481 = ~(P1_U7484 & P1_EBX_REG_15__SCAN_IN); 
assign P1_U6487 = ~(P1_R2096_U85 & P1_U7485); 
assign P1_U6488 = ~(P1_U7484 & P1_EBX_REG_16__SCAN_IN); 
assign P1_U6493 = ~(P1_U2604 & P1_R2099_U78); 
assign P1_U6494 = ~(P1_R2096_U84 & P1_U7485); 
assign P1_U6495 = ~(P1_U7484 & P1_EBX_REG_17__SCAN_IN); 
assign P1_U6500 = ~(P1_U2604 & P1_R2099_U77); 
assign P1_U6501 = ~(P1_R2096_U83 & P1_U7485); 
assign P1_U6502 = ~(P1_U7484 & P1_EBX_REG_18__SCAN_IN); 
assign P1_U6508 = ~(P1_R2096_U82 & P1_U7485); 
assign P1_U6509 = ~(P1_U7484 & P1_EBX_REG_19__SCAN_IN); 
assign P1_U6516 = ~(P1_U7484 & P1_EBX_REG_20__SCAN_IN); 
assign P1_U6523 = ~(P1_U7484 & P1_EBX_REG_21__SCAN_IN); 
assign P1_U6530 = ~(P1_U7484 & P1_EBX_REG_22__SCAN_IN); 
assign P1_U6537 = ~(P1_U7484 & P1_EBX_REG_23__SCAN_IN); 
assign P1_U6544 = ~(P1_U7484 & P1_EBX_REG_24__SCAN_IN); 
assign P1_U6551 = ~(P1_U7484 & P1_EBX_REG_25__SCAN_IN); 
assign P1_U6558 = ~(P1_U7484 & P1_EBX_REG_26__SCAN_IN); 
assign P1_U6565 = ~(P1_U7484 & P1_EBX_REG_27__SCAN_IN); 
assign P1_U6572 = ~(P1_U7484 & P1_EBX_REG_28__SCAN_IN); 
assign P1_U6579 = ~(P1_U7484 & P1_EBX_REG_29__SCAN_IN); 
assign P1_U6586 = ~(P1_U7484 & P1_EBX_REG_30__SCAN_IN); 
assign P1_U6593 = ~(P1_U7484 & P1_EBX_REG_31__SCAN_IN); 
assign P1_U6828 = ~(P1_R2337_U82 & P1_U2352); 
assign P1_U6873 = ~(P1_U4159 & P1_R2144_U10); 
assign P1_U6877 = ~(P1_U4159 & P1_R2144_U45); 
assign P1_U6879 = ~(P1_U4159 & P1_R2144_U47); 
assign P3_ADD_476_U42 = ~(P3_ADD_476_U111 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_476_U162 = ~(P3_ADD_476_U111 & P3_ADD_476_U41); 
assign P3_ADD_531_U43 = ~(P3_ADD_531_U115 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_531_U171 = ~(P3_ADD_531_U115 & P3_ADD_531_U42); 
assign P3_SUB_320_U10 = P3_SUB_320_U118 & P3_SUB_320_U32; 
assign P3_SUB_320_U73 = ~P3_ADD_318_U82; 
assign P3_SUB_320_U97 = ~P3_SUB_320_U32; 
assign P3_SUB_320_U150 = ~(P3_ADD_318_U82 & P3_SUB_320_U32); 
assign P3_ADD_318_U42 = ~(P3_ADD_318_U111 & P3_PHYADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_318_U162 = ~(P3_ADD_318_U111 & P3_ADD_318_U41); 
assign P3_ADD_315_U42 = ~(P3_ADD_315_U108 & P3_PHYADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_315_U154 = ~(P3_ADD_315_U108 & P3_ADD_315_U41); 
assign P3_ADD_360_1242_U82 = ~(P3_ADD_360_1242_U252 & P3_ADD_360_1242_U251); 
assign P3_ADD_360_1242_U83 = ~(P3_ADD_360_1242_U254 & P3_ADD_360_1242_U253); 
assign P3_ADD_360_1242_U157 = ~P3_ADD_360_1242_U53; 
assign P3_ADD_360_1242_U179 = ~(P3_ADD_360_1242_U51 & P3_ADD_360_1242_U178); 
assign P3_ADD_360_1242_U181 = ~(P3_ADD_360_1242_U48 & P3_ADD_360_1242_U180); 
assign P3_ADD_360_1242_U249 = ~(P3_ADD_360_1242_U53 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_467_U42 = ~(P3_ADD_467_U111 & P3_REIP_REG_20__SCAN_IN); 
assign P3_ADD_467_U162 = ~(P3_ADD_467_U111 & P3_ADD_467_U41); 
assign P3_ADD_430_U42 = ~(P3_ADD_430_U111 & P3_REIP_REG_20__SCAN_IN); 
assign P3_ADD_430_U162 = ~(P3_ADD_430_U111 & P3_ADD_430_U41); 
assign P3_ADD_380_U43 = ~(P3_ADD_380_U115 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_380_U171 = ~(P3_ADD_380_U115 & P3_ADD_380_U42); 
assign P3_ADD_344_U43 = ~(P3_ADD_344_U115 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_344_U171 = ~(P3_ADD_344_U115 & P3_ADD_344_U42); 
assign P3_ADD_339_U42 = ~(P3_ADD_339_U111 & P3_PHYADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_339_U162 = ~(P3_ADD_339_U111 & P3_ADD_339_U41); 
assign P3_ADD_541_U42 = ~(P3_ADD_541_U111 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_541_U162 = ~(P3_ADD_541_U111 & P3_ADD_541_U41); 
assign P3_SUB_357_1258_U88 = ~(P3_SUB_357_1258_U449 & P3_SUB_357_1258_U448); 
assign P3_SUB_357_1258_U203 = ~P3_SUB_357_1258_U141; 
assign P3_SUB_357_1258_U249 = ~(P3_SUB_357_1258_U442 & P3_SUB_357_1258_U441 & P3_SUB_357_1258_U67); 
assign P3_SUB_357_1258_U276 = ~(P3_SUB_357_1258_U204 & P3_SUB_357_1258_U141); 
assign P3_SUB_357_1258_U278 = ~(P3_SUB_357_1258_U9 & P3_SUB_357_1258_U141); 
assign P3_SUB_357_1258_U280 = ~(P3_SUB_357_1258_U11 & P3_SUB_357_1258_U141); 
assign P3_SUB_357_1258_U282 = ~(P3_SUB_357_1258_U13 & P3_SUB_357_1258_U141); 
assign P3_SUB_357_1258_U284 = ~(P3_SUB_357_1258_U103 & P3_SUB_357_1258_U141); 
assign P3_SUB_357_1258_U437 = ~(P3_SUB_357_1258_U140 & P3_SUB_357_1258_U141); 
assign P3_SUB_357_1258_U440 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U246); 
assign P3_ADD_515_U42 = ~(P3_ADD_515_U111 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_515_U162 = ~(P3_ADD_515_U111 & P3_ADD_515_U41); 
assign P3_ADD_394_U42 = ~(P3_ADD_394_U114 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_394_U164 = ~(P3_ADD_394_U114 & P3_ADD_394_U41); 
assign P3_ADD_441_U42 = ~(P3_ADD_441_U111 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_441_U162 = ~(P3_ADD_441_U111 & P3_ADD_441_U41); 
assign P3_ADD_349_U43 = ~(P3_ADD_349_U115 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_349_U171 = ~(P3_ADD_349_U115 & P3_ADD_349_U42); 
assign P3_ADD_405_U42 = ~(P3_ADD_405_U114 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_405_U164 = ~(P3_ADD_405_U114 & P3_ADD_405_U41); 
assign P3_ADD_553_U43 = ~(P3_ADD_553_U115 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_553_U171 = ~(P3_ADD_553_U115 & P3_ADD_553_U42); 
assign P3_ADD_558_U43 = ~(P3_ADD_558_U115 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_558_U171 = ~(P3_ADD_558_U115 & P3_ADD_558_U42); 
assign P3_ADD_385_U43 = ~(P3_ADD_385_U115 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_385_U171 = ~(P3_ADD_385_U115 & P3_ADD_385_U42); 
assign P3_ADD_547_U43 = ~(P3_ADD_547_U115 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_ADD_547_U171 = ~(P3_ADD_547_U115 & P3_ADD_547_U42); 
assign P3_ADD_371_1212_U56 = ~(P3_ADD_371_1212_U102 & P3_ADD_371_1212_U165); 
assign P3_ADD_371_1212_U188 = ~(P3_ADD_371_1212_U165 & P3_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P3_ADD_371_1212_U190 = ~(P3_ADD_371_1212_U164 & P3_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P3_ADD_371_1212_U259 = ~(P3_ADD_371_1212_U165 & P3_ADD_371_1212_U55); 
assign P3_ADD_371_1212_U261 = ~(P3_ADD_371_1212_U164 & P3_ADD_371_1212_U52); 
assign P3_ADD_494_U42 = ~(P3_ADD_494_U111 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_494_U162 = ~(P3_ADD_494_U111 & P3_ADD_494_U41); 
assign P3_ADD_536_U42 = ~(P3_ADD_536_U111 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_536_U162 = ~(P3_ADD_536_U111 & P3_ADD_536_U41); 
assign P2_R2099_U67 = ~(P2_R2099_U150 & P2_R2099_U149); 
assign P2_R2099_U125 = ~P2_R2099_U25; 
assign P2_R2099_U222 = ~(P2_U2737 & P2_R2099_U25); 
assign P2_ADD_391_1196_U17 = ~P2_R2182_U74; 
assign P2_ADD_391_1196_U52 = ~P2_R2096_U95; 
assign P2_ADD_391_1196_U115 = P2_ADD_391_1196_U326 & P2_ADD_391_1196_U325; 
assign P2_ADD_391_1196_U173 = ~P2_ADD_391_1196_U116; 
assign P2_ADD_391_1196_U175 = ~(P2_ADD_391_1196_U174 & P2_ADD_391_1196_U116); 
assign P2_ADD_391_1196_U178 = P2_R2096_U73 | P2_R2182_U74; 
assign P2_ADD_391_1196_U180 = ~(P2_R2096_U73 & P2_R2182_U74); 
assign P2_ADD_391_1196_U204 = ~(P2_R2096_U73 & P2_R2182_U74); 
assign P2_ADD_391_1196_U324 = ~(P2_R2182_U74 & P2_ADD_391_1196_U18); 
assign P2_ADD_391_1196_U329 = ~(P2_ADD_391_1196_U328 & P2_ADD_391_1196_U327); 
assign P2_ADD_391_1196_U337 = ~(P2_ADD_391_1196_U117 & P2_ADD_391_1196_U118); 
assign P2_ADD_391_1196_U338 = ~(P2_ADD_391_1196_U169 & P2_ADD_391_1196_U336); 
assign P2_R2182_U19 = P2_U2673 & P2_R2182_U10; 
assign P2_R2182_U73 = ~(P2_R2182_U200 & P2_R2182_U199); 
assign P2_R2182_U139 = ~P2_R2182_U10; 
assign P2_R2182_U195 = ~(P2_R2182_U36 & P2_R2182_U10); 
assign P2_R2182_U198 = ~(P2_R2182_U138 & P2_U2674); 
assign P2_R2027_U43 = ~(P2_R2027_U115 & P2_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P2_R2027_U171 = ~(P2_R2027_U115 & P2_R2027_U42); 
assign P2_R2337_U43 = ~(P2_R2337_U112 & P2_PHYADDRPOINTER_REG_21__SCAN_IN); 
assign P2_R2337_U160 = ~(P2_R2337_U112 & P2_R2337_U42); 
assign P2_R2096_U18 = P2_U2634 & P2_R2096_U17; 
assign P2_R2096_U94 = ~(P2_R2096_U257 & P2_R2096_U256); 
assign P2_R2096_U150 = ~P2_R2096_U17; 
assign P2_R2096_U252 = ~(P2_R2096_U35 & P2_R2096_U17); 
assign P2_R2096_U255 = ~(P2_R2096_U149 & P2_U2635); 
assign P2_R2256_U32 = ~P2_R2256_U30; 
assign P2_R2256_U34 = ~(P2_R2256_U7 & P2_R2256_U33); 
assign P2_R2256_U45 = ~P2_R2256_U29; 
assign P2_R2256_U57 = ~(P2_U7873 & P2_R2256_U8); 
assign P2_R2256_U59 = ~(P2_U7873 & P2_R2256_U8); 
assign P2_R2256_U64 = ~(P2_U2616 & P2_R2256_U29); 
assign P2_R2256_U67 = ~(P2_U3628 & P2_R2256_U33 & P2_U7873); 
assign P2_R2256_U69 = ~(P2_U7873 & P2_R2256_U6); 
assign P2_R1957_U10 = P2_R1957_U118 & P2_R1957_U31; 
assign P2_R1957_U73 = ~P2_U3672; 
assign P2_R1957_U97 = ~P2_R1957_U31; 
assign P2_R1957_U150 = ~(P2_U3672 & P2_R1957_U31); 
assign P2_R2278_U30 = ~P2_U2812; 
assign P2_R2278_U235 = P2_U2812 | P2_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P2_R2278_U236 = ~(P2_U2812 & P2_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P2_R2278_U347 = ~(P2_U2812 & P2_R2278_U29); 
assign P2_R2278_U349 = ~(P2_U2812 & P2_R2278_U29); 
assign P2_ADD_394_U42 = ~(P2_ADD_394_U114 & P2_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P2_ADD_394_U138 = ~(P2_ADD_394_U114 & P2_ADD_394_U41); 
assign P2_R2267_U6 = P2_R2267_U133 & P2_R2267_U31; 
assign P2_R2267_U32 = ~(P2_R2267_U46 & P2_R2267_U102); 
assign P2_R2267_U130 = ~(P2_R2267_U102 & P2_R2267_U84); 
assign P2_R2267_U164 = ~(P2_R2267_U102 & P2_R2267_U84); 
assign P1_R2144_U9 = P1_R2144_U128 & P1_R2144_U127; 
assign P1_R2144_U101 = ~P1_R2144_U24; 
assign P1_R2144_U122 = ~P1_R2144_U78; 
assign P1_R2144_U139 = ~P1_R2144_U97; 
assign P1_R2144_U140 = ~P1_R2144_U96; 
assign P1_R2144_U141 = ~P1_R2144_U25; 
assign P1_R2144_U144 = ~(P1_U2355 & P1_R2144_U24); 
assign P1_R2144_U209 = ~(P1_R2144_U27 & P1_R2144_U78); 
assign P1_R2144_U210 = ~(P1_R2144_U121 & P1_R2144_U204); 
assign P1_R2144_U254 = ~(P1_R2144_U34 & P1_R2144_U25); 
assign P1_R2144_U256 = ~(P1_R2144_U35 & P1_R2144_U96); 
assign P1_R2144_U258 = ~(P1_R2144_U36 & P1_R2144_U97); 
assign P1_R2278_U35 = ~P1_U2798; 
assign P1_R2278_U234 = ~(P1_R2278_U233 & P1_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P1_R2278_U236 = P1_U2798 | P1_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P1_R2278_U238 = ~(P1_U2798 & P1_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P1_R2278_U478 = ~(P1_U2798 & P1_R2278_U34); 
assign P1_R2278_U480 = ~(P1_U2798 & P1_R2278_U34); 
assign P1_R2278_U559 = ~(P1_R2278_U230 & P1_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P1_R2358_U30 = ~P1_U2648; 
assign P1_R2358_U32 = ~P1_U2647; 
assign P1_R2358_U203 = ~(P1_U2647 & P1_R2358_U441); 
assign P1_R2358_U207 = ~(P1_U2648 & P1_R2358_U424); 
assign P1_R2358_U211 = ~(P1_R2358_U120 & P1_R2358_U210); 
assign P1_R2358_U247 = ~P1_R2358_U193; 
assign P1_R2358_U248 = ~(P1_R2358_U193 & P1_R2358_U205); 
assign P1_R2358_U489 = ~(P1_U2352 & P1_R2358_U164); 
assign P1_R2358_U496 = ~(P1_U2352 & P1_R2358_U164); 
assign P1_R2358_U596 = ~(P1_R2358_U346 & P1_R2358_U193); 
assign P1_R2358_U611 = ~(P1_R2358_U331 & P1_R2358_U23); 
assign P1_LT_589_U6 = P1_LT_589_U8 | P1_U2673; 
assign P1_R2099_U16 = ~(P1_R2099_U170 & P1_R2099_U54); 
assign P1_R2099_U325 = ~(P1_R2099_U255 & P1_R2099_U170); 
assign P1_R2337_U42 = ~(P1_R2337_U111 & P1_PHYADDRPOINTER_REG_20__SCAN_IN); 
assign P1_R2337_U162 = ~(P1_R2337_U111 & P1_R2337_U41); 
assign P1_R2096_U42 = ~(P1_R2096_U111 & P1_REIP_REG_20__SCAN_IN); 
assign P1_R2096_U162 = ~(P1_R2096_U111 & P1_R2096_U41); 
assign P1_LT_563_U6 = P1_LT_563_U27 & P1_LT_563_U26; 
assign P1_ADD_405_U42 = ~(P1_ADD_405_U114 & P1_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P1_ADD_405_U138 = ~(P1_ADD_405_U114 & P1_ADD_405_U41); 
assign P1_ADD_515_U42 = ~(P1_ADD_515_U111 & P1_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P1_ADD_515_U136 = ~(P1_ADD_515_U111 & P1_ADD_515_U41); 
assign P3_U2818 = ~(P3_U6502 & P3_U6501 & P3_U6504 & P3_U6503 & P3_U3966); 
assign P3_U2852 = ~(P3_U5895 & P3_U5893 & P3_U5894); 
assign P3_U2853 = ~(P3_U5871 & P3_U5869 & P3_U5870); 
assign P3_U3795 = P3_U3794 & P3_U3793 & P3_U5963; 
assign P3_U3826 = P3_U6068 & P3_U6067; 
assign P3_U3828 = P3_U6070 & P3_U6069 & P3_U6071 & P3_U3827; 
assign P3_U3830 = P3_U6082 & P3_U6081 & P3_U6080 & P3_U6079; 
assign P3_U3834 = P3_U6097 & P3_U6096; 
assign P3_U3835 = P3_U6099 & P3_U6098 & P3_U6100 & P3_U6102 & P3_U6101; 
assign P3_U3967 = P3_U6516 & P3_U6513 & P3_U6514 & P3_U6515; 
assign P3_U4096 = P3_U7261 & P3_U4316 & P3_U7262; 
assign P3_U4625 = ~P3_U3120; 
assign P3_U4639 = ~(P3_U2390 & P3_U3120); 
assign P3_U5918 = ~(P3_U4318 & P3_U5916); 
assign P3_U5940 = ~(P3_U3785 & P3_U5922 & P3_U5921 & P3_U3782 & P3_U3788); 
assign P3_U5968 = ~(P3_ADD_360_1242_U83 & P3_U2395); 
assign P3_U6016 = ~(P3_ADD_360_1242_U82 & P3_U2395); 
assign P3_U6017 = ~(P3_SUB_357_1258_U88 & P3_U2393); 
assign P3_U6519 = ~(P3_U2396 & P3_ADD_360_1242_U83); 
assign P3_U6535 = ~(P3_U2396 & P3_ADD_360_1242_U82); 
assign P3_U6536 = ~(P3_U2394 & P3_SUB_357_1258_U88); 
assign P2_U2367 = P2_U2364 & P2_U4417; 
assign P2_U2369 = P2_U2364 & P2_U4428; 
assign P2_U2375 = P2_U4441 & P2_U3521; 
assign P2_U2379 = P2_U4440 & P2_U7865; 
assign P2_U2380 = P2_U4441 & P2_U7865; 
assign P2_U2393 = P2_U4440 & P2_U3521; 
assign P2_U2397 = P2_U4441 & P2_U4601; 
assign P2_U2407 = U298 & P2_U2362; 
assign P2_U2408 = U307 & P2_U2362; 
assign P2_U2409 = U297 & P2_U2362; 
assign P2_U2410 = U306 & P2_U2362; 
assign P2_U2411 = U296 & P2_U2362; 
assign P2_U2412 = U305 & P2_U2362; 
assign P2_U2413 = U295 & P2_U2362; 
assign P2_U2414 = U304 & P2_U2362; 
assign P2_U2415 = U294 & P2_U2362; 
assign P2_U2416 = U302 & P2_U2362; 
assign P2_U2417 = U293 & P2_U2362; 
assign P2_U2418 = U301 & P2_U2362; 
assign P2_U2419 = U291 & P2_U2362; 
assign P2_U2420 = U300 & P2_U2362; 
assign P2_U2421 = U290 & P2_U2362; 
assign P2_U2422 = U299 & P2_U2362; 
assign P2_U2423 = P2_U2365 & P2_U3255; 
assign P2_U2424 = P2_U2365 & P2_U3278; 
assign P2_U2425 = P2_U2365 & P2_U3521; 
assign P2_U2426 = P2_U2365 & P2_U3279; 
assign P2_U2428 = P2_U2365 & P2_U2616; 
assign P2_U2429 = P2_U2365 & P2_U2617; 
assign P2_U2431 = P2_U2365 & P2_U3253; 
assign P2_U2432 = P2_U2365 & P2_U3280; 
assign P2_U2437 = P2_U2364 & P2_U7871; 
assign P2_U2461 = P2_U3579 & P2_U3426; 
assign P2_U2481 = P2_U8064 & P2_U3426; 
assign P2_U2810 = P2_U3242 & P2_R2267_U6; 
assign P2_U2814 = ~(P2_U4190 & P2_U6861); 
assign P2_U2920 = P2_U6232 & P2_DATAO_REG_31__SCAN_IN; 
assign P2_U3670 = ~(P2_U8396 & P2_U8395); 
assign P2_U4394 = ~(P2_U3872 & P2_U5582); 
assign P2_U4400 = ~(P2_U2374 & P2_U3291); 
assign P2_U4600 = ~P2_U3291; 
assign P2_U4640 = ~P2_U3426; 
assign P2_U5646 = ~(P2_U3426 & P2_U5645); 
assign P2_U5652 = ~(P2_U2398 & P2_U8109); 
assign P2_U6233 = ~(P2_U2430 & P2_EAX_REG_0__SCAN_IN); 
assign P2_U6234 = ~(P2_U2396 & P2_LWORD_REG_0__SCAN_IN); 
assign P2_U6235 = ~(P2_U6232 & P2_DATAO_REG_0__SCAN_IN); 
assign P2_U6236 = ~(P2_U2430 & P2_EAX_REG_1__SCAN_IN); 
assign P2_U6237 = ~(P2_U2396 & P2_LWORD_REG_1__SCAN_IN); 
assign P2_U6238 = ~(P2_U6232 & P2_DATAO_REG_1__SCAN_IN); 
assign P2_U6239 = ~(P2_U2430 & P2_EAX_REG_2__SCAN_IN); 
assign P2_U6240 = ~(P2_U2396 & P2_LWORD_REG_2__SCAN_IN); 
assign P2_U6241 = ~(P2_U6232 & P2_DATAO_REG_2__SCAN_IN); 
assign P2_U6242 = ~(P2_U2430 & P2_EAX_REG_3__SCAN_IN); 
assign P2_U6243 = ~(P2_U2396 & P2_LWORD_REG_3__SCAN_IN); 
assign P2_U6244 = ~(P2_U6232 & P2_DATAO_REG_3__SCAN_IN); 
assign P2_U6245 = ~(P2_U2430 & P2_EAX_REG_4__SCAN_IN); 
assign P2_U6246 = ~(P2_U2396 & P2_LWORD_REG_4__SCAN_IN); 
assign P2_U6247 = ~(P2_U6232 & P2_DATAO_REG_4__SCAN_IN); 
assign P2_U6248 = ~(P2_U2430 & P2_EAX_REG_5__SCAN_IN); 
assign P2_U6249 = ~(P2_U2396 & P2_LWORD_REG_5__SCAN_IN); 
assign P2_U6250 = ~(P2_U6232 & P2_DATAO_REG_5__SCAN_IN); 
assign P2_U6251 = ~(P2_U2430 & P2_EAX_REG_6__SCAN_IN); 
assign P2_U6252 = ~(P2_U2396 & P2_LWORD_REG_6__SCAN_IN); 
assign P2_U6253 = ~(P2_U6232 & P2_DATAO_REG_6__SCAN_IN); 
assign P2_U6254 = ~(P2_U2430 & P2_EAX_REG_7__SCAN_IN); 
assign P2_U6255 = ~(P2_U2396 & P2_LWORD_REG_7__SCAN_IN); 
assign P2_U6256 = ~(P2_U6232 & P2_DATAO_REG_7__SCAN_IN); 
assign P2_U6257 = ~(P2_U2430 & P2_EAX_REG_8__SCAN_IN); 
assign P2_U6258 = ~(P2_U2396 & P2_LWORD_REG_8__SCAN_IN); 
assign P2_U6259 = ~(P2_U6232 & P2_DATAO_REG_8__SCAN_IN); 
assign P2_U6260 = ~(P2_U2430 & P2_EAX_REG_9__SCAN_IN); 
assign P2_U6261 = ~(P2_U2396 & P2_LWORD_REG_9__SCAN_IN); 
assign P2_U6262 = ~(P2_U6232 & P2_DATAO_REG_9__SCAN_IN); 
assign P2_U6263 = ~(P2_U2430 & P2_EAX_REG_10__SCAN_IN); 
assign P2_U6264 = ~(P2_U2396 & P2_LWORD_REG_10__SCAN_IN); 
assign P2_U6265 = ~(P2_U6232 & P2_DATAO_REG_10__SCAN_IN); 
assign P2_U6266 = ~(P2_U2430 & P2_EAX_REG_11__SCAN_IN); 
assign P2_U6267 = ~(P2_U2396 & P2_LWORD_REG_11__SCAN_IN); 
assign P2_U6268 = ~(P2_U6232 & P2_DATAO_REG_11__SCAN_IN); 
assign P2_U6269 = ~(P2_U2430 & P2_EAX_REG_12__SCAN_IN); 
assign P2_U6270 = ~(P2_U2396 & P2_LWORD_REG_12__SCAN_IN); 
assign P2_U6271 = ~(P2_U6232 & P2_DATAO_REG_12__SCAN_IN); 
assign P2_U6272 = ~(P2_U2430 & P2_EAX_REG_13__SCAN_IN); 
assign P2_U6273 = ~(P2_U2396 & P2_LWORD_REG_13__SCAN_IN); 
assign P2_U6274 = ~(P2_U6232 & P2_DATAO_REG_13__SCAN_IN); 
assign P2_U6275 = ~(P2_U2430 & P2_EAX_REG_14__SCAN_IN); 
assign P2_U6276 = ~(P2_U2396 & P2_LWORD_REG_14__SCAN_IN); 
assign P2_U6277 = ~(P2_U6232 & P2_DATAO_REG_14__SCAN_IN); 
assign P2_U6278 = ~(P2_U2430 & P2_EAX_REG_15__SCAN_IN); 
assign P2_U6279 = ~(P2_U2396 & P2_LWORD_REG_15__SCAN_IN); 
assign P2_U6280 = ~(P2_U6232 & P2_DATAO_REG_15__SCAN_IN); 
assign P2_U6281 = ~(P2_U2435 & P2_EAX_REG_16__SCAN_IN); 
assign P2_U6282 = ~(P2_U2396 & P2_UWORD_REG_0__SCAN_IN); 
assign P2_U6283 = ~(P2_U6232 & P2_DATAO_REG_16__SCAN_IN); 
assign P2_U6284 = ~(P2_U2435 & P2_EAX_REG_17__SCAN_IN); 
assign P2_U6285 = ~(P2_U2396 & P2_UWORD_REG_1__SCAN_IN); 
assign P2_U6286 = ~(P2_U6232 & P2_DATAO_REG_17__SCAN_IN); 
assign P2_U6287 = ~(P2_U2435 & P2_EAX_REG_18__SCAN_IN); 
assign P2_U6288 = ~(P2_U2396 & P2_UWORD_REG_2__SCAN_IN); 
assign P2_U6289 = ~(P2_U6232 & P2_DATAO_REG_18__SCAN_IN); 
assign P2_U6290 = ~(P2_U2435 & P2_EAX_REG_19__SCAN_IN); 
assign P2_U6291 = ~(P2_U2396 & P2_UWORD_REG_3__SCAN_IN); 
assign P2_U6292 = ~(P2_U6232 & P2_DATAO_REG_19__SCAN_IN); 
assign P2_U6293 = ~(P2_U2435 & P2_EAX_REG_20__SCAN_IN); 
assign P2_U6294 = ~(P2_U2396 & P2_UWORD_REG_4__SCAN_IN); 
assign P2_U6295 = ~(P2_U6232 & P2_DATAO_REG_20__SCAN_IN); 
assign P2_U6296 = ~(P2_U2435 & P2_EAX_REG_21__SCAN_IN); 
assign P2_U6297 = ~(P2_U2396 & P2_UWORD_REG_5__SCAN_IN); 
assign P2_U6298 = ~(P2_U6232 & P2_DATAO_REG_21__SCAN_IN); 
assign P2_U6299 = ~(P2_U2435 & P2_EAX_REG_22__SCAN_IN); 
assign P2_U6300 = ~(P2_U2396 & P2_UWORD_REG_6__SCAN_IN); 
assign P2_U6301 = ~(P2_U6232 & P2_DATAO_REG_22__SCAN_IN); 
assign P2_U6302 = ~(P2_U2435 & P2_EAX_REG_23__SCAN_IN); 
assign P2_U6303 = ~(P2_U2396 & P2_UWORD_REG_7__SCAN_IN); 
assign P2_U6304 = ~(P2_U6232 & P2_DATAO_REG_23__SCAN_IN); 
assign P2_U6305 = ~(P2_U2435 & P2_EAX_REG_24__SCAN_IN); 
assign P2_U6306 = ~(P2_U2396 & P2_UWORD_REG_8__SCAN_IN); 
assign P2_U6307 = ~(P2_U6232 & P2_DATAO_REG_24__SCAN_IN); 
assign P2_U6308 = ~(P2_U2435 & P2_EAX_REG_25__SCAN_IN); 
assign P2_U6309 = ~(P2_U2396 & P2_UWORD_REG_9__SCAN_IN); 
assign P2_U6310 = ~(P2_U6232 & P2_DATAO_REG_25__SCAN_IN); 
assign P2_U6311 = ~(P2_U2435 & P2_EAX_REG_26__SCAN_IN); 
assign P2_U6312 = ~(P2_U2396 & P2_UWORD_REG_10__SCAN_IN); 
assign P2_U6313 = ~(P2_U6232 & P2_DATAO_REG_26__SCAN_IN); 
assign P2_U6314 = ~(P2_U2435 & P2_EAX_REG_27__SCAN_IN); 
assign P2_U6315 = ~(P2_U2396 & P2_UWORD_REG_11__SCAN_IN); 
assign P2_U6316 = ~(P2_U6232 & P2_DATAO_REG_27__SCAN_IN); 
assign P2_U6317 = ~(P2_U2435 & P2_EAX_REG_28__SCAN_IN); 
assign P2_U6318 = ~(P2_U2396 & P2_UWORD_REG_12__SCAN_IN); 
assign P2_U6319 = ~(P2_U6232 & P2_DATAO_REG_28__SCAN_IN); 
assign P2_U6320 = ~(P2_U2435 & P2_EAX_REG_29__SCAN_IN); 
assign P2_U6321 = ~(P2_U2396 & P2_UWORD_REG_13__SCAN_IN); 
assign P2_U6322 = ~(P2_U6232 & P2_DATAO_REG_29__SCAN_IN); 
assign P2_U6323 = ~(P2_U2435 & P2_EAX_REG_30__SCAN_IN); 
assign P2_U6324 = ~(P2_U2396 & P2_UWORD_REG_14__SCAN_IN); 
assign P2_U6325 = ~(P2_U6232 & P2_DATAO_REG_30__SCAN_IN); 
assign P2_U6580 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_0__SCAN_IN); 
assign P2_U6581 = ~(P2_U6570 & P2_REIP_REG_0__SCAN_IN); 
assign P2_U6589 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_1__SCAN_IN); 
assign P2_U6590 = ~(P2_U6570 & P2_REIP_REG_1__SCAN_IN); 
assign P2_U6598 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_2__SCAN_IN); 
assign P2_U6599 = ~(P2_U6570 & P2_REIP_REG_2__SCAN_IN); 
assign P2_U6607 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_3__SCAN_IN); 
assign P2_U6608 = ~(P2_U6570 & P2_REIP_REG_3__SCAN_IN); 
assign P2_U6616 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_4__SCAN_IN); 
assign P2_U6617 = ~(P2_U6570 & P2_REIP_REG_4__SCAN_IN); 
assign P2_U6625 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_5__SCAN_IN); 
assign P2_U6626 = ~(P2_U6570 & P2_REIP_REG_5__SCAN_IN); 
assign P2_U6633 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_6__SCAN_IN); 
assign P2_U6634 = ~(P2_U6570 & P2_REIP_REG_6__SCAN_IN); 
assign P2_U6641 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_7__SCAN_IN); 
assign P2_U6642 = ~(P2_U6570 & P2_REIP_REG_7__SCAN_IN); 
assign P2_U6649 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_8__SCAN_IN); 
assign P2_U6650 = ~(P2_U6570 & P2_REIP_REG_8__SCAN_IN); 
assign P2_U6657 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_9__SCAN_IN); 
assign P2_U6658 = ~(P2_U6570 & P2_REIP_REG_9__SCAN_IN); 
assign P2_U6665 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_10__SCAN_IN); 
assign P2_U6666 = ~(P2_U6570 & P2_REIP_REG_10__SCAN_IN); 
assign P2_U6673 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_11__SCAN_IN); 
assign P2_U6674 = ~(P2_U6570 & P2_REIP_REG_11__SCAN_IN); 
assign P2_U6681 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_12__SCAN_IN); 
assign P2_U6682 = ~(P2_U6570 & P2_REIP_REG_12__SCAN_IN); 
assign P2_U6689 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_13__SCAN_IN); 
assign P2_U6690 = ~(P2_U6570 & P2_REIP_REG_13__SCAN_IN); 
assign P2_U6697 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_14__SCAN_IN); 
assign P2_U6698 = ~(P2_U6570 & P2_REIP_REG_14__SCAN_IN); 
assign P2_U6705 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_15__SCAN_IN); 
assign P2_U6706 = ~(P2_U6570 & P2_REIP_REG_15__SCAN_IN); 
assign P2_U6713 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_16__SCAN_IN); 
assign P2_U6714 = ~(P2_U6570 & P2_REIP_REG_16__SCAN_IN); 
assign P2_U6721 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_17__SCAN_IN); 
assign P2_U6722 = ~(P2_U6570 & P2_REIP_REG_17__SCAN_IN); 
assign P2_U6729 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_18__SCAN_IN); 
assign P2_U6730 = ~(P2_U6570 & P2_REIP_REG_18__SCAN_IN); 
assign P2_U6737 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_19__SCAN_IN); 
assign P2_U6738 = ~(P2_U6570 & P2_REIP_REG_19__SCAN_IN); 
assign P2_U6745 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_20__SCAN_IN); 
assign P2_U6746 = ~(P2_U6570 & P2_REIP_REG_20__SCAN_IN); 
assign P2_U6753 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_21__SCAN_IN); 
assign P2_U6754 = ~(P2_U6570 & P2_REIP_REG_21__SCAN_IN); 
assign P2_U6761 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_22__SCAN_IN); 
assign P2_U6762 = ~(P2_U6570 & P2_REIP_REG_22__SCAN_IN); 
assign P2_U6769 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_23__SCAN_IN); 
assign P2_U6770 = ~(P2_U6570 & P2_REIP_REG_23__SCAN_IN); 
assign P2_U6777 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_24__SCAN_IN); 
assign P2_U6778 = ~(P2_U6570 & P2_REIP_REG_24__SCAN_IN); 
assign P2_U6785 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_25__SCAN_IN); 
assign P2_U6786 = ~(P2_U6570 & P2_REIP_REG_25__SCAN_IN); 
assign P2_U6793 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_26__SCAN_IN); 
assign P2_U6794 = ~(P2_U6570 & P2_REIP_REG_26__SCAN_IN); 
assign P2_U6801 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_27__SCAN_IN); 
assign P2_U6802 = ~(P2_U6570 & P2_REIP_REG_27__SCAN_IN); 
assign P2_U6809 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_28__SCAN_IN); 
assign P2_U6810 = ~(P2_U6570 & P2_REIP_REG_28__SCAN_IN); 
assign P2_U6817 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_29__SCAN_IN); 
assign P2_U6818 = ~(P2_U6570 & P2_REIP_REG_29__SCAN_IN); 
assign P2_U6825 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_30__SCAN_IN); 
assign P2_U6826 = ~(P2_U6570 & P2_REIP_REG_30__SCAN_IN); 
assign P2_U6833 = ~(P2_U2378 & P2_PHYADDRPOINTER_REG_31__SCAN_IN); 
assign P2_U6834 = ~(P2_U6570 & P2_REIP_REG_31__SCAN_IN); 
assign P2_U6854 = ~(P2_U6853 & P2_CODEFETCH_REG_SCAN_IN); 
assign P2_U8137 = ~(P2_U6843 & P2_REQUESTPENDING_REG_SCAN_IN); 
assign P2_U8143 = ~(P2_U6857 & P2_READREQUEST_REG_SCAN_IN); 
assign P2_U8288 = ~(P2_U5581 & P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P2_U8289 = ~(P2_U5581 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8291 = ~(P2_U5581 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P2_U8293 = ~(P2_U5581 & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P2_U8295 = ~(P2_U5581 & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U2491 = P1_U4529 & P1_U4528; 
assign P1_U2493 = P1_U4529 & P1_U4524; 
assign P1_U2495 = P1_U4529 & P1_U4525; 
assign P1_U2497 = P1_U4529 & P1_U2486; 
assign P1_U2501 = P1_U4524 & P1_U2474; 
assign P1_U2503 = P1_U4525 & P1_U2474; 
assign P1_U2505 = P1_U2486 & P1_U2474; 
assign P1_U2644 = P1_R2144_U9 & P1_U6746; 
assign P1_U2793 = ~(P1_U6874 & P1_U6873); 
assign P1_U2795 = ~(P1_U6878 & P1_U6877); 
assign P1_U2796 = ~(P1_U6880 & P1_U6879); 
assign P1_U3293 = ~(P1_U4178 & P1_U4509 & P1_U7626 & P1_U4225 & P1_LT_563_U6); 
assign P1_U3357 = ~(P1_U2474 & P1_U4528); 
assign P1_U3403 = ~P1_LT_589_U6; 
assign P1_U3823 = P1_U5704 & P1_U5706; 
assign P1_U3825 = P1_U3824 & P1_U5707; 
assign P1_U3920 = P1_U4227 & P1_U6494; 
assign P1_U3922 = P1_U4227 & P1_U6501; 
assign P1_U3924 = P1_U4227 & P1_U6508; 
assign P1_U4022 = P1_U6826 & P1_U6827 & P1_U6828; 
assign P1_U4561 = ~(P1_U2413 & P1_U2477); 
assign P1_U4566 = ~(P1_U2411 & P1_U2477); 
assign P1_U4571 = ~(P1_U2409 & P1_U2477); 
assign P1_U4576 = ~(P1_U2407 & P1_U2477); 
assign P1_U4581 = ~(P1_U2405 & P1_U2477); 
assign P1_U4586 = ~(P1_U2403 & P1_U2477); 
assign P1_U4591 = ~(P1_U2401 & P1_U2477); 
assign P1_U4596 = ~(P1_U2399 & P1_U2477); 
assign P1_U4619 = ~(P1_U2481 & P1_U2413); 
assign P1_U4624 = ~(P1_U2481 & P1_U2411); 
assign P1_U4629 = ~(P1_U2481 & P1_U2409); 
assign P1_U4634 = ~(P1_U2481 & P1_U2407); 
assign P1_U4639 = ~(P1_U2481 & P1_U2405); 
assign P1_U4644 = ~(P1_U2481 & P1_U2403); 
assign P1_U4649 = ~(P1_U2481 & P1_U2401); 
assign P1_U4654 = ~(P1_U2481 & P1_U2399); 
assign P1_U4658 = ~P1_U3333; 
assign P1_U4678 = ~(P1_U2483 & P1_U2413); 
assign P1_U4683 = ~(P1_U2483 & P1_U2411); 
assign P1_U4688 = ~(P1_U2483 & P1_U2409); 
assign P1_U4693 = ~(P1_U2483 & P1_U2407); 
assign P1_U4698 = ~(P1_U2483 & P1_U2405); 
assign P1_U4703 = ~(P1_U2483 & P1_U2403); 
assign P1_U4708 = ~(P1_U2483 & P1_U2401); 
assign P1_U4713 = ~(P1_U2483 & P1_U2399); 
assign P1_U4735 = ~(P1_U2487 & P1_U2413); 
assign P1_U4740 = ~(P1_U2487 & P1_U2411); 
assign P1_U4745 = ~(P1_U2487 & P1_U2409); 
assign P1_U4750 = ~(P1_U2487 & P1_U2407); 
assign P1_U4755 = ~(P1_U2487 & P1_U2405); 
assign P1_U4760 = ~(P1_U2487 & P1_U2403); 
assign P1_U4765 = ~(P1_U2487 & P1_U2401); 
assign P1_U4770 = ~(P1_U2487 & P1_U2399); 
assign P1_U4780 = ~(P1_U4529 & P1_U4528); 
assign P1_U4837 = ~(P1_U4529 & P1_U4524); 
assign P1_U4895 = ~(P1_U4529 & P1_U4525); 
assign P1_U4952 = ~(P1_U4529 & P1_U2486); 
assign P1_U5065 = ~(P1_U4524 & P1_U2474); 
assign P1_U5123 = ~(P1_U4525 & P1_U2474); 
assign P1_U5180 = ~(P1_U2486 & P1_U2474); 
assign P1_U5251 = ~(P1_U2509 & P1_U2413); 
assign P1_U5256 = ~(P1_U2509 & P1_U2411); 
assign P1_U5261 = ~(P1_U2509 & P1_U2409); 
assign P1_U5266 = ~(P1_U2509 & P1_U2407); 
assign P1_U5271 = ~(P1_U2509 & P1_U2405); 
assign P1_U5276 = ~(P1_U2509 & P1_U2403); 
assign P1_U5281 = ~(P1_U2509 & P1_U2401); 
assign P1_U5286 = ~(P1_U2509 & P1_U2399); 
assign P1_U5308 = ~(P1_U2512 & P1_U2413); 
assign P1_U5313 = ~(P1_U2512 & P1_U2411); 
assign P1_U5318 = ~(P1_U2512 & P1_U2409); 
assign P1_U5323 = ~(P1_U2512 & P1_U2407); 
assign P1_U5328 = ~(P1_U2512 & P1_U2405); 
assign P1_U5333 = ~(P1_U2512 & P1_U2403); 
assign P1_U5338 = ~(P1_U2512 & P1_U2401); 
assign P1_U5343 = ~(P1_U2512 & P1_U2399); 
assign P1_U5366 = ~(P1_U2514 & P1_U2413); 
assign P1_U5371 = ~(P1_U2514 & P1_U2411); 
assign P1_U5376 = ~(P1_U2514 & P1_U2409); 
assign P1_U5381 = ~(P1_U2514 & P1_U2407); 
assign P1_U5386 = ~(P1_U2514 & P1_U2405); 
assign P1_U5391 = ~(P1_U2514 & P1_U2403); 
assign P1_U5396 = ~(P1_U2514 & P1_U2401); 
assign P1_U5401 = ~(P1_U2514 & P1_U2399); 
assign P1_U5423 = ~(P1_U2516 & P1_U2413); 
assign P1_U5428 = ~(P1_U2516 & P1_U2411); 
assign P1_U5433 = ~(P1_U2516 & P1_U2409); 
assign P1_U5438 = ~(P1_U2516 & P1_U2407); 
assign P1_U5442 = ~(P1_U2516 & P1_U2405); 
assign P1_U5447 = ~(P1_U2516 & P1_U2403); 
assign P1_U5452 = ~(P1_U2516 & P1_U2401); 
assign P1_U5457 = ~(P1_U2516 & P1_U2399); 
assign P1_U5536 = ~(P1_U2428 & P1_LT_589_U6 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U5539 = ~(P1_U4527 & P1_U3454); 
assign P1_U5550 = ~(P1_U3326 & P1_U3333); 
assign P1_U6875 = ~(P1_U4159 & P1_R2144_U9); 
assign P1_U7693 = ~P1_U3454; 
assign P1_U7732 = ~(P1_U3454 & P1_U3314); 
assign P3_ADD_476_U81 = ~(P3_ADD_476_U162 & P3_ADD_476_U161); 
assign P3_ADD_476_U112 = ~P3_ADD_476_U42; 
assign P3_ADD_476_U159 = ~(P3_ADD_476_U42 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_531_U86 = ~(P3_ADD_531_U171 & P3_ADD_531_U170); 
assign P3_ADD_531_U116 = ~P3_ADD_531_U43; 
assign P3_ADD_531_U166 = ~(P3_ADD_531_U43 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_SUB_320_U115 = ~(P3_SUB_320_U97 & P3_SUB_320_U73); 
assign P3_SUB_320_U151 = ~(P3_SUB_320_U97 & P3_SUB_320_U73); 
assign P3_ADD_318_U81 = ~(P3_ADD_318_U162 & P3_ADD_318_U161); 
assign P3_ADD_318_U112 = ~P3_ADD_318_U42; 
assign P3_ADD_318_U159 = ~(P3_ADD_318_U42 & P3_PHYADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_315_U77 = ~(P3_ADD_315_U154 & P3_ADD_315_U153); 
assign P3_ADD_315_U109 = ~P3_ADD_315_U42; 
assign P3_ADD_315_U151 = ~(P3_ADD_315_U42 & P3_PHYADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_360_1242_U7 = P3_ADD_360_1242_U181 & P3_ADD_360_1242_U50; 
assign P3_ADD_360_1242_U8 = P3_ADD_360_1242_U179 & P3_ADD_360_1242_U53; 
assign P3_ADD_360_1242_U56 = ~(P3_ADD_360_1242_U101 & P3_ADD_360_1242_U157); 
assign P3_ADD_360_1242_U176 = ~(P3_ADD_360_1242_U157 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_360_1242_U250 = ~(P3_ADD_360_1242_U157 & P3_ADD_360_1242_U54); 
assign P3_ADD_467_U81 = ~(P3_ADD_467_U162 & P3_ADD_467_U161); 
assign P3_ADD_467_U112 = ~P3_ADD_467_U42; 
assign P3_ADD_467_U159 = ~(P3_ADD_467_U42 & P3_REIP_REG_21__SCAN_IN); 
assign P3_ADD_430_U81 = ~(P3_ADD_430_U162 & P3_ADD_430_U161); 
assign P3_ADD_430_U112 = ~P3_ADD_430_U42; 
assign P3_ADD_430_U159 = ~(P3_ADD_430_U42 & P3_REIP_REG_21__SCAN_IN); 
assign P3_ADD_380_U86 = ~(P3_ADD_380_U171 & P3_ADD_380_U170); 
assign P3_ADD_380_U116 = ~P3_ADD_380_U43; 
assign P3_ADD_380_U166 = ~(P3_ADD_380_U43 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_344_U86 = ~(P3_ADD_344_U171 & P3_ADD_344_U170); 
assign P3_ADD_344_U116 = ~P3_ADD_344_U43; 
assign P3_ADD_344_U166 = ~(P3_ADD_344_U43 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_339_U81 = ~(P3_ADD_339_U162 & P3_ADD_339_U161); 
assign P3_ADD_339_U112 = ~P3_ADD_339_U42; 
assign P3_ADD_339_U159 = ~(P3_ADD_339_U42 & P3_PHYADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_541_U81 = ~(P3_ADD_541_U162 & P3_ADD_541_U161); 
assign P3_ADD_541_U112 = ~P3_ADD_541_U42; 
assign P3_ADD_541_U159 = ~(P3_ADD_541_U42 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_SUB_357_1258_U63 = ~(P3_SUB_357_1258_U104 & P3_SUB_357_1258_U284); 
assign P3_SUB_357_1258_U64 = ~(P3_SUB_357_1258_U276 & P3_SUB_357_1258_U205); 
assign P3_SUB_357_1258_U133 = ~(P3_SUB_357_1258_U282 & P3_SUB_357_1258_U14); 
assign P3_SUB_357_1258_U135 = ~(P3_SUB_357_1258_U280 & P3_SUB_357_1258_U12); 
assign P3_SUB_357_1258_U137 = ~(P3_SUB_357_1258_U278 & P3_SUB_357_1258_U10); 
assign P3_SUB_357_1258_U248 = ~(P3_SUB_357_1258_U440 & P3_SUB_357_1258_U439 & P3_SUB_357_1258_U247); 
assign P3_SUB_357_1258_U438 = ~(P3_SUB_357_1258_U203 & P3_SUB_357_1258_U436); 
assign P3_ADD_515_U81 = ~(P3_ADD_515_U162 & P3_ADD_515_U161); 
assign P3_ADD_515_U112 = ~P3_ADD_515_U42; 
assign P3_ADD_515_U159 = ~(P3_ADD_515_U42 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_394_U80 = ~(P3_ADD_394_U164 & P3_ADD_394_U163); 
assign P3_ADD_394_U115 = ~P3_ADD_394_U42; 
assign P3_ADD_394_U161 = ~(P3_ADD_394_U42 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_441_U81 = ~(P3_ADD_441_U162 & P3_ADD_441_U161); 
assign P3_ADD_441_U112 = ~P3_ADD_441_U42; 
assign P3_ADD_441_U159 = ~(P3_ADD_441_U42 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_349_U86 = ~(P3_ADD_349_U171 & P3_ADD_349_U170); 
assign P3_ADD_349_U116 = ~P3_ADD_349_U43; 
assign P3_ADD_349_U166 = ~(P3_ADD_349_U43 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_405_U80 = ~(P3_ADD_405_U164 & P3_ADD_405_U163); 
assign P3_ADD_405_U115 = ~P3_ADD_405_U42; 
assign P3_ADD_405_U161 = ~(P3_ADD_405_U42 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_553_U86 = ~(P3_ADD_553_U171 & P3_ADD_553_U170); 
assign P3_ADD_553_U116 = ~P3_ADD_553_U43; 
assign P3_ADD_553_U166 = ~(P3_ADD_553_U43 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_558_U86 = ~(P3_ADD_558_U171 & P3_ADD_558_U170); 
assign P3_ADD_558_U116 = ~P3_ADD_558_U43; 
assign P3_ADD_558_U166 = ~(P3_ADD_558_U43 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_385_U86 = ~(P3_ADD_385_U171 & P3_ADD_385_U170); 
assign P3_ADD_385_U116 = ~P3_ADD_385_U43; 
assign P3_ADD_385_U166 = ~(P3_ADD_385_U43 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_547_U86 = ~(P3_ADD_547_U171 & P3_ADD_547_U170); 
assign P3_ADD_547_U116 = ~P3_ADD_547_U43; 
assign P3_ADD_547_U166 = ~(P3_ADD_547_U43 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_371_1212_U84 = ~(P3_ADD_371_1212_U259 & P3_ADD_371_1212_U258); 
assign P3_ADD_371_1212_U85 = ~(P3_ADD_371_1212_U261 & P3_ADD_371_1212_U260); 
assign P3_ADD_371_1212_U166 = ~P3_ADD_371_1212_U56; 
assign P3_ADD_371_1212_U189 = ~(P3_ADD_371_1212_U54 & P3_ADD_371_1212_U188); 
assign P3_ADD_371_1212_U191 = ~(P3_ADD_371_1212_U51 & P3_ADD_371_1212_U190); 
assign P3_ADD_371_1212_U256 = ~(P3_ADD_371_1212_U56 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_494_U81 = ~(P3_ADD_494_U162 & P3_ADD_494_U161); 
assign P3_ADD_494_U112 = ~P3_ADD_494_U42; 
assign P3_ADD_494_U159 = ~(P3_ADD_494_U42 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_536_U81 = ~(P3_ADD_536_U162 & P3_ADD_536_U161); 
assign P3_ADD_536_U112 = ~P3_ADD_536_U42; 
assign P3_ADD_536_U159 = ~(P3_ADD_536_U42 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P2_R2099_U27 = ~(P2_U2737 & P2_R2099_U125); 
assign P2_R2099_U223 = ~(P2_R2099_U125 & P2_R2099_U26); 
assign P2_ADD_391_1196_U15 = ~P2_R2182_U73; 
assign P2_ADD_391_1196_U38 = ~(P2_ADD_391_1196_U176 & P2_ADD_391_1196_U175); 
assign P2_ADD_391_1196_U45 = ~P2_R2096_U94; 
assign P2_ADD_391_1196_U91 = ~(P2_ADD_391_1196_U338 & P2_ADD_391_1196_U337); 
assign P2_ADD_391_1196_U161 = ~(P2_R2096_U72 & P2_R2182_U73); 
assign P2_ADD_391_1196_U184 = P2_R2096_U72 | P2_R2182_U73; 
assign P2_ADD_391_1196_U197 = P2_R2182_U73 | P2_R2096_U72; 
assign P2_ADD_391_1196_U202 = P2_R2096_U72 | P2_R2182_U73; 
assign P2_ADD_391_1196_U319 = ~(P2_R2182_U73 & P2_ADD_391_1196_U16); 
assign P2_ADD_391_1196_U323 = ~(P2_R2096_U73 & P2_ADD_391_1196_U17); 
assign P2_ADD_391_1196_U330 = ~(P2_ADD_391_1196_U115 & P2_ADD_391_1196_U116); 
assign P2_ADD_391_1196_U331 = ~(P2_ADD_391_1196_U173 & P2_ADD_391_1196_U329); 
assign P2_R2182_U20 = P2_U2672 & P2_R2182_U19; 
assign P2_R2182_U72 = ~(P2_R2182_U198 & P2_R2182_U197); 
assign P2_R2182_U140 = ~P2_R2182_U19; 
assign P2_R2182_U193 = ~(P2_R2182_U34 & P2_R2182_U19); 
assign P2_R2182_U196 = ~(P2_R2182_U139 & P2_U2673); 
assign P2_R2027_U86 = ~(P2_R2027_U171 & P2_R2027_U170); 
assign P2_R2027_U116 = ~P2_R2027_U43; 
assign P2_R2027_U166 = ~(P2_R2027_U43 & P2_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P2_R2337_U79 = ~(P2_R2337_U160 & P2_R2337_U159); 
assign P2_R2337_U113 = ~P2_R2337_U43; 
assign P2_R2337_U157 = ~(P2_R2337_U43 & P2_PHYADDRPOINTER_REG_22__SCAN_IN); 
assign P2_R2096_U5 = P2_U2633 & P2_R2096_U18; 
assign P2_R2096_U93 = ~(P2_R2096_U255 & P2_R2096_U254); 
assign P2_R2096_U151 = ~P2_R2096_U18; 
assign P2_R2096_U250 = ~(P2_R2096_U34 & P2_R2096_U18); 
assign P2_R2096_U253 = ~(P2_R2096_U150 & P2_U2634); 
assign P2_R2256_U21 = ~(P2_R2256_U70 & P2_R2256_U69); 
assign P2_R2256_U27 = P2_R2256_U58 & P2_R2256_U57; 
assign P2_R2256_U35 = ~(P2_U2616 & P2_R2256_U34); 
assign P2_R2256_U61 = ~(P2_R2256_U60 & P2_R2256_U59); 
assign P2_R2256_U65 = ~(P2_R2256_U45 & P2_U7873); 
assign P2_R2256_U68 = ~(P2_R2256_U32 & P2_U2616); 
assign P2_R1957_U115 = ~(P2_R1957_U97 & P2_R1957_U73); 
assign P2_R1957_U151 = ~(P2_R1957_U97 & P2_R1957_U73); 
assign P2_R2278_U50 = ~P2_U2811; 
assign P2_R2278_U52 = ~(P2_U2811 & P2_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P2_R2278_U238 = P2_U2811 | P2_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P2_R2278_U346 = ~(P2_R2278_U30 & P2_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P2_R2278_U348 = ~(P2_R2278_U30 & P2_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P2_R2278_U555 = ~(P2_U2811 & P2_R2278_U51); 
assign P2_R2278_U557 = ~(P2_U2811 & P2_R2278_U51); 
assign P2_ADD_394_U68 = ~(P2_ADD_394_U138 & P2_ADD_394_U137); 
assign P2_ADD_394_U115 = ~P2_ADD_394_U42; 
assign P2_ADD_394_U177 = ~(P2_ADD_394_U42 & P2_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P2_R2267_U85 = P2_R2267_U164 & P2_R2267_U163; 
assign P2_R2267_U103 = ~P2_R2267_U32; 
assign P2_R2267_U131 = ~(P2_U2784 & P2_R2267_U130); 
assign P2_R2267_U161 = ~(P2_U2783 & P2_R2267_U32); 
assign P1_R2144_U26 = ~(P1_R2144_U65 & P1_R2144_U141); 
assign P1_R2144_U80 = P1_R2144_U211 & P1_R2144_U210; 
assign P1_R2144_U95 = ~(P1_R2144_U141 & P1_R2144_U34); 
assign P1_R2144_U145 = ~P1_R2144_U144; 
assign P1_R2144_U146 = ~(P1_R2144_U101 & P1_R2144_U12); 
assign P1_R2144_U208 = ~(P1_R2144_U122 & P1_R2144_U207); 
assign P1_R2144_U253 = ~(P1_R2144_U231 & P1_R2144_U141); 
assign P1_R2144_U255 = ~(P1_R2144_U140 & P1_R2144_U234); 
assign P1_R2144_U257 = ~(P1_R2144_U139 & P1_R2144_U237); 
assign P1_R2278_U37 = ~P1_U2797; 
assign P1_R2278_U192 = ~(P1_R2278_U213 & P1_R2278_U234); 
assign P1_R2278_U214 = P1_R2278_U559 & P1_R2278_U558; 
assign P1_R2278_U240 = P1_U2797 | P1_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P1_R2278_U242 = ~(P1_U2797 & P1_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P1_R2278_U455 = ~(P1_U2797 & P1_R2278_U36); 
assign P1_R2278_U457 = ~(P1_U2797 & P1_R2278_U36); 
assign P1_R2278_U479 = ~(P1_R2278_U35 & P1_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P1_R2278_U481 = ~(P1_R2278_U35 & P1_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P1_R2358_U24 = ~P1_U2643; 
assign P1_R2358_U26 = ~P1_U2645; 
assign P1_R2358_U27 = ~P1_U2646; 
assign P1_R2358_U28 = ~(P1_U2646 & P1_R2358_U413); 
assign P1_R2358_U65 = ~(P1_R2358_U206 & P1_R2358_U248); 
assign P1_R2358_U76 = ~(P1_R2358_U611 & P1_R2358_U610); 
assign P1_R2358_U165 = ~P1_U2664; 
assign P1_R2358_U202 = ~(P1_R2358_U436 & P1_R2358_U435 & P1_R2358_U30); 
assign P1_R2358_U204 = ~(P1_R2358_U438 & P1_R2358_U437 & P1_R2358_U32); 
assign P1_R2358_U212 = ~(P1_R2358_U211 & P1_R2358_U206 & P1_R2358_U207); 
assign P1_R2358_U216 = ~(P1_U2643 & P1_R2358_U421); 
assign P1_R2358_U220 = ~(P1_U2645 & P1_R2358_U416); 
assign P1_R2358_U492 = ~(P1_U2664 & P1_R2358_U23); 
assign P1_R2358_U494 = ~(P1_U2664 & P1_R2358_U23); 
assign P1_R2358_U498 = ~(P1_R2358_U497 & P1_R2358_U496); 
assign P1_R2358_U597 = ~(P1_R2358_U106 & P1_R2358_U247); 
assign P1_R2099_U76 = ~(P1_R2099_U326 & P1_R2099_U325); 
assign P1_R2099_U171 = ~P1_R2099_U16; 
assign P1_R2099_U317 = ~(P1_R2099_U53 & P1_R2099_U16); 
assign P1_R2337_U81 = ~(P1_R2337_U162 & P1_R2337_U161); 
assign P1_R2337_U112 = ~P1_R2337_U42; 
assign P1_R2337_U159 = ~(P1_R2337_U42 & P1_PHYADDRPOINTER_REG_21__SCAN_IN); 
assign P1_R2096_U81 = ~(P1_R2096_U162 & P1_R2096_U161); 
assign P1_R2096_U112 = ~P1_R2096_U42; 
assign P1_R2096_U159 = ~(P1_R2096_U42 & P1_REIP_REG_21__SCAN_IN); 
assign P1_ADD_405_U68 = ~(P1_ADD_405_U138 & P1_ADD_405_U137); 
assign P1_ADD_405_U115 = ~P1_ADD_405_U42; 
assign P1_ADD_405_U177 = ~(P1_ADD_405_U42 & P1_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P1_ADD_515_U68 = ~(P1_ADD_515_U136 & P1_ADD_515_U135); 
assign P1_ADD_515_U112 = ~P1_ADD_515_U42; 
assign P1_ADD_515_U173 = ~(P1_ADD_515_U42 & P1_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_U2817 = ~(P3_U6510 & P3_U6509 & P3_U6512 & P3_U6511 & P3_U3967); 
assign P3_U2851 = ~(P3_U5919 & P3_U5917 & P3_U5918); 
assign P3_U3367 = P3_U3366 & P3_U4639; 
assign P3_U3799 = P3_U3796 & P3_U5970 & P3_U3798 & P3_U5969 & P3_U5968; 
assign P3_U3812 = P3_U3813 & P3_U6017; 
assign P3_U4627 = ~(P3_U3362 & P3_U4625); 
assign P3_U5942 = ~(P3_U4318 & P3_U5940); 
assign P3_U5964 = ~(P3_U3792 & P3_U5946 & P3_U5945 & P3_U3789 & P3_U3795); 
assign P3_U5987 = ~(P3_ADD_371_1212_U85 & P3_U2360); 
assign P3_U5992 = ~(P3_ADD_360_1242_U7 & P3_U2395); 
assign P3_U6035 = ~(P3_ADD_371_1212_U84 & P3_U2360); 
assign P3_U6040 = ~(P3_ADD_360_1242_U8 & P3_U2395); 
assign P3_U6090 = ~(P3_ADD_558_U86 & P3_U3220); 
assign P3_U6091 = ~(P3_ADD_553_U86 & P3_U4298); 
assign P3_U6092 = ~(P3_ADD_547_U86 & P3_U4299); 
assign P3_U6095 = ~(P3_ADD_531_U86 & P3_U2354); 
assign P3_U6103 = ~(P3_ADD_385_U86 & P3_U2358); 
assign P3_U6104 = ~(P3_ADD_380_U86 & P3_U2359); 
assign P3_U6105 = ~(P3_ADD_349_U86 & P3_U4306); 
assign P3_U6106 = ~(P3_ADD_344_U86 & P3_U2362); 
assign P3_U6117 = ~(P3_ADD_541_U81 & P3_U4300); 
assign P3_U6118 = ~(P3_ADD_536_U81 & P3_U4301); 
assign P3_U6121 = ~(P3_ADD_515_U81 & P3_U4302); 
assign P3_U6122 = ~(P3_ADD_494_U81 & P3_U2356); 
assign P3_U6123 = ~(P3_ADD_476_U81 & P3_U4303); 
assign P3_U6124 = ~(P3_ADD_441_U81 & P3_U4304); 
assign P3_U6125 = ~(P3_ADD_405_U80 & P3_U4305); 
assign P3_U6126 = ~(P3_ADD_394_U80 & P3_U2357); 
assign P3_U6523 = ~(P3_U2387 & P3_ADD_371_1212_U85); 
assign P3_U6527 = ~(P3_U2396 & P3_ADD_360_1242_U7); 
assign P3_U6539 = ~(P3_U2387 & P3_ADD_371_1212_U84); 
assign P3_U6543 = ~(P3_U2396 & P3_ADD_360_1242_U8); 
assign P3_U6565 = ~(P3_ADD_318_U81 & P3_U2398); 
assign P3_U6570 = ~(P3_ADD_339_U81 & P3_U2388); 
assign P3_U6574 = ~(P3_ADD_315_U77 & P3_U2397); 
assign P3_U7270 = ~(P3_ADD_467_U81 & P3_U2601); 
assign P3_U7272 = ~(P3_ADD_430_U81 & P3_U2405); 
assign P2_U2377 = P2_U2367 & P2_U4411; 
assign P2_U2391 = P2_U2369 & P2_U3545; 
assign P2_U2392 = P2_U6571 & P2_U2369; 
assign P2_U2427 = P2_U2375 & P2_U3279; 
assign P2_U2433 = P2_U2375 & P2_U3295; 
assign P2_U2434 = P2_U2375 & P2_U7869; 
assign P2_U2491 = P2_U4640 & P2_U3579; 
assign P2_U2500 = P2_U4640 & P2_U8064; 
assign P2_U2809 = P2_U3242 & P2_R2267_U85; 
assign P2_U2816 = ~(P2_U6855 & P2_U6854); 
assign P2_U2921 = ~(P2_U6324 & P2_U6323 & P2_U6325); 
assign P2_U2922 = ~(P2_U6321 & P2_U6320 & P2_U6322); 
assign P2_U2923 = ~(P2_U6318 & P2_U6317 & P2_U6319); 
assign P2_U2924 = ~(P2_U6315 & P2_U6314 & P2_U6316); 
assign P2_U2925 = ~(P2_U6312 & P2_U6311 & P2_U6313); 
assign P2_U2926 = ~(P2_U6309 & P2_U6308 & P2_U6310); 
assign P2_U2927 = ~(P2_U6306 & P2_U6305 & P2_U6307); 
assign P2_U2928 = ~(P2_U6303 & P2_U6302 & P2_U6304); 
assign P2_U2929 = ~(P2_U6300 & P2_U6299 & P2_U6301); 
assign P2_U2930 = ~(P2_U6297 & P2_U6296 & P2_U6298); 
assign P2_U2931 = ~(P2_U6294 & P2_U6293 & P2_U6295); 
assign P2_U2932 = ~(P2_U6291 & P2_U6290 & P2_U6292); 
assign P2_U2933 = ~(P2_U6288 & P2_U6287 & P2_U6289); 
assign P2_U2934 = ~(P2_U6285 & P2_U6284 & P2_U6286); 
assign P2_U2935 = ~(P2_U6282 & P2_U6281 & P2_U6283); 
assign P2_U2936 = ~(P2_U6279 & P2_U6278 & P2_U6280); 
assign P2_U2937 = ~(P2_U6276 & P2_U6275 & P2_U6277); 
assign P2_U2938 = ~(P2_U6273 & P2_U6272 & P2_U6274); 
assign P2_U2939 = ~(P2_U6270 & P2_U6269 & P2_U6271); 
assign P2_U2940 = ~(P2_U6267 & P2_U6266 & P2_U6268); 
assign P2_U2941 = ~(P2_U6264 & P2_U6263 & P2_U6265); 
assign P2_U2942 = ~(P2_U6261 & P2_U6260 & P2_U6262); 
assign P2_U2943 = ~(P2_U6258 & P2_U6257 & P2_U6259); 
assign P2_U2944 = ~(P2_U6255 & P2_U6254 & P2_U6256); 
assign P2_U2945 = ~(P2_U6252 & P2_U6251 & P2_U6253); 
assign P2_U2946 = ~(P2_U6249 & P2_U6248 & P2_U6250); 
assign P2_U2947 = ~(P2_U6246 & P2_U6245 & P2_U6247); 
assign P2_U2948 = ~(P2_U6243 & P2_U6242 & P2_U6244); 
assign P2_U2949 = ~(P2_U6240 & P2_U6239 & P2_U6241); 
assign P2_U2950 = ~(P2_U6237 & P2_U6236 & P2_U6238); 
assign P2_U2951 = ~(P2_U6234 & P2_U6233 & P2_U6235); 
assign P2_U3320 = ~(P2_U4636 & P2_U2461); 
assign P2_U3339 = ~(P2_U4709 & P2_U2461); 
assign P2_U3354 = ~(P2_U4767 & P2_U2461); 
assign P2_U3366 = ~(P2_U2475 & P2_U2461); 
assign P2_U3379 = ~(P2_U2481 & P2_U4636); 
assign P2_U3391 = ~(P2_U2481 & P2_U4709); 
assign P2_U3402 = ~(P2_U2481 & P2_U4767); 
assign P2_U3414 = ~(P2_U2481 & P2_U2475); 
assign P2_U3610 = ~(P2_U8138 & P2_U8137); 
assign P2_U3612 = ~(P2_U8144 & P2_U8143); 
assign P2_U3617 = ~(P2_U8288 & P2_U8287); 
assign P2_U3618 = ~(P2_U8290 & P2_U8289); 
assign P2_U3619 = ~(P2_U8292 & P2_U8291); 
assign P2_U3620 = ~(P2_U8294 & P2_U8293); 
assign P2_U3621 = ~(P2_U8296 & P2_U8295); 
assign P2_U4073 = P2_U6581 & P2_U6580; 
assign P2_U4077 = P2_U6590 & P2_U6589; 
assign P2_U4081 = P2_U6599 & P2_U6598; 
assign P2_U4085 = P2_U6608 & P2_U6607; 
assign P2_U4088 = P2_U6617 & P2_U6616; 
assign P2_U4092 = P2_U6626 & P2_U6625; 
assign P2_U4096 = P2_U6634 & P2_U6633; 
assign P2_U4099 = P2_U6642 & P2_U6641; 
assign P2_U4102 = P2_U6650 & P2_U6649; 
assign P2_U4105 = P2_U6658 & P2_U6657; 
assign P2_U4108 = P2_U6666 & P2_U6665; 
assign P2_U4111 = P2_U6674 & P2_U6673; 
assign P2_U4114 = P2_U6682 & P2_U6681; 
assign P2_U4117 = P2_U6690 & P2_U6689; 
assign P2_U4120 = P2_U6698 & P2_U6697; 
assign P2_U4123 = P2_U6706 & P2_U6705; 
assign P2_U4127 = P2_U6714 & P2_U6713; 
assign P2_U4131 = P2_U6722 & P2_U6721; 
assign P2_U4135 = P2_U6730 & P2_U6729; 
assign P2_U4139 = P2_U6738 & P2_U6737; 
assign P2_U4142 = P2_U6746 & P2_U6745; 
assign P2_U4145 = P2_U6754 & P2_U6753; 
assign P2_U4147 = P2_U6762 & P2_U6761; 
assign P2_U4151 = P2_U6770 & P2_U6769; 
assign P2_U4154 = P2_U6778 & P2_U6777; 
assign P2_U4155 = P2_U6786 & P2_U6785; 
assign P2_U4157 = P2_U6794 & P2_U6793; 
assign P2_U4159 = P2_U6802 & P2_U6801; 
assign P2_U4161 = P2_U6810 & P2_U6809; 
assign P2_U4163 = P2_U6818 & P2_U6817; 
assign P2_U4165 = P2_U6826 & P2_U6825; 
assign P2_U4167 = P2_U6834 & P2_U6833; 
assign P2_U4448 = ~(P2_U2367 & P2_U3290); 
assign P2_U4669 = ~(P2_U2425 & P2_U4643); 
assign P2_U4670 = ~(P2_U2422 & P2_U2463); 
assign P2_U4674 = ~(P2_U2426 & P2_U4643); 
assign P2_U4675 = ~(P2_U2420 & P2_U2463); 
assign P2_U4679 = ~(P2_U2429 & P2_U4643); 
assign P2_U4680 = ~(P2_U2418 & P2_U2463); 
assign P2_U4684 = ~(P2_U2424 & P2_U4643); 
assign P2_U4685 = ~(P2_U2416 & P2_U2463); 
assign P2_U4689 = ~(P2_U2423 & P2_U4643); 
assign P2_U4690 = ~(P2_U2414 & P2_U2463); 
assign P2_U4694 = ~(P2_U2432 & P2_U4643); 
assign P2_U4695 = ~(P2_U2412 & P2_U2463); 
assign P2_U4699 = ~(P2_U2428 & P2_U4643); 
assign P2_U4700 = ~(P2_U2410 & P2_U2463); 
assign P2_U4704 = ~(P2_U2431 & P2_U4643); 
assign P2_U4705 = ~(P2_U2408 & P2_U2463); 
assign P2_U4727 = ~(P2_U4711 & P2_U2425); 
assign P2_U4728 = ~(P2_U2469 & P2_U2422); 
assign P2_U4732 = ~(P2_U4711 & P2_U2426); 
assign P2_U4733 = ~(P2_U2469 & P2_U2420); 
assign P2_U4737 = ~(P2_U4711 & P2_U2429); 
assign P2_U4738 = ~(P2_U2469 & P2_U2418); 
assign P2_U4742 = ~(P2_U4711 & P2_U2424); 
assign P2_U4743 = ~(P2_U2469 & P2_U2416); 
assign P2_U4747 = ~(P2_U4711 & P2_U2423); 
assign P2_U4748 = ~(P2_U2469 & P2_U2414); 
assign P2_U4752 = ~(P2_U4711 & P2_U2432); 
assign P2_U4753 = ~(P2_U2469 & P2_U2412); 
assign P2_U4757 = ~(P2_U4711 & P2_U2428); 
assign P2_U4758 = ~(P2_U2469 & P2_U2410); 
assign P2_U4762 = ~(P2_U4711 & P2_U2431); 
assign P2_U4763 = ~(P2_U2469 & P2_U2408); 
assign P2_U4786 = ~(P2_U4769 & P2_U2425); 
assign P2_U4787 = ~(P2_U2472 & P2_U2422); 
assign P2_U4791 = ~(P2_U4769 & P2_U2426); 
assign P2_U4792 = ~(P2_U2472 & P2_U2420); 
assign P2_U4796 = ~(P2_U4769 & P2_U2429); 
assign P2_U4797 = ~(P2_U2472 & P2_U2418); 
assign P2_U4801 = ~(P2_U4769 & P2_U2424); 
assign P2_U4802 = ~(P2_U2472 & P2_U2416); 
assign P2_U4806 = ~(P2_U4769 & P2_U2423); 
assign P2_U4807 = ~(P2_U2472 & P2_U2414); 
assign P2_U4811 = ~(P2_U4769 & P2_U2432); 
assign P2_U4812 = ~(P2_U2472 & P2_U2412); 
assign P2_U4816 = ~(P2_U4769 & P2_U2428); 
assign P2_U4817 = ~(P2_U2472 & P2_U2410); 
assign P2_U4821 = ~(P2_U4769 & P2_U2431); 
assign P2_U4822 = ~(P2_U2472 & P2_U2408); 
assign P2_U4843 = ~(P2_U4827 & P2_U2425); 
assign P2_U4844 = ~(P2_U2477 & P2_U2422); 
assign P2_U4848 = ~(P2_U4827 & P2_U2426); 
assign P2_U4849 = ~(P2_U2477 & P2_U2420); 
assign P2_U4853 = ~(P2_U4827 & P2_U2429); 
assign P2_U4854 = ~(P2_U2477 & P2_U2418); 
assign P2_U4858 = ~(P2_U4827 & P2_U2424); 
assign P2_U4859 = ~(P2_U2477 & P2_U2416); 
assign P2_U4863 = ~(P2_U4827 & P2_U2423); 
assign P2_U4864 = ~(P2_U2477 & P2_U2414); 
assign P2_U4868 = ~(P2_U4827 & P2_U2432); 
assign P2_U4869 = ~(P2_U2477 & P2_U2412); 
assign P2_U4873 = ~(P2_U4827 & P2_U2428); 
assign P2_U4874 = ~(P2_U2477 & P2_U2410); 
assign P2_U4878 = ~(P2_U4827 & P2_U2431); 
assign P2_U4879 = ~(P2_U2477 & P2_U2408); 
assign P2_U4901 = ~(P2_U4884 & P2_U2425); 
assign P2_U4902 = ~(P2_U2482 & P2_U2422); 
assign P2_U4906 = ~(P2_U4884 & P2_U2426); 
assign P2_U4907 = ~(P2_U2482 & P2_U2420); 
assign P2_U4911 = ~(P2_U4884 & P2_U2429); 
assign P2_U4912 = ~(P2_U2482 & P2_U2418); 
assign P2_U4916 = ~(P2_U4884 & P2_U2424); 
assign P2_U4917 = ~(P2_U2482 & P2_U2416); 
assign P2_U4921 = ~(P2_U4884 & P2_U2423); 
assign P2_U4922 = ~(P2_U2482 & P2_U2414); 
assign P2_U4926 = ~(P2_U4884 & P2_U2432); 
assign P2_U4927 = ~(P2_U2482 & P2_U2412); 
assign P2_U4931 = ~(P2_U4884 & P2_U2428); 
assign P2_U4932 = ~(P2_U2482 & P2_U2410); 
assign P2_U4936 = ~(P2_U4884 & P2_U2431); 
assign P2_U4937 = ~(P2_U2482 & P2_U2408); 
assign P2_U4958 = ~(P2_U4942 & P2_U2425); 
assign P2_U4959 = ~(P2_U2485 & P2_U2422); 
assign P2_U4963 = ~(P2_U4942 & P2_U2426); 
assign P2_U4964 = ~(P2_U2485 & P2_U2420); 
assign P2_U4968 = ~(P2_U4942 & P2_U2429); 
assign P2_U4969 = ~(P2_U2485 & P2_U2418); 
assign P2_U4973 = ~(P2_U4942 & P2_U2424); 
assign P2_U4974 = ~(P2_U2485 & P2_U2416); 
assign P2_U4978 = ~(P2_U4942 & P2_U2423); 
assign P2_U4979 = ~(P2_U2485 & P2_U2414); 
assign P2_U4983 = ~(P2_U4942 & P2_U2432); 
assign P2_U4984 = ~(P2_U2485 & P2_U2412); 
assign P2_U4988 = ~(P2_U4942 & P2_U2428); 
assign P2_U4989 = ~(P2_U2485 & P2_U2410); 
assign P2_U4993 = ~(P2_U4942 & P2_U2431); 
assign P2_U4994 = ~(P2_U2485 & P2_U2408); 
assign P2_U5016 = ~(P2_U4999 & P2_U2425); 
assign P2_U5017 = ~(P2_U2487 & P2_U2422); 
assign P2_U5021 = ~(P2_U4999 & P2_U2426); 
assign P2_U5022 = ~(P2_U2487 & P2_U2420); 
assign P2_U5026 = ~(P2_U4999 & P2_U2429); 
assign P2_U5027 = ~(P2_U2487 & P2_U2418); 
assign P2_U5031 = ~(P2_U4999 & P2_U2424); 
assign P2_U5032 = ~(P2_U2487 & P2_U2416); 
assign P2_U5036 = ~(P2_U4999 & P2_U2423); 
assign P2_U5037 = ~(P2_U2487 & P2_U2414); 
assign P2_U5041 = ~(P2_U4999 & P2_U2432); 
assign P2_U5042 = ~(P2_U2487 & P2_U2412); 
assign P2_U5046 = ~(P2_U4999 & P2_U2428); 
assign P2_U5047 = ~(P2_U2487 & P2_U2410); 
assign P2_U5051 = ~(P2_U4999 & P2_U2431); 
assign P2_U5052 = ~(P2_U2487 & P2_U2408); 
assign P2_U5073 = ~(P2_U5057 & P2_U2425); 
assign P2_U5074 = ~(P2_U2489 & P2_U2422); 
assign P2_U5078 = ~(P2_U5057 & P2_U2426); 
assign P2_U5079 = ~(P2_U2489 & P2_U2420); 
assign P2_U5083 = ~(P2_U5057 & P2_U2429); 
assign P2_U5084 = ~(P2_U2489 & P2_U2418); 
assign P2_U5088 = ~(P2_U5057 & P2_U2424); 
assign P2_U5089 = ~(P2_U2489 & P2_U2416); 
assign P2_U5093 = ~(P2_U5057 & P2_U2423); 
assign P2_U5094 = ~(P2_U2489 & P2_U2414); 
assign P2_U5098 = ~(P2_U5057 & P2_U2432); 
assign P2_U5099 = ~(P2_U2489 & P2_U2412); 
assign P2_U5103 = ~(P2_U5057 & P2_U2428); 
assign P2_U5104 = ~(P2_U2489 & P2_U2410); 
assign P2_U5108 = ~(P2_U5057 & P2_U2431); 
assign P2_U5109 = ~(P2_U2489 & P2_U2408); 
assign P2_U5129 = ~(P2_U4644 & P2_U2425); 
assign P2_U5130 = ~(P2_U4451 & P2_U2422); 
assign P2_U5134 = ~(P2_U4644 & P2_U2426); 
assign P2_U5135 = ~(P2_U4451 & P2_U2420); 
assign P2_U5139 = ~(P2_U4644 & P2_U2429); 
assign P2_U5140 = ~(P2_U4451 & P2_U2418); 
assign P2_U5144 = ~(P2_U4644 & P2_U2424); 
assign P2_U5145 = ~(P2_U4451 & P2_U2416); 
assign P2_U5149 = ~(P2_U4644 & P2_U2423); 
assign P2_U5150 = ~(P2_U4451 & P2_U2414); 
assign P2_U5154 = ~(P2_U4644 & P2_U2432); 
assign P2_U5155 = ~(P2_U4451 & P2_U2412); 
assign P2_U5159 = ~(P2_U4644 & P2_U2428); 
assign P2_U5160 = ~(P2_U4451 & P2_U2410); 
assign P2_U5164 = ~(P2_U4644 & P2_U2431); 
assign P2_U5165 = ~(P2_U4451 & P2_U2408); 
assign P2_U5186 = ~(P2_U5170 & P2_U2425); 
assign P2_U5187 = ~(P2_U2494 & P2_U2422); 
assign P2_U5191 = ~(P2_U5170 & P2_U2426); 
assign P2_U5192 = ~(P2_U2494 & P2_U2420); 
assign P2_U5196 = ~(P2_U5170 & P2_U2429); 
assign P2_U5197 = ~(P2_U2494 & P2_U2418); 
assign P2_U5201 = ~(P2_U5170 & P2_U2424); 
assign P2_U5202 = ~(P2_U2494 & P2_U2416); 
assign P2_U5206 = ~(P2_U5170 & P2_U2423); 
assign P2_U5207 = ~(P2_U2494 & P2_U2414); 
assign P2_U5211 = ~(P2_U5170 & P2_U2432); 
assign P2_U5212 = ~(P2_U2494 & P2_U2412); 
assign P2_U5216 = ~(P2_U5170 & P2_U2428); 
assign P2_U5217 = ~(P2_U2494 & P2_U2410); 
assign P2_U5221 = ~(P2_U5170 & P2_U2431); 
assign P2_U5222 = ~(P2_U2494 & P2_U2408); 
assign P2_U5244 = ~(P2_U5227 & P2_U2425); 
assign P2_U5245 = ~(P2_U2496 & P2_U2422); 
assign P2_U5249 = ~(P2_U5227 & P2_U2426); 
assign P2_U5250 = ~(P2_U2496 & P2_U2420); 
assign P2_U5254 = ~(P2_U5227 & P2_U2429); 
assign P2_U5255 = ~(P2_U2496 & P2_U2418); 
assign P2_U5259 = ~(P2_U5227 & P2_U2424); 
assign P2_U5260 = ~(P2_U2496 & P2_U2416); 
assign P2_U5264 = ~(P2_U5227 & P2_U2423); 
assign P2_U5265 = ~(P2_U2496 & P2_U2414); 
assign P2_U5269 = ~(P2_U5227 & P2_U2432); 
assign P2_U5270 = ~(P2_U2496 & P2_U2412); 
assign P2_U5274 = ~(P2_U5227 & P2_U2428); 
assign P2_U5275 = ~(P2_U2496 & P2_U2410); 
assign P2_U5279 = ~(P2_U5227 & P2_U2431); 
assign P2_U5280 = ~(P2_U2496 & P2_U2408); 
assign P2_U5301 = ~(P2_U5285 & P2_U2425); 
assign P2_U5302 = ~(P2_U2498 & P2_U2422); 
assign P2_U5306 = ~(P2_U5285 & P2_U2426); 
assign P2_U5307 = ~(P2_U2498 & P2_U2420); 
assign P2_U5311 = ~(P2_U5285 & P2_U2429); 
assign P2_U5312 = ~(P2_U2498 & P2_U2418); 
assign P2_U5316 = ~(P2_U5285 & P2_U2424); 
assign P2_U5317 = ~(P2_U2498 & P2_U2416); 
assign P2_U5321 = ~(P2_U5285 & P2_U2423); 
assign P2_U5322 = ~(P2_U2498 & P2_U2414); 
assign P2_U5326 = ~(P2_U5285 & P2_U2432); 
assign P2_U5327 = ~(P2_U2498 & P2_U2412); 
assign P2_U5331 = ~(P2_U5285 & P2_U2428); 
assign P2_U5332 = ~(P2_U2498 & P2_U2410); 
assign P2_U5336 = ~(P2_U5285 & P2_U2431); 
assign P2_U5337 = ~(P2_U2498 & P2_U2408); 
assign P2_U5359 = ~(P2_U5342 & P2_U2425); 
assign P2_U5360 = ~(P2_U2502 & P2_U2422); 
assign P2_U5364 = ~(P2_U5342 & P2_U2426); 
assign P2_U5365 = ~(P2_U2502 & P2_U2420); 
assign P2_U5369 = ~(P2_U5342 & P2_U2429); 
assign P2_U5370 = ~(P2_U2502 & P2_U2418); 
assign P2_U5374 = ~(P2_U5342 & P2_U2424); 
assign P2_U5375 = ~(P2_U2502 & P2_U2416); 
assign P2_U5379 = ~(P2_U5342 & P2_U2423); 
assign P2_U5380 = ~(P2_U2502 & P2_U2414); 
assign P2_U5384 = ~(P2_U5342 & P2_U2432); 
assign P2_U5385 = ~(P2_U2502 & P2_U2412); 
assign P2_U5389 = ~(P2_U5342 & P2_U2428); 
assign P2_U5390 = ~(P2_U2502 & P2_U2410); 
assign P2_U5394 = ~(P2_U5342 & P2_U2431); 
assign P2_U5395 = ~(P2_U2502 & P2_U2408); 
assign P2_U5416 = ~(P2_U5400 & P2_U2425); 
assign P2_U5417 = ~(P2_U2506 & P2_U2422); 
assign P2_U5421 = ~(P2_U5400 & P2_U2426); 
assign P2_U5422 = ~(P2_U2506 & P2_U2420); 
assign P2_U5426 = ~(P2_U5400 & P2_U2429); 
assign P2_U5427 = ~(P2_U2506 & P2_U2418); 
assign P2_U5431 = ~(P2_U5400 & P2_U2424); 
assign P2_U5432 = ~(P2_U2506 & P2_U2416); 
assign P2_U5436 = ~(P2_U5400 & P2_U2423); 
assign P2_U5437 = ~(P2_U2506 & P2_U2414); 
assign P2_U5441 = ~(P2_U5400 & P2_U2432); 
assign P2_U5442 = ~(P2_U2506 & P2_U2412); 
assign P2_U5446 = ~(P2_U5400 & P2_U2428); 
assign P2_U5447 = ~(P2_U2506 & P2_U2410); 
assign P2_U5451 = ~(P2_U5400 & P2_U2431); 
assign P2_U5452 = ~(P2_U2506 & P2_U2408); 
assign P2_U5474 = ~(P2_U5457 & P2_U2425); 
assign P2_U5475 = ~(P2_U2508 & P2_U2422); 
assign P2_U5479 = ~(P2_U5457 & P2_U2426); 
assign P2_U5480 = ~(P2_U2508 & P2_U2420); 
assign P2_U5484 = ~(P2_U5457 & P2_U2429); 
assign P2_U5485 = ~(P2_U2508 & P2_U2418); 
assign P2_U5489 = ~(P2_U5457 & P2_U2424); 
assign P2_U5490 = ~(P2_U2508 & P2_U2416); 
assign P2_U5494 = ~(P2_U5457 & P2_U2423); 
assign P2_U5495 = ~(P2_U2508 & P2_U2414); 
assign P2_U5499 = ~(P2_U5457 & P2_U2432); 
assign P2_U5500 = ~(P2_U2508 & P2_U2412); 
assign P2_U5504 = ~(P2_U5457 & P2_U2428); 
assign P2_U5505 = ~(P2_U2508 & P2_U2410); 
assign P2_U5509 = ~(P2_U5457 & P2_U2431); 
assign P2_U5510 = ~(P2_U2508 & P2_U2408); 
assign P2_U5531 = ~(P2_U5515 & P2_U2425); 
assign P2_U5532 = ~(P2_U2510 & P2_U2422); 
assign P2_U5536 = ~(P2_U5515 & P2_U2426); 
assign P2_U5537 = ~(P2_U2510 & P2_U2420); 
assign P2_U5541 = ~(P2_U5515 & P2_U2429); 
assign P2_U5542 = ~(P2_U2510 & P2_U2418); 
assign P2_U5546 = ~(P2_U5515 & P2_U2424); 
assign P2_U5547 = ~(P2_U2510 & P2_U2416); 
assign P2_U5551 = ~(P2_U5515 & P2_U2423); 
assign P2_U5552 = ~(P2_U2510 & P2_U2414); 
assign P2_U5556 = ~(P2_U5515 & P2_U2432); 
assign P2_U5557 = ~(P2_U2510 & P2_U2412); 
assign P2_U5561 = ~(P2_U5515 & P2_U2428); 
assign P2_U5562 = ~(P2_U2510 & P2_U2410); 
assign P2_U5566 = ~(P2_U5515 & P2_U2431); 
assign P2_U5567 = ~(P2_U2510 & P2_U2408); 
assign P2_U5584 = ~P2_U4394; 
assign P2_U5655 = ~(P2_U3892 & P2_U5652); 
assign P2_U6328 = ~(P2_ADD_391_1196_U87 & P2_U2397); 
assign P2_U6329 = ~(P2_U2380 & P2_R2096_U68); 
assign P2_U6332 = ~(P2_ADD_391_1196_U12 & P2_U2397); 
assign P2_U6333 = ~(P2_U2380 & P2_R2096_U51); 
assign P2_U6336 = ~(P2_ADD_391_1196_U92 & P2_U2397); 
assign P2_U6337 = ~(P2_U2380 & P2_R2096_U77); 
assign P2_U6340 = ~(P2_ADD_391_1196_U91 & P2_U2397); 
assign P2_U6341 = ~(P2_U2380 & P2_R2096_U75); 
assign P2_U6345 = ~(P2_U2380 & P2_R2096_U74); 
assign P2_U6349 = ~(P2_U2380 & P2_R2096_U73); 
assign P2_U6353 = ~(P2_U2380 & P2_R2096_U72); 
assign P2_U6357 = ~(P2_U2380 & P2_R2096_U71); 
assign P2_U6361 = ~(P2_U2380 & P2_R2096_U70); 
assign P2_U6365 = ~(P2_U2380 & P2_R2096_U69); 
assign P2_U6369 = ~(P2_U2380 & P2_R2096_U97); 
assign P2_U6373 = ~(P2_U2380 & P2_R2096_U96); 
assign P2_U6377 = ~(P2_U2380 & P2_R2096_U95); 
assign P2_U6381 = ~(P2_U2380 & P2_R2096_U94); 
assign P2_U6385 = ~(P2_U2380 & P2_R2096_U93); 
assign P2_U6471 = ~(P2_U2393 & P2_R2182_U69); 
assign P2_U6472 = ~(P2_U2379 & P2_R2099_U94); 
assign P2_U6474 = ~(P2_U2393 & P2_R2182_U68); 
assign P2_U6475 = ~(P2_U2379 & P2_R2099_U5); 
assign P2_U6477 = ~(P2_U2393 & P2_R2182_U40); 
assign P2_U6478 = ~(P2_U2379 & P2_R2099_U96); 
assign P2_U6480 = ~(P2_U2393 & P2_R2182_U76); 
assign P2_U6481 = ~(P2_U2379 & P2_R2099_U95); 
assign P2_U6483 = ~(P2_R2182_U75 & P2_U2393); 
assign P2_U6484 = ~(P2_U2379 & P2_R2099_U98); 
assign P2_U6486 = ~(P2_R2182_U74 & P2_U2393); 
assign P2_U6487 = ~(P2_U2379 & P2_R2099_U71); 
assign P2_U6489 = ~(P2_R2182_U73 & P2_U2393); 
assign P2_U6490 = ~(P2_U2379 & P2_R2099_U70); 
assign P2_U6492 = ~(P2_R2182_U72 & P2_U2393); 
assign P2_U6493 = ~(P2_U2379 & P2_R2099_U69); 
assign P2_U6496 = ~(P2_U2379 & P2_R2099_U68); 
assign P2_U6499 = ~(P2_U2379 & P2_R2099_U67); 
assign P2_U6576 = ~(P2_U2437 & P2_R2182_U69); 
assign P2_U6585 = ~(P2_U2437 & P2_R2182_U68); 
assign P2_U6594 = ~(P2_U2437 & P2_R2182_U40); 
assign P2_U6603 = ~(P2_U2437 & P2_R2182_U76); 
assign P2_U6612 = ~(P2_U2437 & P2_R2182_U75); 
assign P2_U6621 = ~(P2_U2437 & P2_R2182_U74); 
assign P2_U6838 = ~P2_U4400; 
assign P2_U6840 = ~(P2_U4400 & P2_FLUSH_REG_SCAN_IN); 
assign P2_U7894 = ~(P2_U4600 & P2_U4615); 
assign P2_U8072 = ~(P2_U3594 & P2_U4394); 
assign P2_U8084 = ~(P2_U5614 & P2_U4394); 
assign P2_U8134 = ~(P2_U4400 & P2_MORE_REG_SCAN_IN); 
assign P2_U8329 = ~(P2_R2256_U21 & P2_U3572); 
assign P2_U8393 = ~(P2_R2337_U79 & P2_U3284); 
assign P1_U2620 = P1_R2144_U145 & P1_U6746; 
assign P1_U2621 = P1_R2144_U145 & P1_U6746; 
assign P1_U2622 = P1_R2144_U145 & P1_U6746; 
assign P1_U2623 = P1_R2144_U145 & P1_U6746; 
assign P1_U2624 = P1_R2144_U145 & P1_U6746; 
assign P1_U2625 = P1_R2144_U145 & P1_U6746; 
assign P1_U2626 = P1_R2144_U145 & P1_U6746; 
assign P1_U2627 = P1_R2144_U145 & P1_U6746; 
assign P1_U2628 = P1_R2144_U145 & P1_U6746; 
assign P1_U2629 = P1_R2144_U145 & P1_U6746; 
assign P1_U2630 = P1_R2144_U145 & P1_U6746; 
assign P1_U2631 = P1_R2144_U145 & P1_U6746; 
assign P1_U2632 = P1_R2144_U145 & P1_U6746; 
assign P1_U2633 = P1_R2144_U145 & P1_U6746; 
assign P1_U2642 = P1_R2144_U80 & P1_U6746; 
assign P1_U2663 = ~(P1_U6825 & P1_U4022); 
assign P1_U2769 = P1_R2144_U145 & P1_U4159; 
assign P1_U2770 = P1_U4159 & P1_R2144_U145; 
assign P1_U2771 = P1_U4159 & P1_R2144_U145; 
assign P1_U2772 = P1_U4159 & P1_R2144_U145; 
assign P1_U2773 = P1_U4159 & P1_R2144_U145; 
assign P1_U2774 = P1_U4159 & P1_R2144_U145; 
assign P1_U2775 = P1_U4159 & P1_R2144_U145; 
assign P1_U2776 = P1_U4159 & P1_R2144_U145; 
assign P1_U2777 = P1_U4159 & P1_R2144_U145; 
assign P1_U2778 = P1_U4159 & P1_R2144_U145; 
assign P1_U2779 = P1_U4159 & P1_R2144_U145; 
assign P1_U2780 = P1_U4159 & P1_R2144_U145; 
assign P1_U2781 = P1_U4159 & P1_R2144_U145; 
assign P1_U2782 = P1_U4159 & P1_R2144_U145; 
assign P1_U2783 = P1_U4159 & P1_R2144_U145; 
assign P1_U2794 = ~(P1_U6876 & P1_U6875); 
assign P1_U3358 = ~(P1_U3342 & P1_U4530 & P1_U3357); 
assign P1_U3404 = ~(P1_U4242 & P1_U3300 & P1_U5536); 
assign P1_U4238 = ~P1_U3357; 
assign P1_U4245 = ~(P1_U2428 & P1_U3403); 
assign P1_U4511 = ~P1_U3293; 
assign P1_U4523 = ~(P1_U2368 & P1_U3293); 
assign P1_U4793 = ~(P1_U2491 & P1_U2413); 
assign P1_U4798 = ~(P1_U2491 & P1_U2411); 
assign P1_U4803 = ~(P1_U2491 & P1_U2409); 
assign P1_U4808 = ~(P1_U2491 & P1_U2407); 
assign P1_U4813 = ~(P1_U2491 & P1_U2405); 
assign P1_U4818 = ~(P1_U2491 & P1_U2403); 
assign P1_U4823 = ~(P1_U2491 & P1_U2401); 
assign P1_U4828 = ~(P1_U2491 & P1_U2399); 
assign P1_U4850 = ~(P1_U2493 & P1_U2413); 
assign P1_U4855 = ~(P1_U2493 & P1_U2411); 
assign P1_U4860 = ~(P1_U2493 & P1_U2409); 
assign P1_U4865 = ~(P1_U2493 & P1_U2407); 
assign P1_U4870 = ~(P1_U2493 & P1_U2405); 
assign P1_U4875 = ~(P1_U2493 & P1_U2403); 
assign P1_U4880 = ~(P1_U2493 & P1_U2401); 
assign P1_U4885 = ~(P1_U2493 & P1_U2399); 
assign P1_U4908 = ~(P1_U2495 & P1_U2413); 
assign P1_U4913 = ~(P1_U2495 & P1_U2411); 
assign P1_U4918 = ~(P1_U2495 & P1_U2409); 
assign P1_U4923 = ~(P1_U2495 & P1_U2407); 
assign P1_U4928 = ~(P1_U2495 & P1_U2405); 
assign P1_U4933 = ~(P1_U2495 & P1_U2403); 
assign P1_U4938 = ~(P1_U2495 & P1_U2401); 
assign P1_U4943 = ~(P1_U2495 & P1_U2399); 
assign P1_U4965 = ~(P1_U2497 & P1_U2413); 
assign P1_U4970 = ~(P1_U2497 & P1_U2411); 
assign P1_U4975 = ~(P1_U2497 & P1_U2409); 
assign P1_U4980 = ~(P1_U2497 & P1_U2407); 
assign P1_U4985 = ~(P1_U2497 & P1_U2405); 
assign P1_U4990 = ~(P1_U2497 & P1_U2403); 
assign P1_U4995 = ~(P1_U2497 & P1_U2401); 
assign P1_U5000 = ~(P1_U2497 & P1_U2399); 
assign P1_U5078 = ~(P1_U2501 & P1_U2413); 
assign P1_U5083 = ~(P1_U2501 & P1_U2411); 
assign P1_U5088 = ~(P1_U2501 & P1_U2409); 
assign P1_U5093 = ~(P1_U2501 & P1_U2407); 
assign P1_U5098 = ~(P1_U2501 & P1_U2405); 
assign P1_U5103 = ~(P1_U2501 & P1_U2403); 
assign P1_U5108 = ~(P1_U2501 & P1_U2401); 
assign P1_U5113 = ~(P1_U2501 & P1_U2399); 
assign P1_U5136 = ~(P1_U2503 & P1_U2413); 
assign P1_U5141 = ~(P1_U2503 & P1_U2411); 
assign P1_U5146 = ~(P1_U2503 & P1_U2409); 
assign P1_U5151 = ~(P1_U2503 & P1_U2407); 
assign P1_U5156 = ~(P1_U2503 & P1_U2405); 
assign P1_U5161 = ~(P1_U2503 & P1_U2403); 
assign P1_U5166 = ~(P1_U2503 & P1_U2401); 
assign P1_U5171 = ~(P1_U2503 & P1_U2399); 
assign P1_U5193 = ~(P1_U2505 & P1_U2413); 
assign P1_U5198 = ~(P1_U2505 & P1_U2411); 
assign P1_U5203 = ~(P1_U2505 & P1_U2409); 
assign P1_U5208 = ~(P1_U2505 & P1_U2407); 
assign P1_U5213 = ~(P1_U2505 & P1_U2405); 
assign P1_U5218 = ~(P1_U2505 & P1_U2403); 
assign P1_U5223 = ~(P1_U2505 & P1_U2401); 
assign P1_U5228 = ~(P1_U2505 & P1_U2399); 
assign P1_U5551 = ~(P1_U2388 & P1_U5550); 
assign P1_U5703 = ~(P1_R2099_U76 & P1_U2380); 
assign P1_U5713 = ~(P1_ADD_405_U68 & P1_U2375); 
assign P1_U5714 = ~(P1_ADD_515_U68 & P1_U2374); 
assign P1_U5802 = ~(P1_R2358_U76 & P1_U2364); 
assign P1_U5899 = ~(P1_R2337_U81 & P1_U2376); 
assign P1_U6155 = ~(P1_U2386 & P1_R2358_U76); 
assign P1_U6265 = ~(P1_U2383 & P1_R2358_U76); 
assign P1_U6323 = ~(P1_U2371 & P1_R2099_U76); 
assign P1_U6507 = ~(P1_U2604 & P1_R2099_U76); 
assign P1_U6515 = ~(P1_R2096_U81 & P1_U7485); 
assign P1_U6819 = ~(P1_R2337_U81 & P1_U2352); 
assign P1_U6871 = ~(P1_U4159 & P1_R2144_U80); 
assign P1_U7731 = ~(P1_U7693 & P1_U4527); 
assign P3_ADD_476_U44 = ~(P3_ADD_476_U112 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_476_U160 = ~(P3_ADD_476_U112 & P3_ADD_476_U43); 
assign P3_ADD_531_U45 = ~(P3_ADD_531_U116 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_531_U167 = ~(P3_ADD_531_U116 & P3_ADD_531_U44); 
assign P3_SUB_320_U44 = ~P3_ADD_318_U81; 
assign P3_SUB_320_U74 = P3_SUB_320_U151 & P3_SUB_320_U150; 
assign P3_SUB_320_U116 = ~(P3_ADD_318_U81 & P3_SUB_320_U115); 
assign P3_ADD_318_U44 = ~(P3_ADD_318_U112 & P3_PHYADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_318_U160 = ~(P3_ADD_318_U112 & P3_ADD_318_U43); 
assign P3_ADD_315_U44 = ~(P3_ADD_315_U109 & P3_PHYADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_315_U152 = ~(P3_ADD_315_U109 & P3_ADD_315_U43); 
assign P3_ADD_360_1242_U81 = ~(P3_ADD_360_1242_U250 & P3_ADD_360_1242_U249); 
assign P3_ADD_360_1242_U158 = ~P3_ADD_360_1242_U56; 
assign P3_ADD_360_1242_U175 = ~(P3_ADD_360_1242_U57 & P3_ADD_360_1242_U56); 
assign P3_ADD_360_1242_U177 = ~(P3_ADD_360_1242_U55 & P3_ADD_360_1242_U176); 
assign P3_ADD_467_U44 = ~(P3_ADD_467_U112 & P3_REIP_REG_21__SCAN_IN); 
assign P3_ADD_467_U160 = ~(P3_ADD_467_U112 & P3_ADD_467_U43); 
assign P3_ADD_430_U44 = ~(P3_ADD_430_U112 & P3_REIP_REG_21__SCAN_IN); 
assign P3_ADD_430_U160 = ~(P3_ADD_430_U112 & P3_ADD_430_U43); 
assign P3_ADD_380_U45 = ~(P3_ADD_380_U116 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_380_U167 = ~(P3_ADD_380_U116 & P3_ADD_380_U44); 
assign P3_ADD_344_U45 = ~(P3_ADD_344_U116 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_344_U167 = ~(P3_ADD_344_U116 & P3_ADD_344_U44); 
assign P3_ADD_339_U44 = ~(P3_ADD_339_U112 & P3_PHYADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_339_U160 = ~(P3_ADD_339_U112 & P3_ADD_339_U43); 
assign P3_ADD_541_U44 = ~(P3_ADD_541_U112 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_541_U160 = ~(P3_ADD_541_U112 & P3_ADD_541_U43); 
assign P3_SUB_357_1258_U16 = P3_SUB_357_1258_U249 & P3_SUB_357_1258_U248; 
assign P3_SUB_357_1258_U87 = ~(P3_SUB_357_1258_U438 & P3_SUB_357_1258_U437); 
assign P3_SUB_357_1258_U218 = ~(P3_SUB_357_1258_U63 & P3_SUB_357_1258_U153); 
assign P3_SUB_357_1258_U229 = ~(P3_SUB_357_1258_U228 & P3_SUB_357_1258_U63); 
assign P3_SUB_357_1258_U237 = ~(P3_SUB_357_1258_U207 & P3_SUB_357_1258_U64); 
assign P3_SUB_357_1258_U240 = ~(P3_SUB_357_1258_U64 & P3_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P3_SUB_357_1258_U277 = ~P3_SUB_357_1258_U64; 
assign P3_SUB_357_1258_U279 = ~P3_SUB_357_1258_U137; 
assign P3_SUB_357_1258_U281 = ~P3_SUB_357_1258_U135; 
assign P3_SUB_357_1258_U283 = ~P3_SUB_357_1258_U133; 
assign P3_SUB_357_1258_U285 = ~P3_SUB_357_1258_U63; 
assign P3_SUB_357_1258_U390 = ~(P3_SUB_357_1258_U63 & P3_SUB_357_1258_U262); 
assign P3_SUB_357_1258_U397 = ~(P3_SUB_357_1258_U132 & P3_SUB_357_1258_U133); 
assign P3_SUB_357_1258_U404 = ~(P3_SUB_357_1258_U134 & P3_SUB_357_1258_U135); 
assign P3_SUB_357_1258_U411 = ~(P3_SUB_357_1258_U136 & P3_SUB_357_1258_U137); 
assign P3_SUB_357_1258_U430 = ~(P3_SUB_357_1258_U64 & P3_SUB_357_1258_U263); 
assign P3_ADD_515_U44 = ~(P3_ADD_515_U112 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_515_U160 = ~(P3_ADD_515_U112 & P3_ADD_515_U43); 
assign P3_ADD_394_U44 = ~(P3_ADD_394_U115 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_394_U162 = ~(P3_ADD_394_U115 & P3_ADD_394_U43); 
assign P3_ADD_441_U44 = ~(P3_ADD_441_U112 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_441_U160 = ~(P3_ADD_441_U112 & P3_ADD_441_U43); 
assign P3_ADD_349_U45 = ~(P3_ADD_349_U116 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_349_U167 = ~(P3_ADD_349_U116 & P3_ADD_349_U44); 
assign P3_ADD_405_U44 = ~(P3_ADD_405_U115 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_405_U162 = ~(P3_ADD_405_U115 & P3_ADD_405_U43); 
assign P3_ADD_553_U45 = ~(P3_ADD_553_U116 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_553_U167 = ~(P3_ADD_553_U116 & P3_ADD_553_U44); 
assign P3_ADD_558_U45 = ~(P3_ADD_558_U116 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_558_U167 = ~(P3_ADD_558_U116 & P3_ADD_558_U44); 
assign P3_ADD_385_U45 = ~(P3_ADD_385_U116 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_385_U167 = ~(P3_ADD_385_U116 & P3_ADD_385_U44); 
assign P3_ADD_547_U45 = ~(P3_ADD_547_U116 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_547_U167 = ~(P3_ADD_547_U116 & P3_ADD_547_U44); 
assign P3_ADD_371_1212_U8 = P3_ADD_371_1212_U191 & P3_ADD_371_1212_U53; 
assign P3_ADD_371_1212_U9 = P3_ADD_371_1212_U189 & P3_ADD_371_1212_U56; 
assign P3_ADD_371_1212_U59 = ~(P3_ADD_371_1212_U103 & P3_ADD_371_1212_U166); 
assign P3_ADD_371_1212_U186 = ~(P3_ADD_371_1212_U166 & P3_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P3_ADD_371_1212_U257 = ~(P3_ADD_371_1212_U166 & P3_ADD_371_1212_U57); 
assign P3_ADD_494_U44 = ~(P3_ADD_494_U112 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_494_U160 = ~(P3_ADD_494_U112 & P3_ADD_494_U43); 
assign P3_ADD_536_U44 = ~(P3_ADD_536_U112 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_536_U160 = ~(P3_ADD_536_U112 & P3_ADD_536_U43); 
assign P2_R2099_U93 = ~(P2_R2099_U223 & P2_R2099_U222); 
assign P2_R2099_U126 = ~P2_R2099_U27; 
assign P2_R2099_U220 = ~(P2_U2736 & P2_R2099_U27); 
assign P2_ADD_391_1196_U13 = ~P2_R2182_U72; 
assign P2_ADD_391_1196_U39 = ~(P2_ADD_391_1196_U38 & P2_ADD_391_1196_U178); 
assign P2_ADD_391_1196_U43 = ~P2_R2096_U93; 
assign P2_ADD_391_1196_U90 = ~(P2_ADD_391_1196_U331 & P2_ADD_391_1196_U330); 
assign P2_ADD_391_1196_U114 = P2_ADD_391_1196_U324 & P2_ADD_391_1196_U323; 
assign P2_ADD_391_1196_U177 = ~P2_ADD_391_1196_U38; 
assign P2_ADD_391_1196_U183 = P2_R2096_U71 | P2_R2182_U72; 
assign P2_ADD_391_1196_U186 = ~(P2_R2096_U71 & P2_R2182_U72); 
assign P2_ADD_391_1196_U200 = ~(P2_R2096_U71 & P2_R2182_U72); 
assign P2_ADD_391_1196_U303 = ~(P2_ADD_391_1196_U202 & P2_ADD_391_1196_U161); 
assign P2_ADD_391_1196_U317 = ~(P2_R2182_U72 & P2_ADD_391_1196_U14); 
assign P2_ADD_391_1196_U318 = ~(P2_R2096_U72 & P2_ADD_391_1196_U15); 
assign P2_R2182_U4 = P2_U2671 & P2_R2182_U20; 
assign P2_R2182_U71 = ~(P2_R2182_U196 & P2_R2182_U195); 
assign P2_R2182_U141 = ~P2_R2182_U20; 
assign P2_R2182_U194 = ~(P2_R2182_U140 & P2_U2672); 
assign P2_R2182_U302 = ~(P2_R2182_U23 & P2_R2182_U20); 
assign P2_R2027_U45 = ~(P2_R2027_U116 & P2_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P2_R2027_U167 = ~(P2_R2027_U116 & P2_R2027_U44); 
assign P2_R2337_U45 = ~(P2_R2337_U113 & P2_PHYADDRPOINTER_REG_22__SCAN_IN); 
assign P2_R2337_U158 = ~(P2_R2337_U113 & P2_R2337_U44); 
assign P2_R2096_U25 = P2_U2632 & P2_R2096_U5; 
assign P2_R2096_U92 = ~(P2_R2096_U253 & P2_R2096_U252); 
assign P2_R2096_U152 = ~P2_R2096_U5; 
assign P2_R2096_U248 = ~(P2_R2096_U48 & P2_R2096_U5); 
assign P2_R2096_U251 = ~(P2_R2096_U151 & P2_U2633); 
assign P2_R2256_U28 = ~(P2_R2256_U30 & P2_R2256_U35); 
assign P2_R2256_U31 = P2_R2256_U68 & P2_R2256_U67; 
assign P2_R2256_U66 = ~(P2_R2256_U65 & P2_R2256_U64); 
assign P2_R1957_U43 = ~P2_U3670; 
assign P2_R1957_U74 = P2_R1957_U151 & P2_R1957_U150; 
assign P2_R1957_U116 = ~(P2_U3670 & P2_R1957_U115); 
assign P2_R2278_U47 = ~P2_U2810; 
assign P2_R2278_U145 = P2_R2278_U347 & P2_R2278_U346; 
assign P2_R2278_U240 = ~P2_R2278_U52; 
assign P2_R2278_U242 = P2_U2810 | P2_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P2_R2278_U243 = ~(P2_U2810 & P2_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P2_R2278_U350 = ~(P2_R2278_U349 & P2_R2278_U348); 
assign P2_R2278_U548 = ~(P2_U2810 & P2_R2278_U48); 
assign P2_R2278_U550 = ~(P2_U2810 & P2_R2278_U48); 
assign P2_R2278_U554 = ~(P2_R2278_U50 & P2_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P2_R2278_U556 = ~(P2_R2278_U50 & P2_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P2_ADD_394_U44 = ~(P2_ADD_394_U115 & P2_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P2_ADD_394_U178 = ~(P2_ADD_394_U115 & P2_ADD_394_U43); 
assign P2_R2267_U7 = P2_R2267_U131 & P2_R2267_U32; 
assign P2_R2267_U33 = ~(P2_R2267_U47 & P2_R2267_U103); 
assign P2_R2267_U128 = ~(P2_R2267_U103 & P2_R2267_U82); 
assign P2_R2267_U162 = ~(P2_R2267_U103 & P2_R2267_U82); 
assign P2_ADD_371_1212_U27 = ~P2_R2256_U21; 
assign P2_ADD_371_1212_U29 = ~(P2_R2256_U21 & P2_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P2_ADD_371_1212_U206 = ~(P2_R2256_U21 & P2_ADD_371_1212_U26); 
assign P1_R2144_U11 = ~(P1_R2144_U144 & P1_R2144_U146); 
assign P1_R2144_U30 = ~(P1_R2144_U209 & P1_R2144_U208); 
assign P1_R2144_U40 = ~(P1_R2144_U254 & P1_R2144_U253); 
assign P1_R2144_U41 = ~(P1_R2144_U256 & P1_R2144_U255); 
assign P1_R2144_U42 = ~(P1_R2144_U258 & P1_R2144_U257); 
assign P1_R2144_U142 = ~P1_R2144_U95; 
assign P1_R2144_U143 = ~P1_R2144_U26; 
assign P1_R2144_U250 = ~(P1_R2144_U32 & P1_R2144_U26); 
assign P1_R2144_U252 = ~(P1_R2144_U33 & P1_R2144_U95); 
assign P1_R2278_U19 = ~(P1_R2278_U214 & P1_R2278_U429); 
assign P1_R2278_U24 = ~P1_U2793; 
assign P1_R2278_U28 = ~P1_U2795; 
assign P1_R2278_U39 = ~P1_U2796; 
assign P1_R2278_U127 = P1_U2793 & P1_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P1_R2278_U191 = P1_R2278_U479 & P1_R2278_U478; 
assign P1_R2278_U235 = ~P1_R2278_U192; 
assign P1_R2278_U237 = ~(P1_R2278_U236 & P1_R2278_U192); 
assign P1_R2278_U244 = P1_U2796 | P1_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P1_R2278_U246 = ~(P1_U2796 & P1_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P1_R2278_U248 = P1_U2795 | P1_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P1_R2278_U250 = ~(P1_U2795 & P1_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P1_R2278_U253 = P1_U2793 | P1_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P1_R2278_U256 = ~(P1_U2793 & P1_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P1_R2278_U267 = ~(P1_U2793 & P1_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P1_R2278_U271 = ~(P1_U2795 & P1_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P1_R2278_U439 = ~(P1_U2793 & P1_R2278_U23); 
assign P1_R2278_U446 = ~(P1_U2795 & P1_R2278_U27); 
assign P1_R2278_U448 = ~(P1_U2796 & P1_R2278_U38); 
assign P1_R2278_U450 = ~(P1_U2796 & P1_R2278_U38); 
assign P1_R2278_U456 = ~(P1_R2278_U37 & P1_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P1_R2278_U458 = ~(P1_R2278_U37 & P1_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P1_R2278_U482 = ~(P1_R2278_U481 & P1_R2278_U480); 
assign P1_R2358_U25 = ~P1_U2644; 
assign P1_R2358_U66 = ~(P1_R2358_U65 & P1_R2358_U202); 
assign P1_R2358_U107 = ~(P1_R2358_U597 & P1_R2358_U596); 
assign P1_R2358_U121 = P1_R2358_U204 & P1_R2358_U202; 
assign P1_R2358_U123 = P1_R2358_U204 & P1_R2358_U203; 
assign P1_R2358_U215 = ~(P1_U2644 & P1_R2358_U408); 
assign P1_R2358_U217 = ~(P1_R2358_U405 & P1_R2358_U404 & P1_R2358_U24); 
assign P1_R2358_U219 = ~(P1_R2358_U410 & P1_R2358_U409 & P1_R2358_U26); 
assign P1_R2358_U221 = ~P1_R2358_U28; 
assign P1_R2358_U225 = ~(P1_R2358_U443 & P1_R2358_U442 & P1_R2358_U27); 
assign P1_R2358_U249 = ~P1_R2358_U65; 
assign P1_R2358_U253 = ~(P1_R2358_U204 & P1_R2358_U203); 
assign P1_R2358_U306 = ~(P1_R2358_U207 & P1_R2358_U202); 
assign P1_R2358_U491 = ~(P1_U2352 & P1_R2358_U165); 
assign P1_R2358_U493 = ~(P1_U2352 & P1_R2358_U165); 
assign P1_R2099_U17 = ~(P1_R2099_U171 & P1_R2099_U53); 
assign P1_R2099_U316 = ~(P1_R2099_U252 & P1_R2099_U171); 
assign P1_R2337_U44 = ~(P1_R2337_U112 & P1_PHYADDRPOINTER_REG_21__SCAN_IN); 
assign P1_R2337_U160 = ~(P1_R2337_U112 & P1_R2337_U43); 
assign P1_R2096_U44 = ~(P1_R2096_U112 & P1_REIP_REG_21__SCAN_IN); 
assign P1_R2096_U160 = ~(P1_R2096_U112 & P1_R2096_U43); 
assign P1_ADD_405_U44 = ~(P1_ADD_405_U115 & P1_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P1_ADD_405_U178 = ~(P1_ADD_405_U115 & P1_ADD_405_U43); 
assign P1_ADD_515_U44 = ~(P1_ADD_515_U112 & P1_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P1_ADD_515_U174 = ~(P1_ADD_515_U112 & P1_ADD_515_U43); 
assign P3_U2850 = ~(P3_U5943 & P3_U5941 & P3_U5942); 
assign P3_U3802 = P3_U3801 & P3_U3800 & P3_U5987; 
assign P3_U3807 = P3_U3804 & P3_U5994 & P3_U3806 & P3_U5993 & P3_U5992; 
assign P3_U3818 = P3_U3817 & P3_U3816 & P3_U6035; 
assign P3_U3832 = P3_U6092 & P3_U6091; 
assign P3_U3836 = P3_U6106 & P3_U6105 & P3_U6104 & P3_U6103; 
assign P3_U3839 = P3_U6121 & P3_U6120; 
assign P3_U3842 = P3_U6123 & P3_U6122 & P3_U6124 & P3_U6126 & P3_U6125; 
assign P3_U3968 = P3_U6524 & P3_U6521 & P3_U6522 & P3_U6523; 
assign P3_U3970 = P3_U6540 & P3_U6537 & P3_U6538 & P3_U6539; 
assign P3_U4099 = P3_U7270 & P3_U7269; 
assign P3_U5966 = ~(P3_U4318 & P3_U5964); 
assign P3_U6011 = ~(P3_ADD_371_1212_U8 & P3_U2360); 
assign P3_U6041 = ~(P3_SUB_357_1258_U16 & P3_U2393); 
assign P3_U6059 = ~(P3_ADD_371_1212_U9 & P3_U2360); 
assign P3_U6064 = ~(P3_ADD_360_1242_U81 & P3_U2395); 
assign P3_U6065 = ~(P3_SUB_357_1258_U87 & P3_U2393); 
assign P3_U6531 = ~(P3_U2387 & P3_ADD_371_1212_U8); 
assign P3_U6544 = ~(P3_U2394 & P3_SUB_357_1258_U16); 
assign P3_U6547 = ~(P3_U2387 & P3_ADD_371_1212_U9); 
assign P3_U6551 = ~(P3_U2396 & P3_ADD_360_1242_U81); 
assign P3_U6552 = ~(P3_U2394 & P3_SUB_357_1258_U87); 
assign P3_U7952 = ~(P3_U4627 & P3_STATE2_REG_0__SCAN_IN); 
assign P2_U2468 = P2_U3320 & P2_U4657; 
assign P2_U2471 = P2_U3339 & P2_U4715; 
assign P2_U2474 = P2_U3354 & P2_U4774; 
assign P2_U2480 = P2_U3366 & P2_U4831; 
assign P2_U2484 = P2_U3379 & P2_U4889; 
assign P2_U2486 = P2_U3391 & P2_U4946; 
assign P2_U2488 = P2_U3402 & P2_U5004; 
assign P2_U2490 = P2_U3414 & P2_U5061; 
assign P2_U2587 = P2_U2391 & P2_EBX_REG_31__SCAN_IN; 
assign P2_U2588 = P2_U2377 & P2_U2360; 
assign P2_U2808 = P2_U3242 & P2_R2267_U7; 
assign P2_U2880 = ~(P2_U6493 & P2_U6492 & P2_U6494); 
assign P2_U2881 = ~(P2_U6490 & P2_U6489 & P2_U6491); 
assign P2_U2882 = ~(P2_U6487 & P2_U6486 & P2_U6488); 
assign P2_U2883 = ~(P2_U6484 & P2_U6483 & P2_U6485); 
assign P2_U2884 = ~(P2_U6481 & P2_U6480 & P2_U6482); 
assign P2_U2885 = ~(P2_U6478 & P2_U6477 & P2_U6479); 
assign P2_U2886 = ~(P2_U6475 & P2_U6474 & P2_U6476); 
assign P2_U2887 = ~(P2_U6472 & P2_U6471 & P2_U6473); 
assign P2_U3427 = ~(P2_U2491 & P2_U4636); 
assign P2_U3440 = ~(P2_U2491 & P2_U4709); 
assign P2_U3451 = ~(P2_U2491 & P2_U4767); 
assign P2_U3463 = ~(P2_U2491 & P2_U2475); 
assign P2_U3474 = ~(P2_U2500 & P2_U4636); 
assign P2_U3486 = ~(P2_U2500 & P2_U4709); 
assign P2_U3497 = ~(P2_U2500 & P2_U4767); 
assign P2_U3509 = ~(P2_U2500 & P2_U2475); 
assign P2_U3638 = ~(P2_U8330 & P2_U8329); 
assign P2_U3669 = ~(P2_U8394 & P2_U8393); 
assign P2_U4059 = P2_U6330 & P2_U6329; 
assign P2_U4060 = P2_U6334 & P2_U6333; 
assign P2_U4061 = P2_U6338 & P2_U6337; 
assign P2_U4062 = P2_U6342 & P2_U6341; 
assign P2_U4063 = P2_U6346 & P2_U6345; 
assign P2_U4064 = P2_U6350 & P2_U6349; 
assign P2_U4065 = P2_U6354 & P2_U6353; 
assign P2_U4066 = P2_U6358 & P2_U6357; 
assign P2_U4067 = P2_U6362 & P2_U6361; 
assign P2_U4068 = P2_U6366 & P2_U6365; 
assign P2_U4641 = ~P2_U3320; 
assign P2_U4710 = ~P2_U3339; 
assign P2_U4768 = ~P2_U3354; 
assign P2_U4826 = ~P2_U3366; 
assign P2_U4883 = ~P2_U3379; 
assign P2_U4941 = ~P2_U3391; 
assign P2_U4998 = ~P2_U3402; 
assign P2_U5056 = ~P2_U3414; 
assign P2_U6327 = ~(P2_U2433 & U314); 
assign P2_U6331 = ~(P2_U2433 & U303); 
assign P2_U6335 = ~(P2_U2433 & U292); 
assign P2_U6339 = ~(P2_U2433 & U289); 
assign P2_U6343 = ~(P2_U2433 & U288); 
assign P2_U6344 = ~(P2_ADD_391_1196_U90 & P2_U2397); 
assign P2_U6347 = ~(P2_U2433 & U287); 
assign P2_U6351 = ~(P2_U2433 & U286); 
assign P2_U6355 = ~(P2_U2433 & U285); 
assign P2_U6359 = ~(P2_U2433 & U284); 
assign P2_U6363 = ~(P2_U2433 & U283); 
assign P2_U6367 = ~(P2_U2433 & U313); 
assign P2_U6371 = ~(P2_U2433 & U312); 
assign P2_U6375 = ~(P2_U2433 & U311); 
assign P2_U6379 = ~(P2_U2433 & U310); 
assign P2_U6383 = ~(P2_U2433 & U309); 
assign P2_U6387 = ~(P2_U2433 & U308); 
assign P2_U6389 = ~(P2_U2380 & P2_R2096_U92); 
assign P2_U6391 = ~(P2_U2434 & U314); 
assign P2_U6392 = ~(P2_U2427 & U307); 
assign P2_U6396 = ~(P2_U2434 & U303); 
assign P2_U6397 = ~(P2_U2427 & U306); 
assign P2_U6401 = ~(P2_U2434 & U292); 
assign P2_U6402 = ~(P2_U2427 & U305); 
assign P2_U6406 = ~(P2_U2434 & U289); 
assign P2_U6407 = ~(P2_U2427 & U304); 
assign P2_U6411 = ~(P2_U2434 & U288); 
assign P2_U6412 = ~(P2_U2427 & U302); 
assign P2_U6416 = ~(P2_U2434 & U287); 
assign P2_U6417 = ~(P2_U2427 & U301); 
assign P2_U6421 = ~(P2_U2434 & U286); 
assign P2_U6422 = ~(P2_U2427 & U300); 
assign P2_U6426 = ~(P2_U2434 & U285); 
assign P2_U6427 = ~(P2_U2427 & U299); 
assign P2_U6431 = ~(P2_U2434 & U284); 
assign P2_U6432 = ~(P2_U2427 & U298); 
assign P2_U6436 = ~(P2_U2434 & U283); 
assign P2_U6437 = ~(P2_U2427 & U297); 
assign P2_U6441 = ~(P2_U2434 & U313); 
assign P2_U6442 = ~(P2_U2427 & U296); 
assign P2_U6446 = ~(P2_U2434 & U312); 
assign P2_U6447 = ~(P2_U2427 & U295); 
assign P2_U6451 = ~(P2_U2434 & U311); 
assign P2_U6452 = ~(P2_U2427 & U294); 
assign P2_U6456 = ~(P2_U2434 & U310); 
assign P2_U6457 = ~(P2_U2427 & U293); 
assign P2_U6461 = ~(P2_U2434 & U309); 
assign P2_U6462 = ~(P2_U2427 & U291); 
assign P2_U6466 = ~(P2_U2427 & U290); 
assign P2_U6495 = ~(P2_R2182_U71 & P2_U2393); 
assign P2_U6502 = ~(P2_U2379 & P2_R2099_U93); 
assign P2_U6577 = ~(P2_U2392 & P2_R2099_U94); 
assign P2_U6586 = ~(P2_U2392 & P2_R2099_U5); 
assign P2_U6595 = ~(P2_U2392 & P2_R2099_U96); 
assign P2_U6604 = ~(P2_U2392 & P2_R2099_U95); 
assign P2_U6613 = ~(P2_U2392 & P2_R2099_U98); 
assign P2_U6622 = ~(P2_U2392 & P2_R2099_U71); 
assign P2_U6630 = ~(P2_U2392 & P2_R2099_U70); 
assign P2_U6638 = ~(P2_U2392 & P2_R2099_U69); 
assign P2_U6646 = ~(P2_U2392 & P2_R2099_U68); 
assign P2_U6654 = ~(P2_U2392 & P2_R2099_U67); 
assign P2_U6662 = ~(P2_U2392 & P2_R2099_U93); 
assign P2_U7741 = ~(P2_U2391 & P2_U3544); 
assign P2_U7742 = ~(P2_U2377 & P2_U6572); 
assign P2_U8073 = ~(P2_U5584 & P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign P2_U8083 = ~(P2_U5584 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign P2_U8093 = ~(P2_U5584 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign P2_U8101 = ~(P2_U5584 & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign P2_U8103 = ~(P2_U5584 & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign P1_U2475 = P1_U3454 & P1_U3358; 
assign P1_U2490 = P1_U7693 & P1_U3358; 
assign P1_U2634 = P1_R2144_U11 & P1_U6746; 
assign P1_U2638 = P1_R2144_U40 & P1_U6746; 
assign P1_U2639 = P1_R2144_U41 & P1_U6746; 
assign P1_U2640 = P1_R2144_U42 & P1_U6746; 
assign P1_U2641 = P1_R2144_U30 & P1_U6746; 
assign P1_U2784 = P1_U4159 & P1_R2144_U11; 
assign P1_U2788 = P1_U4159 & P1_R2144_U40; 
assign P1_U2789 = P1_U4159 & P1_R2144_U41; 
assign P1_U2790 = P1_U4159 & P1_R2144_U42; 
assign P1_U2791 = P1_U4159 & P1_R2144_U30; 
assign P1_U2792 = ~(P1_U6872 & P1_U6871); 
assign P1_U2872 = ~(P1_U6266 & P1_U6265 & P1_U6267); 
assign P1_U2904 = ~(P1_U6155 & P1_U6154 & P1_U6156); 
assign P1_U2999 = ~(P1_U5800 & P1_U5799 & P1_U5801 & P1_U5803 & P1_U5802); 
assign P1_U3586 = P1_U3585 & P1_U4523; 
assign P1_U3826 = P1_U5711 & P1_U5713; 
assign P1_U3828 = P1_U3827 & P1_U5714; 
assign P1_U3926 = P1_U6517 & P1_U6515; 
assign P1_U4020 = P1_U6817 & P1_U6818 & P1_U6819; 
assign P1_U4512 = ~(P1_U4511 & P1_U3262); 
assign P1_U4531 = ~P1_U3358; 
assign P1_U5021 = ~(P1_U4238 & P1_U2413); 
assign P1_U5026 = ~(P1_U4238 & P1_U2411); 
assign P1_U5031 = ~(P1_U4238 & P1_U2409); 
assign P1_U5036 = ~(P1_U4238 & P1_U2407); 
assign P1_U5041 = ~(P1_U4238 & P1_U2405); 
assign P1_U5046 = ~(P1_U4238 & P1_U2403); 
assign P1_U5051 = ~(P1_U4238 & P1_U2401); 
assign P1_U5056 = ~(P1_U4238 & P1_U2399); 
assign P1_U5537 = ~P1_U3404; 
assign P1_U5540 = ~(P1_U3358 & P1_U5539); 
assign P1_U5554 = ~(P1_U3753 & P1_U5551); 
assign P1_U5557 = ~(P1_U5555 & P1_U5556 & P1_U4245); 
assign P1_U5579 = ~(P1_R2278_U19 & P1_U2377); 
assign P1_U5805 = ~(P1_U2372 & P1_R2278_U19); 
assign P1_U5807 = ~(P1_R2358_U107 & P1_U2364); 
assign P1_U6158 = ~(P1_U2386 & P1_R2358_U107); 
assign P1_U6268 = ~(P1_U2383 & P1_R2358_U107); 
assign P1_U7733 = ~(P1_U7732 & P1_U7731); 
assign P3_ADD_476_U80 = ~(P3_ADD_476_U160 & P3_ADD_476_U159); 
assign P3_ADD_476_U113 = ~P3_ADD_476_U44; 
assign P3_ADD_476_U157 = ~(P3_ADD_476_U44 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_531_U84 = ~(P3_ADD_531_U167 & P3_ADD_531_U166); 
assign P3_ADD_531_U117 = ~P3_ADD_531_U45; 
assign P3_ADD_531_U164 = ~(P3_ADD_531_U45 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_SUB_320_U33 = ~(P3_SUB_320_U44 & P3_SUB_320_U73 & P3_SUB_320_U97); 
assign P3_ADD_318_U80 = ~(P3_ADD_318_U160 & P3_ADD_318_U159); 
assign P3_ADD_318_U113 = ~P3_ADD_318_U44; 
assign P3_ADD_318_U157 = ~(P3_ADD_318_U44 & P3_PHYADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_315_U76 = ~(P3_ADD_315_U152 & P3_ADD_315_U151); 
assign P3_ADD_315_U110 = ~P3_ADD_315_U44; 
assign P3_ADD_315_U149 = ~(P3_ADD_315_U44 & P3_PHYADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_360_1242_U9 = P3_ADD_360_1242_U177 & P3_ADD_360_1242_U56; 
assign P3_ADD_360_1242_U58 = ~(P3_ADD_360_1242_U158 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_467_U80 = ~(P3_ADD_467_U160 & P3_ADD_467_U159); 
assign P3_ADD_467_U113 = ~P3_ADD_467_U44; 
assign P3_ADD_467_U157 = ~(P3_ADD_467_U44 & P3_REIP_REG_22__SCAN_IN); 
assign P3_ADD_430_U80 = ~(P3_ADD_430_U160 & P3_ADD_430_U159); 
assign P3_ADD_430_U113 = ~P3_ADD_430_U44; 
assign P3_ADD_430_U157 = ~(P3_ADD_430_U44 & P3_REIP_REG_22__SCAN_IN); 
assign P3_ADD_380_U84 = ~(P3_ADD_380_U167 & P3_ADD_380_U166); 
assign P3_ADD_380_U117 = ~P3_ADD_380_U45; 
assign P3_ADD_380_U164 = ~(P3_ADD_380_U45 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_344_U84 = ~(P3_ADD_344_U167 & P3_ADD_344_U166); 
assign P3_ADD_344_U117 = ~P3_ADD_344_U45; 
assign P3_ADD_344_U164 = ~(P3_ADD_344_U45 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_339_U80 = ~(P3_ADD_339_U160 & P3_ADD_339_U159); 
assign P3_ADD_339_U113 = ~P3_ADD_339_U44; 
assign P3_ADD_339_U157 = ~(P3_ADD_339_U44 & P3_PHYADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_541_U80 = ~(P3_ADD_541_U160 & P3_ADD_541_U159); 
assign P3_ADD_541_U113 = ~P3_ADD_541_U44; 
assign P3_ADD_541_U157 = ~(P3_ADD_541_U44 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_SUB_357_1258_U62 = ~(P3_SUB_357_1258_U105 & P3_SUB_357_1258_U218); 
assign P3_SUB_357_1258_U65 = ~(P3_SUB_357_1258_U277 & P3_SUB_357_1258_U47); 
assign P3_SUB_357_1258_U111 = P3_SUB_357_1258_U237 & P3_SUB_357_1258_U156; 
assign P3_SUB_357_1258_U131 = ~(P3_SUB_357_1258_U106 & P3_SUB_357_1258_U218); 
assign P3_SUB_357_1258_U230 = ~(P3_SUB_357_1258_U109 & P3_SUB_357_1258_U229); 
assign P3_SUB_357_1258_U231 = ~(P3_SUB_357_1258_U285 & P3_SUB_357_1258_U157); 
assign P3_SUB_357_1258_U242 = ~(P3_SUB_357_1258_U277 & P3_SUB_357_1258_U206); 
assign P3_SUB_357_1258_U391 = ~(P3_SUB_357_1258_U389 & P3_SUB_357_1258_U285); 
assign P3_SUB_357_1258_U398 = ~(P3_SUB_357_1258_U283 & P3_SUB_357_1258_U396); 
assign P3_SUB_357_1258_U405 = ~(P3_SUB_357_1258_U281 & P3_SUB_357_1258_U403); 
assign P3_SUB_357_1258_U412 = ~(P3_SUB_357_1258_U279 & P3_SUB_357_1258_U410); 
assign P3_SUB_357_1258_U431 = ~(P3_SUB_357_1258_U429 & P3_SUB_357_1258_U277); 
assign P3_ADD_515_U80 = ~(P3_ADD_515_U160 & P3_ADD_515_U159); 
assign P3_ADD_515_U113 = ~P3_ADD_515_U44; 
assign P3_ADD_515_U157 = ~(P3_ADD_515_U44 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_394_U79 = ~(P3_ADD_394_U162 & P3_ADD_394_U161); 
assign P3_ADD_394_U116 = ~P3_ADD_394_U44; 
assign P3_ADD_394_U159 = ~(P3_ADD_394_U44 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_441_U80 = ~(P3_ADD_441_U160 & P3_ADD_441_U159); 
assign P3_ADD_441_U113 = ~P3_ADD_441_U44; 
assign P3_ADD_441_U157 = ~(P3_ADD_441_U44 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_349_U84 = ~(P3_ADD_349_U167 & P3_ADD_349_U166); 
assign P3_ADD_349_U117 = ~P3_ADD_349_U45; 
assign P3_ADD_349_U164 = ~(P3_ADD_349_U45 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_405_U79 = ~(P3_ADD_405_U162 & P3_ADD_405_U161); 
assign P3_ADD_405_U116 = ~P3_ADD_405_U44; 
assign P3_ADD_405_U159 = ~(P3_ADD_405_U44 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_553_U84 = ~(P3_ADD_553_U167 & P3_ADD_553_U166); 
assign P3_ADD_553_U117 = ~P3_ADD_553_U45; 
assign P3_ADD_553_U164 = ~(P3_ADD_553_U45 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_558_U84 = ~(P3_ADD_558_U167 & P3_ADD_558_U166); 
assign P3_ADD_558_U117 = ~P3_ADD_558_U45; 
assign P3_ADD_558_U164 = ~(P3_ADD_558_U45 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_385_U84 = ~(P3_ADD_385_U167 & P3_ADD_385_U166); 
assign P3_ADD_385_U117 = ~P3_ADD_385_U45; 
assign P3_ADD_385_U164 = ~(P3_ADD_385_U45 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_547_U84 = ~(P3_ADD_547_U167 & P3_ADD_547_U166); 
assign P3_ADD_547_U117 = ~P3_ADD_547_U45; 
assign P3_ADD_547_U164 = ~(P3_ADD_547_U45 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_371_1212_U83 = ~(P3_ADD_371_1212_U257 & P3_ADD_371_1212_U256); 
assign P3_ADD_371_1212_U167 = ~P3_ADD_371_1212_U59; 
assign P3_ADD_371_1212_U185 = ~(P3_ADD_371_1212_U60 & P3_ADD_371_1212_U59); 
assign P3_ADD_371_1212_U187 = ~(P3_ADD_371_1212_U58 & P3_ADD_371_1212_U186); 
assign P3_ADD_494_U80 = ~(P3_ADD_494_U160 & P3_ADD_494_U159); 
assign P3_ADD_494_U113 = ~P3_ADD_494_U44; 
assign P3_ADD_494_U157 = ~(P3_ADD_494_U44 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_536_U80 = ~(P3_ADD_536_U160 & P3_ADD_536_U159); 
assign P3_ADD_536_U113 = ~P3_ADD_536_U44; 
assign P3_ADD_536_U157 = ~(P3_ADD_536_U44 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P2_R2099_U29 = ~(P2_U2736 & P2_R2099_U126); 
assign P2_R2099_U221 = ~(P2_R2099_U126 & P2_R2099_U28); 
assign P2_ADD_391_1196_U30 = ~(P2_ADD_391_1196_U39 & P2_ADD_391_1196_U180); 
assign P2_ADD_391_1196_U31 = ~P2_R2182_U71; 
assign P2_ADD_391_1196_U41 = ~P2_R2096_U92; 
assign P2_ADD_391_1196_U179 = ~P2_ADD_391_1196_U39; 
assign P2_ADD_391_1196_U188 = P2_R2182_U71 | P2_R2096_U70; 
assign P2_ADD_391_1196_U190 = ~(P2_R2096_U70 & P2_R2182_U71); 
assign P2_ADD_391_1196_U203 = ~(P2_ADD_391_1196_U114 & P2_ADD_391_1196_U177); 
assign P2_ADD_391_1196_U310 = ~(P2_R2182_U71 & P2_ADD_391_1196_U32); 
assign P2_ADD_391_1196_U312 = ~(P2_R2182_U71 & P2_ADD_391_1196_U32); 
assign P2_ADD_391_1196_U316 = ~(P2_R2096_U71 & P2_ADD_391_1196_U13); 
assign P2_ADD_391_1196_U320 = ~(P2_ADD_391_1196_U319 & P2_ADD_391_1196_U318); 
assign P2_SUB_563_U6 = ~P2_U3618; 
assign P2_SUB_563_U7 = ~P2_U3619; 
assign P2_R2182_U5 = P2_U2670 & P2_R2182_U4; 
assign P2_R2182_U70 = ~(P2_R2182_U194 & P2_R2182_U193); 
assign P2_R2182_U142 = ~P2_R2182_U4; 
assign P2_R2182_U300 = ~(P2_R2182_U33 & P2_R2182_U4); 
assign P2_R2182_U303 = ~(P2_R2182_U141 & P2_U2671); 
assign P2_R2027_U84 = ~(P2_R2027_U167 & P2_R2027_U166); 
assign P2_R2027_U117 = ~P2_R2027_U45; 
assign P2_R2027_U164 = ~(P2_R2027_U45 & P2_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P2_R2337_U78 = ~(P2_R2337_U158 & P2_R2337_U157); 
assign P2_R2337_U114 = ~P2_R2337_U45; 
assign P2_R2337_U155 = ~(P2_R2337_U45 & P2_PHYADDRPOINTER_REG_23__SCAN_IN); 
assign P2_R2096_U6 = P2_U2631 & P2_R2096_U25; 
assign P2_R2096_U91 = ~(P2_R2096_U251 & P2_R2096_U250); 
assign P2_R2096_U153 = ~P2_R2096_U25; 
assign P2_R2096_U246 = ~(P2_R2096_U26 & P2_R2096_U25); 
assign P2_R2096_U249 = ~(P2_R2096_U152 & P2_U2632); 
assign P2_LT_563_U7 = ~P2_U3620; 
assign P2_LT_563_U10 = ~P2_U3619; 
assign P2_LT_563_U11 = ~P2_U3618; 
assign P2_LT_563_U14 = ~P2_U3617; 
assign P2_LT_563_U15 = ~P2_U3621; 
assign P2_LT_563_U16 = ~(P2_U3620 & P2_LT_563_U8); 
assign P2_LT_563_U21 = ~(P2_U3619 & P2_LT_563_U9); 
assign P2_LT_563_U22 = ~(P2_U3618 & P2_LT_563_U12); 
assign P2_LT_563_U27 = ~(P2_U3617 & P2_LT_563_U13); 
assign P2_R2256_U36 = ~P2_R2256_U28; 
assign P2_R2256_U38 = ~(P2_R2256_U37 & P2_R2256_U28); 
assign P2_R2256_U46 = ~(P2_R2256_U66 & P2_R2256_U7); 
assign P2_R2256_U62 = ~(P2_R2256_U27 & P2_R2256_U28); 
assign P2_R1957_U32 = ~(P2_R1957_U97 & P2_R1957_U73 & P2_R1957_U43); 
assign P2_R2278_U53 = ~P2_U2809; 
assign P2_R2278_U55 = ~(P2_U2809 & P2_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P2_R2278_U121 = P2_R2278_U238 & P2_R2278_U242; 
assign P2_R2278_U203 = P2_R2278_U555 & P2_R2278_U554; 
assign P2_R2278_U245 = P2_U2809 | P2_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P2_R2278_U322 = ~(P2_R2278_U240 & P2_R2278_U242); 
assign P2_R2278_U541 = ~(P2_U2809 & P2_R2278_U54); 
assign P2_R2278_U543 = ~(P2_U2809 & P2_R2278_U54); 
assign P2_R2278_U547 = ~(P2_R2278_U47 & P2_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P2_R2278_U549 = ~(P2_R2278_U47 & P2_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P2_R2278_U558 = ~(P2_R2278_U557 & P2_R2278_U556); 
assign P2_ADD_394_U87 = ~(P2_ADD_394_U178 & P2_ADD_394_U177); 
assign P2_ADD_394_U116 = ~P2_ADD_394_U44; 
assign P2_ADD_394_U143 = ~(P2_ADD_394_U44 & P2_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P2_R2267_U83 = P2_R2267_U162 & P2_R2267_U161; 
assign P2_R2267_U104 = ~P2_R2267_U33; 
assign P2_R2267_U129 = ~(P2_U2782 & P2_R2267_U128); 
assign P2_R2267_U159 = ~(P2_U2781 & P2_R2267_U33); 
assign P2_ADD_371_1212_U137 = ~P2_ADD_371_1212_U29; 
assign P2_ADD_371_1212_U205 = ~(P2_ADD_371_1212_U27 & P2_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P2_ADD_371_1212_U265 = ~(P2_ADD_371_1212_U29 & P2_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P1_R2144_U94 = ~(P1_R2144_U143 & P1_R2144_U32); 
assign P1_R2144_U249 = ~(P1_R2144_U222 & P1_R2144_U143); 
assign P1_R2144_U251 = ~(P1_R2144_U142 & P1_R2144_U228); 
assign P1_R2278_U26 = ~P1_U2794; 
assign P1_R2278_U45 = ~P1_U2775; 
assign P1_R2278_U47 = ~P1_U2774; 
assign P1_R2278_U49 = ~P1_U2776; 
assign P1_R2278_U51 = ~P1_U2777; 
assign P1_R2278_U53 = ~P1_U2779; 
assign P1_R2278_U55 = ~P1_U2780; 
assign P1_R2278_U57 = ~P1_U2781; 
assign P1_R2278_U72 = ~P1_U2783; 
assign P1_R2278_U75 = ~P1_U2778; 
assign P1_R2278_U76 = ~(P1_U2778 & P1_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P1_R2278_U78 = ~P1_U2782; 
assign P1_R2278_U79 = ~(P1_U2782 & P1_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P1_R2278_U81 = ~P1_U2772; 
assign P1_R2278_U84 = ~P1_U2773; 
assign P1_R2278_U85 = ~(P1_U2773 & P1_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P1_R2278_U88 = ~P1_U2770; 
assign P1_R2278_U90 = ~P1_U2771; 
assign P1_R2278_U130 = P1_U2777 & P1_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P1_R2278_U133 = P1_U2781 & P1_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P1_R2278_U183 = P1_R2278_U456 & P1_R2278_U455; 
assign P1_R2278_U184 = ~(P1_R2278_U238 & P1_R2278_U237); 
assign P1_R2278_U186 = ~P1_U2769; 
assign P1_R2278_U187 = ~(P1_U2771 & P1_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P1_R2278_U231 = ~(P1_U2794 & P1_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P1_R2278_U254 = P1_U2794 | P1_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P1_R2278_U264 = P1_U2794 | P1_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P1_R2278_U269 = P1_U2794 | P1_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P1_R2278_U292 = P1_U2783 | P1_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P1_R2278_U293 = ~(P1_U2783 & P1_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P1_R2278_U295 = P1_U2782 | P1_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P1_R2278_U298 = P1_U2781 | P1_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P1_R2278_U300 = ~(P1_U2781 & P1_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P1_R2278_U302 = P1_U2780 | P1_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P1_R2278_U303 = ~(P1_U2780 & P1_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P1_R2278_U305 = P1_U2779 | P1_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P1_R2278_U306 = ~(P1_U2779 & P1_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P1_R2278_U308 = P1_U2778 | P1_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P1_R2278_U311 = P1_U2777 | P1_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P1_R2278_U312 = ~(P1_U2777 & P1_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P1_R2278_U313 = P1_U2776 | P1_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P1_R2278_U314 = ~(P1_U2776 & P1_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P1_R2278_U315 = P1_U2775 | P1_INSTADDRPOINTER_REG_25__SCAN_IN; 
assign P1_R2278_U316 = ~(P1_U2775 & P1_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P1_R2278_U317 = P1_U2774 | P1_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P1_R2278_U318 = ~(P1_U2774 & P1_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P1_R2278_U319 = P1_U2773 | P1_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P1_R2278_U321 = P1_U2772 | P1_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P1_R2278_U322 = ~(P1_U2772 & P1_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P1_R2278_U324 = P1_U2771 | P1_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P1_R2278_U327 = P1_U2770 | P1_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P1_R2278_U393 = ~(P1_U2770 & P1_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P1_R2278_U440 = ~(P1_R2278_U24 & P1_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P1_R2278_U441 = ~(P1_U2794 & P1_R2278_U25); 
assign P1_R2278_U447 = ~(P1_R2278_U28 & P1_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P1_R2278_U449 = ~(P1_R2278_U39 & P1_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P1_R2278_U451 = ~(P1_R2278_U39 & P1_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P1_R2278_U459 = ~(P1_R2278_U458 & P1_R2278_U457); 
assign P1_R2278_U463 = ~(P1_U2769 & P1_R2278_U185); 
assign P1_R2278_U465 = ~(P1_U2769 & P1_R2278_U185); 
assign P1_R2278_U472 = ~(P1_U2770 & P1_R2278_U89); 
assign P1_R2278_U474 = ~(P1_U2770 & P1_R2278_U89); 
assign P1_R2278_U483 = ~(P1_R2278_U191 & P1_R2278_U192); 
assign P1_R2278_U484 = ~(P1_R2278_U235 & P1_R2278_U482); 
assign P1_R2278_U486 = ~(P1_U2771 & P1_R2278_U91); 
assign P1_R2278_U488 = ~(P1_U2771 & P1_R2278_U91); 
assign P1_R2278_U493 = ~(P1_U2772 & P1_R2278_U82); 
assign P1_R2278_U495 = ~(P1_U2772 & P1_R2278_U82); 
assign P1_R2278_U499 = ~(P1_U2773 & P1_R2278_U83); 
assign P1_R2278_U501 = ~(P1_U2773 & P1_R2278_U83); 
assign P1_R2278_U506 = ~(P1_U2774 & P1_R2278_U46); 
assign P1_R2278_U508 = ~(P1_U2774 & P1_R2278_U46); 
assign P1_R2278_U513 = ~(P1_U2775 & P1_R2278_U44); 
assign P1_R2278_U515 = ~(P1_U2775 & P1_R2278_U44); 
assign P1_R2278_U520 = ~(P1_U2776 & P1_R2278_U48); 
assign P1_R2278_U522 = ~(P1_U2776 & P1_R2278_U48); 
assign P1_R2278_U527 = ~(P1_U2777 & P1_R2278_U50); 
assign P1_R2278_U529 = ~(P1_U2777 & P1_R2278_U50); 
assign P1_R2278_U534 = ~(P1_U2778 & P1_R2278_U74); 
assign P1_R2278_U536 = ~(P1_U2778 & P1_R2278_U74); 
assign P1_R2278_U541 = ~(P1_U2779 & P1_R2278_U52); 
assign P1_R2278_U543 = ~(P1_U2779 & P1_R2278_U52); 
assign P1_R2278_U548 = ~(P1_U2780 & P1_R2278_U54); 
assign P1_R2278_U550 = ~(P1_U2780 & P1_R2278_U54); 
assign P1_R2278_U560 = ~(P1_U2781 & P1_R2278_U56); 
assign P1_R2278_U562 = ~(P1_U2781 & P1_R2278_U56); 
assign P1_R2278_U567 = ~(P1_U2782 & P1_R2278_U77); 
assign P1_R2278_U569 = ~(P1_U2782 & P1_R2278_U77); 
assign P1_R2278_U574 = ~(P1_U2783 & P1_R2278_U71); 
assign P1_R2278_U576 = ~(P1_U2783 & P1_R2278_U71); 
assign P1_R2358_U33 = ~P1_U2642; 
assign P1_R2358_U37 = ~P1_U2623; 
assign P1_R2358_U38 = ~P1_U2624; 
assign P1_R2358_U39 = ~P1_U2625; 
assign P1_R2358_U40 = ~P1_U2626; 
assign P1_R2358_U41 = ~P1_U2627; 
assign P1_R2358_U43 = ~P1_U2628; 
assign P1_R2358_U44 = ~P1_U2629; 
assign P1_R2358_U45 = ~P1_U2630; 
assign P1_R2358_U46 = ~P1_U2631; 
assign P1_R2358_U48 = ~P1_U2632; 
assign P1_R2358_U49 = ~P1_U2633; 
assign P1_R2358_U62 = ~P1_U2622; 
assign P1_R2358_U63 = ~P1_U2620; 
assign P1_R2358_U64 = ~P1_U2621; 
assign P1_R2358_U81 = P1_R2358_U220 & P1_R2358_U219; 
assign P1_R2358_U83 = P1_R2358_U225 & P1_R2358_U28; 
assign P1_R2358_U122 = P1_R2358_U217 & P1_R2358_U216; 
assign P1_R2358_U168 = ~P1_U2663; 
assign P1_R2358_U213 = ~(P1_R2358_U121 & P1_R2358_U212); 
assign P1_R2358_U218 = ~(P1_R2358_U418 & P1_R2358_U417 & P1_R2358_U25); 
assign P1_R2358_U222 = ~(P1_R2358_U221 & P1_R2358_U219); 
assign P1_R2358_U228 = ~(P1_U2642 & P1_R2358_U448); 
assign P1_R2358_U241 = ~(P1_R2358_U217 & P1_R2358_U216); 
assign P1_R2358_U250 = ~P1_R2358_U66; 
assign P1_R2358_U251 = ~(P1_R2358_U66 & P1_R2358_U207); 
assign P1_R2358_U254 = ~(P1_R2358_U66 & P1_R2358_U207 & P1_R2358_U253); 
assign P1_R2358_U275 = ~(P1_U2633 & P1_R2358_U498); 
assign P1_R2358_U307 = ~(P1_R2358_U249 & P1_R2358_U306); 
assign P1_R2358_U334 = ~(P1_R2358_U220 & P1_R2358_U219); 
assign P1_R2358_U335 = ~(P1_R2358_U225 & P1_R2358_U28); 
assign P1_R2358_U495 = ~(P1_R2358_U494 & P1_R2358_U493); 
assign P1_R2358_U507 = ~(P1_U2663 & P1_R2358_U23); 
assign P1_R2358_U520 = ~(P1_U2663 & P1_R2358_U23); 
assign P1_R2099_U75 = ~(P1_R2099_U317 & P1_R2099_U316); 
assign P1_R2099_U172 = ~P1_R2099_U17; 
assign P1_R2099_U315 = ~(P1_R2099_U52 & P1_R2099_U17); 
assign P1_R2337_U80 = ~(P1_R2337_U160 & P1_R2337_U159); 
assign P1_R2337_U113 = ~P1_R2337_U44; 
assign P1_R2337_U157 = ~(P1_R2337_U44 & P1_PHYADDRPOINTER_REG_22__SCAN_IN); 
assign P1_R2096_U80 = ~(P1_R2096_U160 & P1_R2096_U159); 
assign P1_R2096_U113 = ~P1_R2096_U44; 
assign P1_R2096_U157 = ~(P1_R2096_U44 & P1_REIP_REG_22__SCAN_IN); 
assign P1_ADD_405_U87 = ~(P1_ADD_405_U178 & P1_ADD_405_U177); 
assign P1_ADD_405_U116 = ~P1_ADD_405_U44; 
assign P1_ADD_405_U143 = ~(P1_ADD_405_U44 & P1_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P1_ADD_515_U87 = ~(P1_ADD_515_U174 & P1_ADD_515_U173); 
assign P1_ADD_515_U113 = ~P1_ADD_515_U44; 
assign P1_ADD_515_U141 = ~(P1_ADD_515_U44 & P1_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_U2814 = ~(P3_U6534 & P3_U6533 & P3_U6535 & P3_U6536 & P3_U3970); 
assign P3_U2816 = ~(P3_U6518 & P3_U6517 & P3_U6520 & P3_U6519 & P3_U3968); 
assign P3_U2849 = ~(P3_U5967 & P3_U5965 & P3_U5966); 
assign P3_U3810 = P3_U3809 & P3_U3808 & P3_U6011; 
assign P3_U3820 = P3_U6046 & P3_U6045 & P3_U6047 & P3_U3821 & P3_U6041; 
assign P3_U3824 = P3_U3823 & P3_U3822 & P3_U6059; 
assign P3_U3825 = P3_U3826 & P3_U6065; 
assign P3_U3969 = P3_U6532 & P3_U6529 & P3_U6530 & P3_U6531; 
assign P3_U3971 = P3_U6548 & P3_U6545 & P3_U6546 & P3_U6547; 
assign P3_U4629 = ~(P3_U7953 & P3_U7952 & P3_STATE2_REG_2__SCAN_IN); 
assign P3_U5988 = ~(P3_U3802 & P3_U3799); 
assign P3_U6036 = ~(P3_U6018 & P3_U3815 & P3_U6016 & P3_U3812 & P3_U3818); 
assign P3_U6083 = ~(P3_ADD_371_1212_U83 & P3_U2360); 
assign P3_U6088 = ~(P3_ADD_360_1242_U9 & P3_U2395); 
assign P3_U6114 = ~(P3_ADD_558_U84 & P3_U3220); 
assign P3_U6115 = ~(P3_ADD_553_U84 & P3_U4298); 
assign P3_U6116 = ~(P3_ADD_547_U84 & P3_U4299); 
assign P3_U6119 = ~(P3_ADD_531_U84 & P3_U2354); 
assign P3_U6127 = ~(P3_ADD_385_U84 & P3_U2358); 
assign P3_U6128 = ~(P3_ADD_380_U84 & P3_U2359); 
assign P3_U6129 = ~(P3_ADD_349_U84 & P3_U4306); 
assign P3_U6130 = ~(P3_ADD_344_U84 & P3_U2362); 
assign P3_U6141 = ~(P3_ADD_541_U80 & P3_U4300); 
assign P3_U6142 = ~(P3_ADD_536_U80 & P3_U4301); 
assign P3_U6145 = ~(P3_ADD_515_U80 & P3_U4302); 
assign P3_U6146 = ~(P3_ADD_494_U80 & P3_U2356); 
assign P3_U6147 = ~(P3_ADD_476_U80 & P3_U4303); 
assign P3_U6148 = ~(P3_ADD_441_U80 & P3_U4304); 
assign P3_U6149 = ~(P3_ADD_405_U79 & P3_U4305); 
assign P3_U6150 = ~(P3_ADD_394_U79 & P3_U2357); 
assign P3_U6555 = ~(P3_U2387 & P3_ADD_371_1212_U83); 
assign P3_U6559 = ~(P3_U2396 & P3_ADD_360_1242_U9); 
assign P3_U6573 = ~(P3_ADD_318_U80 & P3_U2398); 
assign P3_U6578 = ~(P3_ADD_339_U80 & P3_U2388); 
assign P3_U6582 = ~(P3_ADD_315_U76 & P3_U2397); 
assign P3_U7278 = ~(P3_ADD_467_U80 & P3_U2601); 
assign P3_U7280 = ~(P3_ADD_430_U80 & P3_U2405); 
assign P2_U2493 = P2_U3427 & P2_U3425; 
assign P2_U2495 = P2_U3440 & P2_U5174; 
assign P2_U2497 = P2_U3451 & P2_U5232; 
assign P2_U2499 = P2_U3463 & P2_U5289; 
assign P2_U2505 = P2_U3474 & P2_U5347; 
assign P2_U2507 = P2_U3486 & P2_U5404; 
assign P2_U2509 = P2_U3497 & P2_U5462; 
assign P2_U2511 = P2_U3509 & P2_U5519; 
assign P2_U2807 = P2_U3242 & P2_R2267_U83; 
assign P2_U2879 = ~(P2_U6496 & P2_U6497 & P2_U6495); 
assign P2_U2915 = ~(P2_U6344 & P2_U6343 & P2_U4063); 
assign P2_U2916 = ~(P2_U6340 & P2_U6339 & P2_U4062); 
assign P2_U2917 = ~(P2_U6336 & P2_U6335 & P2_U4061); 
assign P2_U2918 = ~(P2_U6332 & P2_U6331 & P2_U4060); 
assign P2_U2919 = ~(P2_U6328 & P2_U6327 & P2_U4059); 
assign P2_U3595 = ~(P2_U8073 & P2_U8072); 
assign P2_U3596 = ~(P2_U8084 & P2_U8083); 
assign P2_U4071 = P2_U6577 & P2_U6576; 
assign P2_U4075 = P2_U6586 & P2_U6585; 
assign P2_U4079 = P2_U6595 & P2_U6594; 
assign P2_U4083 = P2_U6604 & P2_U6603; 
assign P2_U4658 = ~(P2_U2468 & P2_U2362); 
assign P2_U4664 = ~(P2_U2468 & P2_U2398); 
assign P2_U4671 = ~(P2_U2421 & P2_U4641); 
assign P2_U4676 = ~(P2_U2419 & P2_U4641); 
assign P2_U4681 = ~(P2_U2417 & P2_U4641); 
assign P2_U4686 = ~(P2_U2415 & P2_U4641); 
assign P2_U4691 = ~(P2_U2413 & P2_U4641); 
assign P2_U4696 = ~(P2_U2411 & P2_U4641); 
assign P2_U4701 = ~(P2_U2409 & P2_U4641); 
assign P2_U4706 = ~(P2_U2407 & P2_U4641); 
assign P2_U4716 = ~(P2_U2471 & P2_U2362); 
assign P2_U4722 = ~(P2_U2471 & P2_U2398); 
assign P2_U4729 = ~(P2_U4710 & P2_U2421); 
assign P2_U4734 = ~(P2_U4710 & P2_U2419); 
assign P2_U4739 = ~(P2_U4710 & P2_U2417); 
assign P2_U4744 = ~(P2_U4710 & P2_U2415); 
assign P2_U4749 = ~(P2_U4710 & P2_U2413); 
assign P2_U4754 = ~(P2_U4710 & P2_U2411); 
assign P2_U4759 = ~(P2_U4710 & P2_U2409); 
assign P2_U4764 = ~(P2_U4710 & P2_U2407); 
assign P2_U4775 = ~(P2_U2474 & P2_U2362); 
assign P2_U4781 = ~(P2_U2474 & P2_U2398); 
assign P2_U4788 = ~(P2_U4768 & P2_U2421); 
assign P2_U4793 = ~(P2_U4768 & P2_U2419); 
assign P2_U4798 = ~(P2_U4768 & P2_U2417); 
assign P2_U4803 = ~(P2_U4768 & P2_U2415); 
assign P2_U4808 = ~(P2_U4768 & P2_U2413); 
assign P2_U4813 = ~(P2_U4768 & P2_U2411); 
assign P2_U4818 = ~(P2_U4768 & P2_U2409); 
assign P2_U4823 = ~(P2_U4768 & P2_U2407); 
assign P2_U4832 = ~(P2_U2480 & P2_U2362); 
assign P2_U4838 = ~(P2_U2480 & P2_U2398); 
assign P2_U4845 = ~(P2_U4826 & P2_U2421); 
assign P2_U4850 = ~(P2_U4826 & P2_U2419); 
assign P2_U4855 = ~(P2_U4826 & P2_U2417); 
assign P2_U4860 = ~(P2_U4826 & P2_U2415); 
assign P2_U4865 = ~(P2_U4826 & P2_U2413); 
assign P2_U4870 = ~(P2_U4826 & P2_U2411); 
assign P2_U4875 = ~(P2_U4826 & P2_U2409); 
assign P2_U4880 = ~(P2_U4826 & P2_U2407); 
assign P2_U4890 = ~(P2_U2484 & P2_U2362); 
assign P2_U4896 = ~(P2_U2484 & P2_U2398); 
assign P2_U4903 = ~(P2_U4883 & P2_U2421); 
assign P2_U4908 = ~(P2_U4883 & P2_U2419); 
assign P2_U4913 = ~(P2_U4883 & P2_U2417); 
assign P2_U4918 = ~(P2_U4883 & P2_U2415); 
assign P2_U4923 = ~(P2_U4883 & P2_U2413); 
assign P2_U4928 = ~(P2_U4883 & P2_U2411); 
assign P2_U4933 = ~(P2_U4883 & P2_U2409); 
assign P2_U4938 = ~(P2_U4883 & P2_U2407); 
assign P2_U4947 = ~(P2_U2486 & P2_U2362); 
assign P2_U4953 = ~(P2_U2486 & P2_U2398); 
assign P2_U4960 = ~(P2_U4941 & P2_U2421); 
assign P2_U4965 = ~(P2_U4941 & P2_U2419); 
assign P2_U4970 = ~(P2_U4941 & P2_U2417); 
assign P2_U4975 = ~(P2_U4941 & P2_U2415); 
assign P2_U4980 = ~(P2_U4941 & P2_U2413); 
assign P2_U4985 = ~(P2_U4941 & P2_U2411); 
assign P2_U4990 = ~(P2_U4941 & P2_U2409); 
assign P2_U4995 = ~(P2_U4941 & P2_U2407); 
assign P2_U5005 = ~(P2_U2488 & P2_U2362); 
assign P2_U5011 = ~(P2_U2488 & P2_U2398); 
assign P2_U5018 = ~(P2_U4998 & P2_U2421); 
assign P2_U5023 = ~(P2_U4998 & P2_U2419); 
assign P2_U5028 = ~(P2_U4998 & P2_U2417); 
assign P2_U5033 = ~(P2_U4998 & P2_U2415); 
assign P2_U5038 = ~(P2_U4998 & P2_U2413); 
assign P2_U5043 = ~(P2_U4998 & P2_U2411); 
assign P2_U5048 = ~(P2_U4998 & P2_U2409); 
assign P2_U5053 = ~(P2_U4998 & P2_U2407); 
assign P2_U5062 = ~(P2_U2490 & P2_U2362); 
assign P2_U5068 = ~(P2_U2490 & P2_U2398); 
assign P2_U5075 = ~(P2_U5056 & P2_U2421); 
assign P2_U5080 = ~(P2_U5056 & P2_U2419); 
assign P2_U5085 = ~(P2_U5056 & P2_U2417); 
assign P2_U5090 = ~(P2_U5056 & P2_U2415); 
assign P2_U5095 = ~(P2_U5056 & P2_U2413); 
assign P2_U5100 = ~(P2_U5056 & P2_U2411); 
assign P2_U5105 = ~(P2_U5056 & P2_U2409); 
assign P2_U5110 = ~(P2_U5056 & P2_U2407); 
assign P2_U5113 = ~P2_U3427; 
assign P2_U5169 = ~P2_U3440; 
assign P2_U5226 = ~P2_U3451; 
assign P2_U5284 = ~P2_U3463; 
assign P2_U5341 = ~P2_U3474; 
assign P2_U5399 = ~P2_U3486; 
assign P2_U5456 = ~P2_U3497; 
assign P2_U5514 = ~P2_U3509; 
assign P2_U5647 = ~(P2_U3427 & P2_U5646); 
assign P2_U6394 = ~(P2_U2380 & P2_R2096_U91); 
assign P2_U6498 = ~(P2_R2182_U70 & P2_U2393); 
assign P2_U6573 = ~(P2_R2267_U21 & P2_U2587); 
assign P2_U6574 = ~(P2_U2588 & P2_R2096_U68); 
assign P2_U6582 = ~(P2_R2267_U43 & P2_U2587); 
assign P2_U6583 = ~(P2_U2588 & P2_R2096_U51); 
assign P2_U6591 = ~(P2_R2267_U65 & P2_U2587); 
assign P2_U6592 = ~(P2_U2588 & P2_R2096_U77); 
assign P2_U6600 = ~(P2_R2267_U17 & P2_U2587); 
assign P2_U6601 = ~(P2_U2588 & P2_R2096_U75); 
assign P2_U6609 = ~(P2_R2267_U60 & P2_U2587); 
assign P2_U6610 = ~(P2_U2588 & P2_R2096_U74); 
assign P2_U6618 = ~(P2_R2267_U18 & P2_U2587); 
assign P2_U6619 = ~(P2_U2588 & P2_R2096_U73); 
assign P2_U6627 = ~(P2_R2267_U58 & P2_U2587); 
assign P2_U6628 = ~(P2_U2588 & P2_R2096_U72); 
assign P2_U6635 = ~(P2_R2267_U19 & P2_U2587); 
assign P2_U6636 = ~(P2_U2588 & P2_R2096_U71); 
assign P2_U6643 = ~(P2_R2267_U56 & P2_U2587); 
assign P2_U6644 = ~(P2_U2588 & P2_R2096_U70); 
assign P2_U6651 = ~(P2_R2267_U20 & P2_U2587); 
assign P2_U6652 = ~(P2_U2588 & P2_R2096_U69); 
assign P2_U6659 = ~(P2_R2267_U87 & P2_U2587); 
assign P2_U6660 = ~(P2_U2588 & P2_R2096_U97); 
assign P2_U6667 = ~(P2_R2267_U6 & P2_U2587); 
assign P2_U6668 = ~(P2_U2588 & P2_R2096_U96); 
assign P2_U6675 = ~(P2_R2267_U85 & P2_U2587); 
assign P2_U6676 = ~(P2_U2588 & P2_R2096_U95); 
assign P2_U6683 = ~(P2_R2267_U7 & P2_U2587); 
assign P2_U6684 = ~(P2_U2588 & P2_R2096_U94); 
assign P2_U6691 = ~(P2_R2267_U83 & P2_U2587); 
assign P2_U6692 = ~(P2_U2588 & P2_R2096_U93); 
assign P2_U6700 = ~(P2_U2588 & P2_R2096_U92); 
assign P2_U6708 = ~(P2_U2588 & P2_R2096_U91); 
assign P2_U7743 = ~(P2_U7741 & P2_U4448 & P2_U7742); 
assign P2_U8391 = ~(P2_R2337_U78 & P2_U3284); 
assign P1_U2499 = P1_U4531 & P1_U3454; 
assign P1_U2507 = P1_U4531 & P1_U7693; 
assign P1_U2662 = ~(P1_U6816 & P1_U4020); 
assign P1_U2871 = ~(P1_U6269 & P1_U6270 & P1_U6268); 
assign P1_U2903 = ~(P1_U6158 & P1_U6157 & P1_U6159); 
assign P1_U2998 = ~(P1_U5805 & P1_U5804 & P1_U5806 & P1_U5808 & P1_U5807); 
assign P1_U3032 = P1_U5537 & P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign P1_U3315 = ~(P1_U4527 & P1_U2475); 
assign P1_U3327 = ~(P1_U4600 & P1_U2475); 
assign P1_U3334 = ~(P1_U4658 & P1_U2475); 
assign P1_U3338 = ~(P1_U2485 & P1_U2475); 
assign P1_U3343 = ~(P1_U2490 & P1_U4527); 
assign P1_U3347 = ~(P1_U2490 & P1_U4600); 
assign P1_U3350 = ~(P1_U2490 & P1_U4658); 
assign P1_U3354 = ~(P1_U2490 & P1_U2485); 
assign P1_U3768 = P1_U5580 & P1_U5579; 
assign P1_U5546 = ~(P1_U2388 & P1_U7733); 
assign P1_U5710 = ~(P1_R2099_U75 & P1_U2380); 
assign P1_U5720 = ~(P1_ADD_405_U87 & P1_U2375); 
assign P1_U5721 = ~(P1_ADD_515_U87 & P1_U2374); 
assign P1_U5904 = ~(P1_R2337_U80 & P1_U2376); 
assign P1_U6326 = ~(P1_U2371 & P1_R2099_U75); 
assign P1_U6514 = ~(P1_U2604 & P1_R2099_U75); 
assign P1_U6522 = ~(P1_R2096_U80 & P1_U7485); 
assign P1_U6815 = ~(P1_R2337_U80 & P1_U2352); 
assign P1_U7683 = ~(P1_U4512 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U7729 = ~(P1_U5537 & P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P1_U7734 = ~(P1_U5537 & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P1_U7736 = ~(P1_U5537 & P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P1_U7737 = ~(P1_U5554 & P1_U3404); 
assign P1_U7738 = ~(P1_U5537 & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P1_U7739 = ~(P1_U5557 & P1_U3404); 
assign P3_ADD_476_U46 = ~(P3_ADD_476_U113 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_476_U158 = ~(P3_ADD_476_U113 & P3_ADD_476_U45); 
assign P3_ADD_531_U47 = ~(P3_ADD_531_U117 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_531_U165 = ~(P3_ADD_531_U117 & P3_ADD_531_U46); 
assign P3_SUB_320_U11 = P3_SUB_320_U116 & P3_SUB_320_U33; 
assign P3_SUB_320_U69 = ~P3_ADD_318_U80; 
assign P3_SUB_320_U98 = ~P3_SUB_320_U33; 
assign P3_SUB_320_U146 = ~(P3_ADD_318_U80 & P3_SUB_320_U33); 
assign P3_ADD_318_U46 = ~(P3_ADD_318_U113 & P3_PHYADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_318_U158 = ~(P3_ADD_318_U113 & P3_ADD_318_U45); 
assign P3_ADD_315_U46 = ~(P3_ADD_315_U110 & P3_PHYADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_315_U150 = ~(P3_ADD_315_U110 & P3_ADD_315_U45); 
assign P3_ADD_360_1242_U10 = P3_ADD_360_1242_U175 & P3_ADD_360_1242_U58; 
assign P3_ADD_360_1242_U159 = ~P3_ADD_360_1242_U58; 
assign P3_ADD_360_1242_U174 = ~(P3_ADD_360_1242_U59 & P3_ADD_360_1242_U58); 
assign P3_ADD_467_U46 = ~(P3_ADD_467_U113 & P3_REIP_REG_22__SCAN_IN); 
assign P3_ADD_467_U158 = ~(P3_ADD_467_U113 & P3_ADD_467_U45); 
assign P3_ADD_430_U46 = ~(P3_ADD_430_U113 & P3_REIP_REG_22__SCAN_IN); 
assign P3_ADD_430_U158 = ~(P3_ADD_430_U113 & P3_ADD_430_U45); 
assign P3_ADD_380_U47 = ~(P3_ADD_380_U117 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_380_U165 = ~(P3_ADD_380_U117 & P3_ADD_380_U46); 
assign P3_ADD_344_U47 = ~(P3_ADD_344_U117 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_344_U165 = ~(P3_ADD_344_U117 & P3_ADD_344_U46); 
assign P3_ADD_339_U46 = ~(P3_ADD_339_U113 & P3_PHYADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_339_U158 = ~(P3_ADD_339_U113 & P3_ADD_339_U45); 
assign P3_ADD_541_U46 = ~(P3_ADD_541_U113 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_541_U158 = ~(P3_ADD_541_U113 & P3_ADD_541_U45); 
assign P3_SUB_357_1258_U81 = ~(P3_SUB_357_1258_U391 & P3_SUB_357_1258_U390); 
assign P3_SUB_357_1258_U82 = ~(P3_SUB_357_1258_U398 & P3_SUB_357_1258_U397); 
assign P3_SUB_357_1258_U83 = ~(P3_SUB_357_1258_U405 & P3_SUB_357_1258_U404); 
assign P3_SUB_357_1258_U84 = ~(P3_SUB_357_1258_U412 & P3_SUB_357_1258_U411); 
assign P3_SUB_357_1258_U86 = ~(P3_SUB_357_1258_U431 & P3_SUB_357_1258_U430); 
assign P3_SUB_357_1258_U220 = ~P3_SUB_357_1258_U131; 
assign P3_SUB_357_1258_U221 = ~P3_SUB_357_1258_U62; 
assign P3_SUB_357_1258_U233 = ~(P3_SUB_357_1258_U110 & P3_SUB_357_1258_U231); 
assign P3_SUB_357_1258_U235 = ~P3_SUB_357_1258_U65; 
assign P3_SUB_357_1258_U236 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U65); 
assign P3_SUB_357_1258_U244 = ~(P3_SUB_357_1258_U112 & P3_SUB_357_1258_U242); 
assign P3_SUB_357_1258_U274 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U62); 
assign P3_SUB_357_1258_U302 = ~(P3_SUB_357_1258_U131 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_SUB_357_1258_U304 = ~(P3_SUB_357_1258_U4 & P3_SUB_357_1258_U131); 
assign P3_SUB_357_1258_U306 = ~(P3_SUB_357_1258_U4 & P3_SUB_357_1258_U131); 
assign P3_SUB_357_1258_U383 = ~(P3_SUB_357_1258_U130 & P3_SUB_357_1258_U131); 
assign P3_ADD_515_U46 = ~(P3_ADD_515_U113 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_515_U158 = ~(P3_ADD_515_U113 & P3_ADD_515_U45); 
assign P3_ADD_394_U46 = ~(P3_ADD_394_U116 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_394_U160 = ~(P3_ADD_394_U116 & P3_ADD_394_U45); 
assign P3_ADD_441_U46 = ~(P3_ADD_441_U113 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_441_U158 = ~(P3_ADD_441_U113 & P3_ADD_441_U45); 
assign P3_ADD_349_U47 = ~(P3_ADD_349_U117 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_349_U165 = ~(P3_ADD_349_U117 & P3_ADD_349_U46); 
assign P3_ADD_405_U46 = ~(P3_ADD_405_U116 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_405_U160 = ~(P3_ADD_405_U116 & P3_ADD_405_U45); 
assign P3_ADD_553_U47 = ~(P3_ADD_553_U117 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_553_U165 = ~(P3_ADD_553_U117 & P3_ADD_553_U46); 
assign P3_ADD_558_U47 = ~(P3_ADD_558_U117 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_558_U165 = ~(P3_ADD_558_U117 & P3_ADD_558_U46); 
assign P3_ADD_385_U47 = ~(P3_ADD_385_U117 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_385_U165 = ~(P3_ADD_385_U117 & P3_ADD_385_U46); 
assign P3_ADD_547_U47 = ~(P3_ADD_547_U117 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_547_U165 = ~(P3_ADD_547_U117 & P3_ADD_547_U46); 
assign P3_ADD_371_1212_U10 = P3_ADD_371_1212_U187 & P3_ADD_371_1212_U59; 
assign P3_ADD_371_1212_U62 = ~(P3_ADD_371_1212_U104 & P3_ADD_371_1212_U167); 
assign P3_ADD_371_1212_U168 = ~(P3_ADD_371_1212_U167 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_ADD_494_U46 = ~(P3_ADD_494_U113 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_494_U158 = ~(P3_ADD_494_U113 & P3_ADD_494_U45); 
assign P3_ADD_536_U46 = ~(P3_ADD_536_U113 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_536_U158 = ~(P3_ADD_536_U113 & P3_ADD_536_U45); 
assign P2_R2099_U92 = ~(P2_R2099_U221 & P2_R2099_U220); 
assign P2_R2099_U127 = ~P2_R2099_U29; 
assign P2_R2099_U218 = ~(P2_U2735 & P2_R2099_U29); 
assign P2_ADD_391_1196_U34 = ~P2_R2182_U70; 
assign P2_ADD_391_1196_U55 = ~P2_R2096_U91; 
assign P2_ADD_391_1196_U113 = P2_ADD_391_1196_U317 & P2_ADD_391_1196_U316; 
assign P2_ADD_391_1196_U181 = ~P2_ADD_391_1196_U30; 
assign P2_ADD_391_1196_U193 = P2_R2096_U69 | P2_R2182_U70; 
assign P2_ADD_391_1196_U195 = ~(P2_R2182_U70 & P2_R2096_U69); 
assign P2_ADD_391_1196_U198 = ~(P2_ADD_391_1196_U197 & P2_ADD_391_1196_U30); 
assign P2_ADD_391_1196_U205 = ~(P2_ADD_391_1196_U179 & P2_ADD_391_1196_U204); 
assign P2_ADD_391_1196_U206 = ~(P2_R2182_U70 & P2_R2096_U69); 
assign P2_ADD_391_1196_U308 = ~(P2_R2182_U70 & P2_ADD_391_1196_U33); 
assign P2_ADD_391_1196_U309 = ~(P2_R2096_U70 & P2_ADD_391_1196_U31); 
assign P2_ADD_391_1196_U311 = ~(P2_R2096_U70 & P2_ADD_391_1196_U31); 
assign P2_ADD_391_1196_U321 = ~(P2_ADD_391_1196_U303 & P2_ADD_391_1196_U30); 
assign P2_R2182_U6 = P2_U2669 & P2_R2182_U5; 
assign P2_R2182_U96 = ~(P2_R2182_U303 & P2_R2182_U302); 
assign P2_R2182_U143 = ~P2_R2182_U5; 
assign P2_R2182_U298 = ~(P2_R2182_U39 & P2_R2182_U5); 
assign P2_R2182_U301 = ~(P2_R2182_U142 & P2_U2670); 
assign P2_R2027_U47 = ~(P2_R2027_U117 & P2_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P2_R2027_U165 = ~(P2_R2027_U117 & P2_R2027_U46); 
assign P2_LT_563_1260_U7 = ~(P2_SUB_563_U6 | P2_SUB_563_U7); 
assign P2_R2337_U47 = ~(P2_R2337_U114 & P2_PHYADDRPOINTER_REG_23__SCAN_IN); 
assign P2_R2337_U156 = ~(P2_R2337_U114 & P2_R2337_U46); 
assign P2_R2096_U16 = P2_U2630 & P2_R2096_U6; 
assign P2_R2096_U90 = ~(P2_R2096_U249 & P2_R2096_U248); 
assign P2_R2096_U154 = ~P2_R2096_U6; 
assign P2_R2096_U244 = ~(P2_R2096_U47 & P2_R2096_U6); 
assign P2_R2096_U247 = ~(P2_R2096_U153 & P2_U2631); 
assign P2_LT_563_U17 = ~(P2_LT_563_U15 & P2_LT_563_U16 & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P2_LT_563_U18 = ~(P2_LT_563_U7 & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P2_LT_563_U19 = ~(P2_LT_563_U10 & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P2_LT_563_U24 = ~(P2_LT_563_U11 & P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P2_LT_563_U25 = ~(P2_LT_563_U14 & P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign P2_R2256_U4 = ~(P2_R2256_U31 & P2_R2256_U46); 
assign P2_R2256_U25 = ~(P2_R2256_U39 & P2_R2256_U38); 
assign P2_R2256_U63 = ~(P2_R2256_U36 & P2_R2256_U61); 
assign P2_R1957_U11 = P2_R1957_U116 & P2_R1957_U32; 
assign P2_R1957_U69 = ~P2_U3669; 
assign P2_R1957_U98 = ~P2_R1957_U32; 
assign P2_R1957_U146 = ~(P2_U3669 & P2_R1957_U32); 
assign P2_R2278_U13 = ~P2_U3638; 
assign P2_R2278_U15 = ~(P2_U3638 & P2_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P2_R2278_U45 = ~P2_U2808; 
assign P2_R2278_U122 = P2_R2278_U322 & P2_R2278_U243; 
assign P2_R2278_U201 = P2_R2278_U548 & P2_R2278_U547; 
assign P2_R2278_U247 = ~P2_R2278_U55; 
assign P2_R2278_U249 = P2_U2808 | P2_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P2_R2278_U250 = ~(P2_U2808 & P2_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P2_R2278_U534 = ~(P2_U2808 & P2_R2278_U46); 
assign P2_R2278_U536 = ~(P2_U2808 & P2_R2278_U46); 
assign P2_R2278_U540 = ~(P2_R2278_U53 & P2_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P2_R2278_U542 = ~(P2_R2278_U53 & P2_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P2_R2278_U551 = ~(P2_R2278_U550 & P2_R2278_U549); 
assign P2_R2278_U562 = ~(P2_U3638 & P2_R2278_U14); 
assign P2_ADD_394_U46 = ~(P2_ADD_394_U116 & P2_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P2_ADD_394_U144 = ~(P2_ADD_394_U116 & P2_ADD_394_U45); 
assign P2_R2267_U8 = P2_R2267_U129 & P2_R2267_U33; 
assign P2_R2267_U34 = ~(P2_R2267_U48 & P2_R2267_U104); 
assign P2_R2267_U126 = ~(P2_R2267_U104 & P2_R2267_U80); 
assign P2_R2267_U160 = ~(P2_R2267_U104 & P2_R2267_U80); 
assign P2_ADD_371_1212_U68 = ~(P2_ADD_371_1212_U206 & P2_ADD_371_1212_U205); 
assign P2_ADD_371_1212_U266 = ~(P2_ADD_371_1212_U137 & P2_ADD_371_1212_U28); 
assign P1_R2144_U38 = ~(P1_R2144_U250 & P1_R2144_U249); 
assign P1_R2144_U39 = ~(P1_R2144_U252 & P1_R2144_U251); 
assign P1_R2144_U147 = ~P1_R2144_U94; 
assign P1_R2144_U248 = ~(P1_R2144_U31 & P1_R2144_U94); 
assign P1_R2278_U8 = P1_R2278_U302 & P1_R2278_U298 & P1_R2278_U305; 
assign P1_R2278_U10 = P1_R2278_U313 & P1_R2278_U311 & P1_R2278_U315; 
assign P1_R2278_U12 = P1_R2278_U295 & P1_R2278_U292; 
assign P1_R2278_U22 = ~P1_U2792; 
assign P1_R2278_U59 = ~P1_U2789; 
assign P1_R2278_U61 = ~P1_U2790; 
assign P1_R2278_U68 = ~(P1_U2788 & P1_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P1_R2278_U70 = ~P1_U2784; 
assign P1_R2278_U107 = ~(P1_R2278_U484 & P1_R2278_U483); 
assign P1_R2278_U131 = P1_R2278_U318 & P1_R2278_U316; 
assign P1_R2278_U132 = P1_R2278_U319 & P1_R2278_U317 & P1_R2278_U321; 
assign P1_R2278_U134 = P1_R2278_U319 & P1_R2278_U317; 
assign P1_R2278_U135 = P1_R2278_U321 & P1_R2278_U308; 
assign P1_R2278_U148 = P1_R2278_U324 & P1_R2278_U321 & P1_R2278_U319 & P1_R2278_U317; 
assign P1_R2278_U149 = P1_R2278_U321 & P1_R2278_U308 & P1_R2278_U324; 
assign P1_R2278_U154 = P1_R2278_U324 & P1_R2278_U321; 
assign P1_R2278_U166 = P1_R2278_U311 & P1_R2278_U313; 
assign P1_R2278_U171 = P1_R2278_U298 & P1_R2278_U302; 
assign P1_R2278_U179 = P1_R2278_U440 & P1_R2278_U439; 
assign P1_R2278_U180 = P1_R2278_U447 & P1_R2278_U446; 
assign P1_R2278_U181 = P1_R2278_U449 & P1_R2278_U448; 
assign P1_R2278_U228 = ~(P1_U2790 & P1_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P1_R2278_U239 = ~P1_R2278_U184; 
assign P1_R2278_U241 = ~(P1_R2278_U240 & P1_R2278_U184); 
assign P1_R2278_U258 = P1_U2792 | P1_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P1_R2278_U259 = ~(P1_U2792 & P1_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P1_R2278_U261 = P1_U2791 | P1_INSTADDRPOINTER_REG_9__SCAN_IN; 
assign P1_R2278_U262 = ~(P1_U2791 & P1_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P1_R2278_U263 = ~(P1_U2791 & P1_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P1_R2278_U273 = ~(P1_U2791 & P1_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P1_R2278_U276 = P1_U2789 | P1_INSTADDRPOINTER_REG_11__SCAN_IN; 
assign P1_R2278_U277 = P1_U2790 | P1_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P1_R2278_U279 = ~(P1_U2789 & P1_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P1_R2278_U281 = P1_U2788 | P1_INSTADDRPOINTER_REG_12__SCAN_IN; 
assign P1_R2278_U288 = P1_U2784 | P1_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P1_R2278_U290 = ~(P1_U2784 & P1_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P1_R2278_U296 = ~P1_R2278_U79; 
assign P1_R2278_U309 = ~P1_R2278_U76; 
assign P1_R2278_U320 = ~P1_R2278_U85; 
assign P1_R2278_U325 = ~P1_R2278_U187; 
assign P1_R2278_U340 = P1_U2790 | P1_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P1_R2278_U343 = ~(P1_U2789 & P1_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P1_R2278_U345 = P1_U2790 | P1_INSTADDRPOINTER_REG_10__SCAN_IN; 
assign P1_R2278_U347 = ~(P1_R2278_U269 & P1_R2278_U231); 
assign P1_R2278_U364 = ~(P1_R2278_U133 & P1_R2278_U302); 
assign P1_R2278_U370 = ~(P1_R2278_U130 & P1_R2278_U313); 
assign P1_R2278_U432 = ~(P1_U2792 & P1_R2278_U21); 
assign P1_R2278_U434 = ~(P1_U2792 & P1_R2278_U21); 
assign P1_R2278_U442 = ~(P1_R2278_U26 & P1_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P1_R2278_U452 = ~(P1_R2278_U451 & P1_R2278_U450); 
assign P1_R2278_U460 = ~(P1_R2278_U183 & P1_R2278_U184); 
assign P1_R2278_U462 = ~(P1_R2278_U186 & P1_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P1_R2278_U464 = ~(P1_R2278_U186 & P1_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P1_R2278_U471 = ~(P1_R2278_U88 & P1_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P1_R2278_U473 = ~(P1_R2278_U88 & P1_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P1_R2278_U485 = ~(P1_R2278_U90 & P1_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P1_R2278_U487 = ~(P1_R2278_U90 & P1_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P1_R2278_U492 = ~(P1_R2278_U81 & P1_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P1_R2278_U494 = ~(P1_R2278_U81 & P1_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P1_R2278_U500 = ~(P1_R2278_U84 & P1_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P1_R2278_U502 = ~(P1_R2278_U84 & P1_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P1_R2278_U507 = ~(P1_R2278_U47 & P1_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P1_R2278_U509 = ~(P1_R2278_U47 & P1_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P1_R2278_U514 = ~(P1_R2278_U45 & P1_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P1_R2278_U516 = ~(P1_R2278_U45 & P1_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P1_R2278_U521 = ~(P1_R2278_U49 & P1_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P1_R2278_U523 = ~(P1_R2278_U49 & P1_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P1_R2278_U528 = ~(P1_R2278_U51 & P1_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P1_R2278_U530 = ~(P1_R2278_U51 & P1_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P1_R2278_U535 = ~(P1_R2278_U75 & P1_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P1_R2278_U537 = ~(P1_R2278_U75 & P1_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P1_R2278_U542 = ~(P1_R2278_U53 & P1_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P1_R2278_U544 = ~(P1_R2278_U53 & P1_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P1_R2278_U549 = ~(P1_R2278_U55 & P1_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P1_R2278_U551 = ~(P1_R2278_U55 & P1_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P1_R2278_U561 = ~(P1_R2278_U57 & P1_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P1_R2278_U563 = ~(P1_R2278_U57 & P1_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P1_R2278_U568 = ~(P1_R2278_U78 & P1_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P1_R2278_U570 = ~(P1_R2278_U78 & P1_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P1_R2278_U575 = ~(P1_R2278_U72 & P1_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P1_R2278_U577 = ~(P1_R2278_U72 & P1_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P1_R2278_U581 = ~(P1_U2784 & P1_R2278_U69); 
assign P1_R2278_U583 = ~(P1_U2784 & P1_R2278_U69); 
assign P1_R2278_U602 = ~(P1_U2789 & P1_R2278_U58); 
assign P1_R2278_U604 = ~(P1_U2790 & P1_R2278_U60); 
assign P1_R2358_U34 = ~P1_U2641; 
assign P1_R2358_U50 = ~P1_U2634; 
assign P1_R2358_U51 = ~(P1_U2634 & P1_R2358_U501); 
assign P1_R2358_U52 = ~P1_U2639; 
assign P1_R2358_U53 = ~P1_U2640; 
assign P1_R2358_U56 = ~P1_U2638; 
assign P1_R2358_U57 = ~(P1_U2638 & P1_R2358_U471); 
assign P1_R2358_U156 = ~(P1_R2358_U203 & P1_R2358_U213); 
assign P1_R2358_U223 = ~(P1_R2358_U220 & P1_R2358_U222 & P1_R2358_U215); 
assign P1_R2358_U229 = ~(P1_R2358_U445 & P1_R2358_U444 & P1_R2358_U33); 
assign P1_R2358_U233 = ~(P1_U2641 & P1_R2358_U403); 
assign P1_R2358_U243 = ~(P1_R2358_U218 & P1_R2358_U215); 
assign P1_R2358_U252 = ~(P1_R2358_U123 & P1_R2358_U251); 
assign P1_R2358_U263 = ~(P1_U2640 & P1_R2358_U479); 
assign P1_R2358_U264 = ~(P1_U2639 & P1_R2358_U484); 
assign P1_R2358_U274 = ~(P1_R2358_U490 & P1_R2358_U489 & P1_R2358_U49); 
assign P1_R2358_U276 = ~(P1_R2358_U492 & P1_R2358_U491 & P1_R2358_U48); 
assign P1_R2358_U277 = ~(P1_U2632 & P1_R2358_U495); 
assign P1_R2358_U308 = ~(P1_R2358_U250 & P1_R2358_U207); 
assign P1_R2358_U506 = ~(P1_U2352 & P1_R2358_U168); 
assign P1_R2358_U519 = ~(P1_U2352 & P1_R2358_U168); 
assign P1_R2099_U18 = ~(P1_R2099_U172 & P1_R2099_U52); 
assign P1_R2099_U314 = ~(P1_R2099_U249 & P1_R2099_U172); 
assign P1_R2337_U46 = ~(P1_R2337_U113 & P1_PHYADDRPOINTER_REG_22__SCAN_IN); 
assign P1_R2337_U158 = ~(P1_R2337_U113 & P1_R2337_U45); 
assign P1_R2096_U46 = ~(P1_R2096_U113 & P1_REIP_REG_22__SCAN_IN); 
assign P1_R2096_U158 = ~(P1_R2096_U113 & P1_R2096_U45); 
assign P1_ADD_405_U46 = ~(P1_ADD_405_U116 & P1_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P1_ADD_405_U144 = ~(P1_ADD_405_U116 & P1_ADD_405_U45); 
assign P1_ADD_515_U46 = ~(P1_ADD_515_U113 & P1_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P1_ADD_515_U142 = ~(P1_ADD_515_U113 & P1_ADD_515_U45); 
assign P3_U2813 = ~(P3_U6542 & P3_U6541 & P3_U6543 & P3_U6544 & P3_U3971); 
assign P3_U2815 = ~(P3_U6526 & P3_U6525 & P3_U6528 & P3_U6527 & P3_U3969); 
assign P3_U3122 = ~(P3_U4629 & P3_STATE2_REG_0__SCAN_IN); 
assign P3_U3831 = P3_U3830 & P3_U3829 & P3_U6083; 
assign P3_U3838 = P3_U6116 & P3_U6115; 
assign P3_U3840 = P3_U6118 & P3_U6117 & P3_U6119 & P3_U3839; 
assign P3_U3843 = P3_U6130 & P3_U6129 & P3_U6128 & P3_U6127; 
assign P3_U3847 = P3_U6145 & P3_U6144; 
assign P3_U3850 = P3_U6147 & P3_U6146 & P3_U6148 & P3_U6150 & P3_U6149; 
assign P3_U3972 = P3_U6556 & P3_U6553 & P3_U6554 & P3_U6555; 
assign P3_U4102 = P3_U7278 & P3_U7277; 
assign P3_U4633 = ~(P3_U4629 & P3_U4338); 
assign P3_U4636 = ~(P3_U2390 & P3_U4629); 
assign P3_U4638 = ~(P3_U4629 & P3_U4337); 
assign P3_U5990 = ~(P3_U4318 & P3_U5988); 
assign P3_U6012 = ~(P3_U3810 & P3_U3807); 
assign P3_U6038 = ~(P3_U4318 & P3_U6036); 
assign P3_U6060 = ~(P3_U6042 & P3_U3819 & P3_U6040 & P3_U3824 & P3_U3820); 
assign P3_U6089 = ~(P3_SUB_357_1258_U86 & P3_U2393); 
assign P3_U6107 = ~(P3_ADD_371_1212_U10 & P3_U2360); 
assign P3_U6112 = ~(P3_ADD_360_1242_U10 & P3_U2395); 
assign P3_U6161 = ~(P3_SUB_357_1258_U84 & P3_U2393); 
assign P3_U6185 = ~(P3_SUB_357_1258_U83 & P3_U2393); 
assign P3_U6209 = ~(P3_SUB_357_1258_U82 & P3_U2393); 
assign P3_U6233 = ~(P3_SUB_357_1258_U81 & P3_U2393); 
assign P3_U6560 = ~(P3_U2394 & P3_SUB_357_1258_U86); 
assign P3_U6563 = ~(P3_U2387 & P3_ADD_371_1212_U10); 
assign P3_U6567 = ~(P3_U2396 & P3_ADD_360_1242_U10); 
assign P3_U6584 = ~(P3_U2394 & P3_SUB_357_1258_U84); 
assign P3_U6592 = ~(P3_U2394 & P3_SUB_357_1258_U83); 
assign P3_U6600 = ~(P3_U2394 & P3_SUB_357_1258_U82); 
assign P3_U6608 = ~(P3_U2394 & P3_SUB_357_1258_U81); 
assign P3_U7959 = ~(P3_U4637 & P3_U4629 & P3_U3121); 
assign P2_U2806 = P2_U3242 & P2_R2267_U8; 
assign P2_U2878 = ~(P2_U6499 & P2_U6500 & P2_U6498); 
assign P2_U3668 = ~(P2_U8392 & P2_U8391); 
assign P2_U3723 = P2_U4670 & P2_U4669 & P2_U4671; 
assign P2_U3724 = P2_U4675 & P2_U4674 & P2_U4676; 
assign P2_U3725 = P2_U4680 & P2_U4679 & P2_U4681; 
assign P2_U3726 = P2_U4685 & P2_U4684 & P2_U4686; 
assign P2_U3727 = P2_U4690 & P2_U4689 & P2_U4691; 
assign P2_U3728 = P2_U4695 & P2_U4694 & P2_U4696; 
assign P2_U3729 = P2_U4700 & P2_U4699 & P2_U4701; 
assign P2_U3730 = P2_U4705 & P2_U4704 & P2_U4706; 
assign P2_U3732 = P2_U4728 & P2_U4727 & P2_U4729; 
assign P2_U3733 = P2_U4733 & P2_U4732 & P2_U4734; 
assign P2_U3734 = P2_U4738 & P2_U4737 & P2_U4739; 
assign P2_U3735 = P2_U4743 & P2_U4742 & P2_U4744; 
assign P2_U3736 = P2_U4748 & P2_U4747 & P2_U4749; 
assign P2_U3737 = P2_U4753 & P2_U4752 & P2_U4754; 
assign P2_U3738 = P2_U4758 & P2_U4757 & P2_U4759; 
assign P2_U3739 = P2_U4763 & P2_U4762 & P2_U4764; 
assign P2_U3741 = P2_U4787 & P2_U4786 & P2_U4788; 
assign P2_U3742 = P2_U4792 & P2_U4791 & P2_U4793; 
assign P2_U3743 = P2_U4797 & P2_U4796 & P2_U4798; 
assign P2_U3744 = P2_U4802 & P2_U4801 & P2_U4803; 
assign P2_U3745 = P2_U4807 & P2_U4806 & P2_U4808; 
assign P2_U3746 = P2_U4812 & P2_U4811 & P2_U4813; 
assign P2_U3747 = P2_U4817 & P2_U4816 & P2_U4818; 
assign P2_U3748 = P2_U4822 & P2_U4821 & P2_U4823; 
assign P2_U3750 = P2_U4844 & P2_U4843 & P2_U4845; 
assign P2_U3751 = P2_U4849 & P2_U4848 & P2_U4850; 
assign P2_U3752 = P2_U4854 & P2_U4853 & P2_U4855; 
assign P2_U3753 = P2_U4859 & P2_U4858 & P2_U4860; 
assign P2_U3754 = P2_U4864 & P2_U4863 & P2_U4865; 
assign P2_U3755 = P2_U4869 & P2_U4868 & P2_U4870; 
assign P2_U3756 = P2_U4874 & P2_U4873 & P2_U4875; 
assign P2_U3757 = P2_U4879 & P2_U4878 & P2_U4880; 
assign P2_U3759 = P2_U4902 & P2_U4901 & P2_U4903; 
assign P2_U3760 = P2_U4907 & P2_U4906 & P2_U4908; 
assign P2_U3761 = P2_U4912 & P2_U4911 & P2_U4913; 
assign P2_U3762 = P2_U4917 & P2_U4916 & P2_U4918; 
assign P2_U3763 = P2_U4922 & P2_U4921 & P2_U4923; 
assign P2_U3764 = P2_U4927 & P2_U4926 & P2_U4928; 
assign P2_U3765 = P2_U4932 & P2_U4931 & P2_U4933; 
assign P2_U3766 = P2_U4937 & P2_U4936 & P2_U4938; 
assign P2_U3768 = P2_U4959 & P2_U4958 & P2_U4960; 
assign P2_U3769 = P2_U4964 & P2_U4963 & P2_U4965; 
assign P2_U3770 = P2_U4969 & P2_U4968 & P2_U4970; 
assign P2_U3771 = P2_U4974 & P2_U4973 & P2_U4975; 
assign P2_U3772 = P2_U4979 & P2_U4978 & P2_U4980; 
assign P2_U3773 = P2_U4984 & P2_U4983 & P2_U4985; 
assign P2_U3774 = P2_U4989 & P2_U4988 & P2_U4990; 
assign P2_U3775 = P2_U4994 & P2_U4993 & P2_U4995; 
assign P2_U3777 = P2_U5017 & P2_U5016 & P2_U5018; 
assign P2_U3778 = P2_U5022 & P2_U5021 & P2_U5023; 
assign P2_U3779 = P2_U5027 & P2_U5026 & P2_U5028; 
assign P2_U3780 = P2_U5032 & P2_U5031 & P2_U5033; 
assign P2_U3781 = P2_U5037 & P2_U5036 & P2_U5038; 
assign P2_U3782 = P2_U5042 & P2_U5041 & P2_U5043; 
assign P2_U3783 = P2_U5047 & P2_U5046 & P2_U5048; 
assign P2_U3784 = P2_U5052 & P2_U5051 & P2_U5053; 
assign P2_U3786 = P2_U5074 & P2_U5073 & P2_U5075; 
assign P2_U3787 = P2_U5079 & P2_U5078 & P2_U5080; 
assign P2_U3788 = P2_U5084 & P2_U5083 & P2_U5085; 
assign P2_U3789 = P2_U5089 & P2_U5088 & P2_U5090; 
assign P2_U3790 = P2_U5094 & P2_U5093 & P2_U5095; 
assign P2_U3791 = P2_U5099 & P2_U5098 & P2_U5100; 
assign P2_U3792 = P2_U5104 & P2_U5103 & P2_U5105; 
assign P2_U3793 = P2_U5109 & P2_U5108 & P2_U5110; 
assign P2_U4070 = P2_U6574 & P2_U6573 & P2_U4071; 
assign P2_U4074 = P2_U6583 & P2_U6582 & P2_U4075; 
assign P2_U4078 = P2_U6592 & P2_U6591 & P2_U4079; 
assign P2_U4082 = P2_U6601 & P2_U6600 & P2_U4083; 
assign P2_U4086 = P2_U6609 & P2_U4446 & P2_U6610; 
assign P2_U4090 = P2_U6618 & P2_U4446 & P2_U6619; 
assign P2_U4094 = P2_U6627 & P2_U4446 & P2_U6628; 
assign P2_U4097 = P2_U6635 & P2_U4446 & P2_U6636; 
assign P2_U4100 = P2_U6643 & P2_U4446 & P2_U6644; 
assign P2_U4103 = P2_U6651 & P2_U4446 & P2_U6652; 
assign P2_U4106 = P2_U6659 & P2_U4446 & P2_U6660; 
assign P2_U4109 = P2_U6667 & P2_U4446 & P2_U6668; 
assign P2_U4659 = ~(P2_U4445 & P2_U4658); 
assign P2_U4665 = ~(P2_U4445 & P2_U4664); 
assign P2_U4717 = ~(P2_U4445 & P2_U4716); 
assign P2_U4723 = ~(P2_U4445 & P2_U4722); 
assign P2_U4776 = ~(P2_U4445 & P2_U4775); 
assign P2_U4782 = ~(P2_U4445 & P2_U4781); 
assign P2_U4833 = ~(P2_U4445 & P2_U4832); 
assign P2_U4839 = ~(P2_U4445 & P2_U4838); 
assign P2_U4891 = ~(P2_U4445 & P2_U4890); 
assign P2_U4897 = ~(P2_U4445 & P2_U4896); 
assign P2_U4948 = ~(P2_U4445 & P2_U4947); 
assign P2_U4954 = ~(P2_U4445 & P2_U4953); 
assign P2_U5006 = ~(P2_U4445 & P2_U5005); 
assign P2_U5012 = ~(P2_U4445 & P2_U5011); 
assign P2_U5063 = ~(P2_U4445 & P2_U5062); 
assign P2_U5069 = ~(P2_U4445 & P2_U5068); 
assign P2_U5118 = ~(P2_U2493 & P2_U2362); 
assign P2_U5124 = ~(P2_U2493 & P2_U2398); 
assign P2_U5131 = ~(P2_U5113 & P2_U2421); 
assign P2_U5136 = ~(P2_U5113 & P2_U2419); 
assign P2_U5141 = ~(P2_U5113 & P2_U2417); 
assign P2_U5146 = ~(P2_U5113 & P2_U2415); 
assign P2_U5151 = ~(P2_U5113 & P2_U2413); 
assign P2_U5156 = ~(P2_U5113 & P2_U2411); 
assign P2_U5161 = ~(P2_U5113 & P2_U2409); 
assign P2_U5166 = ~(P2_U5113 & P2_U2407); 
assign P2_U5175 = ~(P2_U2495 & P2_U2362); 
assign P2_U5181 = ~(P2_U2495 & P2_U2398); 
assign P2_U5188 = ~(P2_U5169 & P2_U2421); 
assign P2_U5193 = ~(P2_U5169 & P2_U2419); 
assign P2_U5198 = ~(P2_U5169 & P2_U2417); 
assign P2_U5203 = ~(P2_U5169 & P2_U2415); 
assign P2_U5208 = ~(P2_U5169 & P2_U2413); 
assign P2_U5213 = ~(P2_U5169 & P2_U2411); 
assign P2_U5218 = ~(P2_U5169 & P2_U2409); 
assign P2_U5223 = ~(P2_U5169 & P2_U2407); 
assign P2_U5233 = ~(P2_U2497 & P2_U2362); 
assign P2_U5239 = ~(P2_U2497 & P2_U2398); 
assign P2_U5246 = ~(P2_U5226 & P2_U2421); 
assign P2_U5251 = ~(P2_U5226 & P2_U2419); 
assign P2_U5256 = ~(P2_U5226 & P2_U2417); 
assign P2_U5261 = ~(P2_U5226 & P2_U2415); 
assign P2_U5266 = ~(P2_U5226 & P2_U2413); 
assign P2_U5271 = ~(P2_U5226 & P2_U2411); 
assign P2_U5276 = ~(P2_U5226 & P2_U2409); 
assign P2_U5281 = ~(P2_U5226 & P2_U2407); 
assign P2_U5290 = ~(P2_U2499 & P2_U2362); 
assign P2_U5296 = ~(P2_U2499 & P2_U2398); 
assign P2_U5303 = ~(P2_U5284 & P2_U2421); 
assign P2_U5308 = ~(P2_U5284 & P2_U2419); 
assign P2_U5313 = ~(P2_U5284 & P2_U2417); 
assign P2_U5318 = ~(P2_U5284 & P2_U2415); 
assign P2_U5323 = ~(P2_U5284 & P2_U2413); 
assign P2_U5328 = ~(P2_U5284 & P2_U2411); 
assign P2_U5333 = ~(P2_U5284 & P2_U2409); 
assign P2_U5338 = ~(P2_U5284 & P2_U2407); 
assign P2_U5348 = ~(P2_U2505 & P2_U2362); 
assign P2_U5354 = ~(P2_U2505 & P2_U2398); 
assign P2_U5361 = ~(P2_U5341 & P2_U2421); 
assign P2_U5366 = ~(P2_U5341 & P2_U2419); 
assign P2_U5371 = ~(P2_U5341 & P2_U2417); 
assign P2_U5376 = ~(P2_U5341 & P2_U2415); 
assign P2_U5381 = ~(P2_U5341 & P2_U2413); 
assign P2_U5386 = ~(P2_U5341 & P2_U2411); 
assign P2_U5391 = ~(P2_U5341 & P2_U2409); 
assign P2_U5396 = ~(P2_U5341 & P2_U2407); 
assign P2_U5405 = ~(P2_U2507 & P2_U2362); 
assign P2_U5411 = ~(P2_U2507 & P2_U2398); 
assign P2_U5418 = ~(P2_U5399 & P2_U2421); 
assign P2_U5423 = ~(P2_U5399 & P2_U2419); 
assign P2_U5428 = ~(P2_U5399 & P2_U2417); 
assign P2_U5433 = ~(P2_U5399 & P2_U2415); 
assign P2_U5438 = ~(P2_U5399 & P2_U2413); 
assign P2_U5443 = ~(P2_U5399 & P2_U2411); 
assign P2_U5448 = ~(P2_U5399 & P2_U2409); 
assign P2_U5453 = ~(P2_U5399 & P2_U2407); 
assign P2_U5463 = ~(P2_U2509 & P2_U2362); 
assign P2_U5469 = ~(P2_U2509 & P2_U2398); 
assign P2_U5476 = ~(P2_U5456 & P2_U2421); 
assign P2_U5481 = ~(P2_U5456 & P2_U2419); 
assign P2_U5486 = ~(P2_U5456 & P2_U2417); 
assign P2_U5491 = ~(P2_U5456 & P2_U2415); 
assign P2_U5496 = ~(P2_U5456 & P2_U2413); 
assign P2_U5501 = ~(P2_U5456 & P2_U2411); 
assign P2_U5506 = ~(P2_U5456 & P2_U2409); 
assign P2_U5511 = ~(P2_U5456 & P2_U2407); 
assign P2_U5520 = ~(P2_U2511 & P2_U2362); 
assign P2_U5526 = ~(P2_U2511 & P2_U2398); 
assign P2_U5533 = ~(P2_U5514 & P2_U2421); 
assign P2_U5538 = ~(P2_U5514 & P2_U2419); 
assign P2_U5543 = ~(P2_U5514 & P2_U2417); 
assign P2_U5548 = ~(P2_U5514 & P2_U2415); 
assign P2_U5553 = ~(P2_U5514 & P2_U2413); 
assign P2_U5558 = ~(P2_U5514 & P2_U2411); 
assign P2_U5563 = ~(P2_U5514 & P2_U2409); 
assign P2_U5568 = ~(P2_U5514 & P2_U2407); 
assign P2_U5648 = ~(P2_U2398 & P2_U5647); 
assign P2_U6399 = ~(P2_U2380 & P2_R2096_U90); 
assign P2_U6501 = ~(P2_R2182_U96 & P2_U2393); 
assign P2_U6505 = ~(P2_U2379 & P2_R2099_U92); 
assign P2_U6575 = ~(P2_U7743 & P2_EBX_REG_0__SCAN_IN); 
assign P2_U6584 = ~(P2_U7743 & P2_EBX_REG_1__SCAN_IN); 
assign P2_U6593 = ~(P2_U7743 & P2_EBX_REG_2__SCAN_IN); 
assign P2_U6602 = ~(P2_U7743 & P2_EBX_REG_3__SCAN_IN); 
assign P2_U6611 = ~(P2_U7743 & P2_EBX_REG_4__SCAN_IN); 
assign P2_U6620 = ~(P2_U7743 & P2_EBX_REG_5__SCAN_IN); 
assign P2_U6629 = ~(P2_U7743 & P2_EBX_REG_6__SCAN_IN); 
assign P2_U6637 = ~(P2_U7743 & P2_EBX_REG_7__SCAN_IN); 
assign P2_U6645 = ~(P2_U7743 & P2_EBX_REG_8__SCAN_IN); 
assign P2_U6653 = ~(P2_U7743 & P2_EBX_REG_9__SCAN_IN); 
assign P2_U6661 = ~(P2_U7743 & P2_EBX_REG_10__SCAN_IN); 
assign P2_U6669 = ~(P2_U7743 & P2_EBX_REG_11__SCAN_IN); 
assign P2_U6670 = ~(P2_U2392 & P2_R2099_U92); 
assign P2_U6677 = ~(P2_U7743 & P2_EBX_REG_12__SCAN_IN); 
assign P2_U6685 = ~(P2_U7743 & P2_EBX_REG_13__SCAN_IN); 
assign P2_U6693 = ~(P2_U7743 & P2_EBX_REG_14__SCAN_IN); 
assign P2_U6699 = ~(P2_R2267_U8 & P2_U2587); 
assign P2_U6701 = ~(P2_U7743 & P2_EBX_REG_15__SCAN_IN); 
assign P2_U6709 = ~(P2_U7743 & P2_EBX_REG_16__SCAN_IN); 
assign P2_U6716 = ~(P2_U2588 & P2_R2096_U90); 
assign P2_U6717 = ~(P2_U7743 & P2_EBX_REG_17__SCAN_IN); 
assign P2_U6725 = ~(P2_U7743 & P2_EBX_REG_18__SCAN_IN); 
assign P2_U6733 = ~(P2_U7743 & P2_EBX_REG_19__SCAN_IN); 
assign P2_U6741 = ~(P2_U7743 & P2_EBX_REG_20__SCAN_IN); 
assign P2_U6749 = ~(P2_U7743 & P2_EBX_REG_21__SCAN_IN); 
assign P2_U6757 = ~(P2_U7743 & P2_EBX_REG_22__SCAN_IN); 
assign P2_U6765 = ~(P2_U7743 & P2_EBX_REG_23__SCAN_IN); 
assign P2_U6773 = ~(P2_U7743 & P2_EBX_REG_24__SCAN_IN); 
assign P2_U6781 = ~(P2_U7743 & P2_EBX_REG_25__SCAN_IN); 
assign P2_U6789 = ~(P2_U7743 & P2_EBX_REG_26__SCAN_IN); 
assign P2_U6797 = ~(P2_U7743 & P2_EBX_REG_27__SCAN_IN); 
assign P2_U6805 = ~(P2_U7743 & P2_EBX_REG_28__SCAN_IN); 
assign P2_U6813 = ~(P2_U7743 & P2_EBX_REG_29__SCAN_IN); 
assign P2_U6821 = ~(P2_U7743 & P2_EBX_REG_30__SCAN_IN); 
assign P2_U6829 = ~(P2_U7743 & P2_EBX_REG_31__SCAN_IN); 
assign P2_U8327 = ~(P2_R2256_U4 & P2_U3572); 
assign P1_U2480 = P1_U3315 & P1_U4548; 
assign P1_U2482 = P1_U3327 & P1_U4606; 
assign P1_U2484 = P1_U3334 & P1_U4665; 
assign P1_U2489 = P1_U3338 & P1_U4722; 
assign P1_U2492 = P1_U3343 & P1_U4780; 
assign P1_U2494 = P1_U3347 & P1_U4837; 
assign P1_U2496 = P1_U3350 & P1_U4895; 
assign P1_U2498 = P1_U3354 & P1_U4952; 
assign P1_U2636 = P1_R2144_U38 & P1_U6746; 
assign P1_U2637 = P1_R2144_U39 & P1_U6746; 
assign P1_U2786 = P1_U4159 & P1_R2144_U38; 
assign P1_U2787 = P1_U4159 & P1_R2144_U39; 
assign P1_U3030 = ~(P1_U3768 & P1_U3767 & P1_U3770); 
assign P1_U3359 = ~(P1_U2499 & P1_U4527); 
assign P1_U3364 = ~(P1_U2499 & P1_U4600); 
assign P1_U3367 = ~(P1_U2499 & P1_U4658); 
assign P1_U3371 = ~(P1_U2499 & P1_U2485); 
assign P1_U3374 = ~(P1_U2507 & P1_U4527); 
assign P1_U3378 = ~(P1_U2507 & P1_U4600); 
assign P1_U3381 = ~(P1_U2507 & P1_U4658); 
assign P1_U3385 = ~(P1_U2507 & P1_U2485); 
assign P1_U3477 = ~(P1_U7737 & P1_U7736); 
assign P1_U3478 = ~(P1_U7739 & P1_U7738); 
assign P1_U3829 = P1_U5718 & P1_U5720; 
assign P1_U3831 = P1_U3830 & P1_U5721; 
assign P1_U3928 = P1_U6524 & P1_U6522; 
assign P1_U4019 = P1_U6813 & P1_U6814 & P1_U6815; 
assign P1_U4532 = ~P1_U3315; 
assign P1_U4601 = ~P1_U3327; 
assign P1_U4659 = ~P1_U3334; 
assign P1_U4717 = ~P1_U3338; 
assign P1_U4774 = ~P1_U3343; 
assign P1_U4832 = ~P1_U3347; 
assign P1_U4889 = ~P1_U3350; 
assign P1_U4947 = ~P1_U3354; 
assign P1_U5549 = ~(P1_U3752 & P1_U5546); 
assign P1_U5586 = ~(P1_R2278_U107 & P1_U2377); 
assign P1_U5810 = ~(P1_U2372 & P1_R2278_U107); 
assign P1_U7604 = ~(P1_U7684 & P1_U7683 & P1_U3581); 
assign P3_ADD_476_U79 = ~(P3_ADD_476_U158 & P3_ADD_476_U157); 
assign P3_ADD_476_U114 = ~P3_ADD_476_U46; 
assign P3_ADD_476_U155 = ~(P3_ADD_476_U46 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_531_U83 = ~(P3_ADD_531_U165 & P3_ADD_531_U164); 
assign P3_ADD_531_U118 = ~P3_ADD_531_U47; 
assign P3_ADD_531_U162 = ~(P3_ADD_531_U47 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_SUB_320_U113 = ~(P3_SUB_320_U98 & P3_SUB_320_U69); 
assign P3_SUB_320_U147 = ~(P3_SUB_320_U98 & P3_SUB_320_U69); 
assign P3_ADD_318_U79 = ~(P3_ADD_318_U158 & P3_ADD_318_U157); 
assign P3_ADD_318_U114 = ~P3_ADD_318_U46; 
assign P3_ADD_318_U155 = ~(P3_ADD_318_U46 & P3_PHYADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_315_U75 = ~(P3_ADD_315_U150 & P3_ADD_315_U149); 
assign P3_ADD_315_U111 = ~P3_ADD_315_U46; 
assign P3_ADD_315_U147 = ~(P3_ADD_315_U46 & P3_PHYADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_360_1242_U60 = ~(P3_ADD_360_1242_U159 & P3_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P3_ADD_467_U79 = ~(P3_ADD_467_U158 & P3_ADD_467_U157); 
assign P3_ADD_467_U114 = ~P3_ADD_467_U46; 
assign P3_ADD_467_U155 = ~(P3_ADD_467_U46 & P3_REIP_REG_23__SCAN_IN); 
assign P3_ADD_430_U79 = ~(P3_ADD_430_U158 & P3_ADD_430_U157); 
assign P3_ADD_430_U114 = ~P3_ADD_430_U46; 
assign P3_ADD_430_U155 = ~(P3_ADD_430_U46 & P3_REIP_REG_23__SCAN_IN); 
assign P3_ADD_380_U83 = ~(P3_ADD_380_U165 & P3_ADD_380_U164); 
assign P3_ADD_380_U118 = ~P3_ADD_380_U47; 
assign P3_ADD_380_U162 = ~(P3_ADD_380_U47 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_344_U83 = ~(P3_ADD_344_U165 & P3_ADD_344_U164); 
assign P3_ADD_344_U118 = ~P3_ADD_344_U47; 
assign P3_ADD_344_U162 = ~(P3_ADD_344_U47 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_339_U79 = ~(P3_ADD_339_U158 & P3_ADD_339_U157); 
assign P3_ADD_339_U114 = ~P3_ADD_339_U46; 
assign P3_ADD_339_U155 = ~(P3_ADD_339_U46 & P3_PHYADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_541_U79 = ~(P3_ADD_541_U158 & P3_ADD_541_U157); 
assign P3_ADD_541_U114 = ~P3_ADD_541_U46; 
assign P3_ADD_541_U155 = ~(P3_ADD_541_U46 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_SUB_357_1258_U18 = P3_SUB_357_1258_U233 & P3_SUB_357_1258_U230; 
assign P3_SUB_357_1258_U129 = ~(P3_SUB_357_1258_U275 & P3_SUB_357_1258_U274 & P3_SUB_357_1258_U304); 
assign P3_SUB_357_1258_U139 = ~(P3_SUB_357_1258_U111 & P3_SUB_357_1258_U236); 
assign P3_SUB_357_1258_U226 = ~(P3_SUB_357_1258_U221 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_SUB_357_1258_U239 = ~(P3_SUB_357_1258_U235 & P3_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P3_SUB_357_1258_U377 = ~(P3_SUB_357_1258_U306 & P3_SUB_357_1258_U39); 
assign P3_SUB_357_1258_U384 = ~(P3_SUB_357_1258_U220 & P3_SUB_357_1258_U382); 
assign P3_ADD_515_U79 = ~(P3_ADD_515_U158 & P3_ADD_515_U157); 
assign P3_ADD_515_U114 = ~P3_ADD_515_U46; 
assign P3_ADD_515_U155 = ~(P3_ADD_515_U46 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_394_U78 = ~(P3_ADD_394_U160 & P3_ADD_394_U159); 
assign P3_ADD_394_U117 = ~P3_ADD_394_U46; 
assign P3_ADD_394_U157 = ~(P3_ADD_394_U46 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_441_U79 = ~(P3_ADD_441_U158 & P3_ADD_441_U157); 
assign P3_ADD_441_U114 = ~P3_ADD_441_U46; 
assign P3_ADD_441_U155 = ~(P3_ADD_441_U46 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_349_U83 = ~(P3_ADD_349_U165 & P3_ADD_349_U164); 
assign P3_ADD_349_U118 = ~P3_ADD_349_U47; 
assign P3_ADD_349_U162 = ~(P3_ADD_349_U47 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_405_U78 = ~(P3_ADD_405_U160 & P3_ADD_405_U159); 
assign P3_ADD_405_U117 = ~P3_ADD_405_U46; 
assign P3_ADD_405_U157 = ~(P3_ADD_405_U46 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_553_U83 = ~(P3_ADD_553_U165 & P3_ADD_553_U164); 
assign P3_ADD_553_U118 = ~P3_ADD_553_U47; 
assign P3_ADD_553_U162 = ~(P3_ADD_553_U47 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_558_U83 = ~(P3_ADD_558_U165 & P3_ADD_558_U164); 
assign P3_ADD_558_U118 = ~P3_ADD_558_U47; 
assign P3_ADD_558_U162 = ~(P3_ADD_558_U47 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_385_U83 = ~(P3_ADD_385_U165 & P3_ADD_385_U164); 
assign P3_ADD_385_U118 = ~P3_ADD_385_U47; 
assign P3_ADD_385_U162 = ~(P3_ADD_385_U47 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_547_U83 = ~(P3_ADD_547_U165 & P3_ADD_547_U164); 
assign P3_ADD_547_U118 = ~P3_ADD_547_U47; 
assign P3_ADD_547_U162 = ~(P3_ADD_547_U47 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_371_1212_U11 = P3_ADD_371_1212_U185 & P3_ADD_371_1212_U168; 
assign P3_ADD_371_1212_U169 = ~P3_ADD_371_1212_U62; 
assign P3_ADD_371_1212_U184 = ~(P3_ADD_371_1212_U61 & P3_ADD_371_1212_U168); 
assign P3_ADD_371_1212_U249 = ~(P3_ADD_371_1212_U62 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_494_U79 = ~(P3_ADD_494_U158 & P3_ADD_494_U157); 
assign P3_ADD_494_U114 = ~P3_ADD_494_U46; 
assign P3_ADD_494_U155 = ~(P3_ADD_494_U46 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_536_U79 = ~(P3_ADD_536_U158 & P3_ADD_536_U157); 
assign P3_ADD_536_U114 = ~P3_ADD_536_U46; 
assign P3_ADD_536_U155 = ~(P3_ADD_536_U46 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P2_R2099_U31 = ~(P2_U2735 & P2_R2099_U127); 
assign P2_R2099_U219 = ~(P2_R2099_U127 & P2_R2099_U30); 
assign P2_ADD_391_1196_U9 = P2_ADD_391_1196_U205 & P2_ADD_391_1196_U203; 
assign P2_ADD_391_1196_U48 = ~P2_R2182_U96; 
assign P2_ADD_391_1196_U57 = ~P2_R2096_U90; 
assign P2_ADD_391_1196_U111 = P2_ADD_391_1196_U310 & P2_ADD_391_1196_U309; 
assign P2_ADD_391_1196_U158 = ~(P2_R2096_U97 & P2_R2182_U96); 
assign P2_ADD_391_1196_U182 = ~(P2_ADD_391_1196_U181 & P2_ADD_391_1196_U161); 
assign P2_ADD_391_1196_U199 = ~(P2_ADD_391_1196_U198 & P2_ADD_391_1196_U161 & P2_ADD_391_1196_U113); 
assign P2_ADD_391_1196_U210 = P2_R2096_U97 | P2_R2182_U96; 
assign P2_ADD_391_1196_U297 = P2_R2182_U96 | P2_R2096_U97; 
assign P2_ADD_391_1196_U302 = P2_R2096_U97 | P2_R2182_U96; 
assign P2_ADD_391_1196_U307 = ~(P2_R2096_U69 & P2_ADD_391_1196_U34); 
assign P2_ADD_391_1196_U313 = ~(P2_ADD_391_1196_U312 & P2_ADD_391_1196_U311); 
assign P2_ADD_391_1196_U322 = ~(P2_ADD_391_1196_U320 & P2_ADD_391_1196_U181); 
assign P2_ADD_391_1196_U473 = ~(P2_R2182_U96 & P2_ADD_391_1196_U49); 
assign P2_R2182_U14 = P2_U2668 & P2_R2182_U6; 
assign P2_R2182_U95 = ~(P2_R2182_U301 & P2_R2182_U300); 
assign P2_R2182_U144 = ~P2_R2182_U6; 
assign P2_R2182_U296 = ~(P2_R2182_U38 & P2_R2182_U6); 
assign P2_R2182_U299 = ~(P2_R2182_U143 & P2_U2669); 
assign P2_R2027_U83 = ~(P2_R2027_U165 & P2_R2027_U164); 
assign P2_R2027_U118 = ~P2_R2027_U47; 
assign P2_R2027_U162 = ~(P2_R2027_U47 & P2_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P2_LT_563_1260_U6 = P2_LT_563_1260_U7 | P2_U3617; 
assign P2_R2337_U77 = ~(P2_R2337_U156 & P2_R2337_U155); 
assign P2_R2337_U115 = ~P2_R2337_U47; 
assign P2_R2337_U153 = ~(P2_R2337_U47 & P2_PHYADDRPOINTER_REG_24__SCAN_IN); 
assign P2_R2096_U7 = P2_U2629 & P2_R2096_U16; 
assign P2_R2096_U89 = ~(P2_R2096_U247 & P2_R2096_U246); 
assign P2_R2096_U155 = ~P2_R2096_U16; 
assign P2_R2096_U237 = ~(P2_R2096_U36 & P2_R2096_U16); 
assign P2_R2096_U245 = ~(P2_R2096_U154 & P2_U2630); 
assign P2_LT_563_U20 = ~(P2_LT_563_U18 & P2_LT_563_U19 & P2_LT_563_U17); 
assign P2_R2256_U10 = ~(P2_U3626 & P2_R2256_U25); 
assign P2_R2256_U22 = ~(P2_R2256_U63 & P2_R2256_U62); 
assign P2_R2256_U40 = ~P2_R2256_U25; 
assign P2_R2256_U55 = ~(P2_U3626 & P2_R2256_U25); 
assign P2_R1957_U113 = ~(P2_R1957_U98 & P2_R1957_U69); 
assign P2_R1957_U147 = ~(P2_R1957_U98 & P2_R1957_U69); 
assign P2_R2278_U56 = ~P2_U2807; 
assign P2_R2278_U58 = ~(P2_U2807 & P2_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P2_R2278_U123 = P2_R2278_U245 & P2_R2278_U249; 
assign P2_R2278_U199 = P2_R2278_U541 & P2_R2278_U540; 
assign P2_R2278_U208 = ~P2_R2278_U15; 
assign P2_R2278_U252 = P2_U2807 | P2_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P2_R2278_U324 = ~(P2_R2278_U247 & P2_R2278_U249); 
assign P2_R2278_U486 = ~(P2_R2278_U15 & P2_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P2_R2278_U527 = ~(P2_U2807 & P2_R2278_U57); 
assign P2_R2278_U529 = ~(P2_U2807 & P2_R2278_U57); 
assign P2_R2278_U533 = ~(P2_R2278_U45 & P2_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P2_R2278_U535 = ~(P2_R2278_U45 & P2_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P2_R2278_U544 = ~(P2_R2278_U543 & P2_R2278_U542); 
assign P2_R2278_U561 = ~(P2_R2278_U13 & P2_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P2_ADD_394_U71 = ~(P2_ADD_394_U144 & P2_ADD_394_U143); 
assign P2_ADD_394_U117 = ~P2_ADD_394_U46; 
assign P2_ADD_394_U163 = ~(P2_ADD_394_U46 & P2_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P2_R2267_U81 = P2_R2267_U160 & P2_R2267_U159; 
assign P2_R2267_U105 = ~P2_R2267_U34; 
assign P2_R2267_U127 = ~(P2_U2780 & P2_R2267_U126); 
assign P2_R2267_U157 = ~(P2_U2779 & P2_R2267_U34); 
assign P2_ADD_371_1212_U30 = ~P2_R2256_U4; 
assign P2_ADD_371_1212_U67 = ~(P2_R2256_U4 & P2_ADD_371_1212_U137); 
assign P2_ADD_371_1212_U267 = ~(P2_ADD_371_1212_U266 & P2_ADD_371_1212_U265); 
assign P2_ADD_371_1212_U268 = ~(P2_ADD_371_1212_U29 & P2_ADD_371_1212_U28 & P2_R2256_U4); 
assign P1_R2144_U247 = ~(P1_R2144_U147 & P1_R2144_U225); 
assign P1_R2278_U6 = P1_R2278_U292 & P1_R2278_U288; 
assign P1_R2278_U9 = P1_R2278_U8 & P1_R2278_U308; 
assign P1_R2278_U11 = P1_R2278_U134 & P1_R2278_U10; 
assign P1_R2278_U14 = P1_R2278_U463 & P1_R2278_U462; 
assign P1_R2278_U100 = P1_R2278_U262 & P1_R2278_U261; 
assign P1_R2278_U124 = P1_R2278_U68 & P1_R2278_U281; 
assign P1_R2278_U128 = P1_R2278_U258 & P1_R2278_U254; 
assign P1_R2278_U137 = P1_R2278_U259 & P1_R2278_U228 & P1_R2278_U273; 
assign P1_R2278_U143 = P1_R2278_U309 & P1_R2278_U321; 
assign P1_R2278_U144 = P1_R2278_U296 & P1_R2278_U308; 
assign P1_R2278_U164 = P1_R2278_U317 & P1_R2278_U10; 
assign P1_R2278_U167 = P1_R2278_U370 & P1_R2278_U314; 
assign P1_R2278_U172 = P1_R2278_U364 & P1_R2278_U303; 
assign P1_R2278_U182 = ~(P1_R2278_U242 & P1_R2278_U241); 
assign P1_R2278_U189 = P1_R2278_U472 & P1_R2278_U471; 
assign P1_R2278_U193 = P1_R2278_U486 & P1_R2278_U485; 
assign P1_R2278_U195 = P1_R2278_U493 & P1_R2278_U492; 
assign P1_R2278_U197 = P1_R2278_U500 & P1_R2278_U499; 
assign P1_R2278_U199 = P1_R2278_U507 & P1_R2278_U506; 
assign P1_R2278_U201 = P1_R2278_U514 & P1_R2278_U513; 
assign P1_R2278_U203 = P1_R2278_U521 & P1_R2278_U520; 
assign P1_R2278_U205 = P1_R2278_U528 & P1_R2278_U527; 
assign P1_R2278_U207 = P1_R2278_U535 & P1_R2278_U534; 
assign P1_R2278_U209 = P1_R2278_U542 & P1_R2278_U541; 
assign P1_R2278_U211 = P1_R2278_U549 & P1_R2278_U548; 
assign P1_R2278_U215 = P1_R2278_U561 & P1_R2278_U560; 
assign P1_R2278_U217 = P1_R2278_U568 & P1_R2278_U567; 
assign P1_R2278_U219 = P1_R2278_U575 & P1_R2278_U574; 
assign P1_R2278_U282 = ~P1_R2278_U68; 
assign P1_R2278_U346 = ~(P1_R2278_U263 & P1_R2278_U261); 
assign P1_R2278_U350 = ~(P1_R2278_U68 & P1_R2278_U281); 
assign P1_R2278_U351 = ~(P1_R2278_U345 & P1_R2278_U228); 
assign P1_R2278_U352 = ~(P1_R2278_U127 & P1_R2278_U258); 
assign P1_R2278_U359 = ~(P1_R2278_U293 & P1_R2278_U290); 
assign P1_R2278_U366 = ~(P1_R2278_U364 & P1_R2278_U303); 
assign P1_R2278_U379 = ~(P1_R2278_U320 & P1_R2278_U321); 
assign P1_R2278_U381 = ~(P1_R2278_U370 & P1_R2278_U314); 
assign P1_R2278_U388 = ~(P1_R2278_U277 & P1_R2278_U261); 
assign P1_R2278_U433 = ~(P1_R2278_U22 & P1_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P1_R2278_U435 = ~(P1_R2278_U22 & P1_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P1_R2278_U443 = ~(P1_R2278_U442 & P1_R2278_U441); 
assign P1_R2278_U461 = ~(P1_R2278_U239 & P1_R2278_U459); 
assign P1_R2278_U466 = ~(P1_R2278_U465 & P1_R2278_U464); 
assign P1_R2278_U475 = ~(P1_R2278_U474 & P1_R2278_U473); 
assign P1_R2278_U489 = ~(P1_R2278_U488 & P1_R2278_U487); 
assign P1_R2278_U496 = ~(P1_R2278_U495 & P1_R2278_U494); 
assign P1_R2278_U503 = ~(P1_R2278_U502 & P1_R2278_U501); 
assign P1_R2278_U510 = ~(P1_R2278_U509 & P1_R2278_U508); 
assign P1_R2278_U517 = ~(P1_R2278_U516 & P1_R2278_U515); 
assign P1_R2278_U524 = ~(P1_R2278_U523 & P1_R2278_U522); 
assign P1_R2278_U531 = ~(P1_R2278_U530 & P1_R2278_U529); 
assign P1_R2278_U538 = ~(P1_R2278_U537 & P1_R2278_U536); 
assign P1_R2278_U545 = ~(P1_R2278_U544 & P1_R2278_U543); 
assign P1_R2278_U552 = ~(P1_R2278_U551 & P1_R2278_U550); 
assign P1_R2278_U564 = ~(P1_R2278_U563 & P1_R2278_U562); 
assign P1_R2278_U571 = ~(P1_R2278_U570 & P1_R2278_U569); 
assign P1_R2278_U578 = ~(P1_R2278_U577 & P1_R2278_U576); 
assign P1_R2278_U582 = ~(P1_R2278_U70 & P1_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P1_R2278_U584 = ~(P1_R2278_U70 & P1_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P1_R2278_U603 = ~(P1_R2278_U59 & P1_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P1_R2278_U605 = ~(P1_R2278_U61 & P1_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P1_R2358_U18 = P1_R2358_U308 & P1_R2358_U307; 
assign P1_R2358_U19 = P1_R2358_U254 & P1_R2358_U252; 
assign P1_R2358_U54 = ~(P1_R2358_U400 & P1_R2358_U399 & P1_R2358_U34); 
assign P1_R2358_U79 = P1_R2358_U229 & P1_R2358_U228; 
assign P1_R2358_U110 = P1_R2358_U277 & P1_R2358_U276; 
assign P1_R2358_U112 = P1_R2358_U275 & P1_R2358_U274; 
assign P1_R2358_U169 = ~P1_U2662; 
assign P1_R2358_U214 = ~P1_R2358_U156; 
assign P1_R2358_U224 = ~(P1_R2358_U218 & P1_R2358_U223 & P1_R2358_U217); 
assign P1_R2358_U226 = ~(P1_R2358_U225 & P1_R2358_U156 & P1_R2358_U219 & P1_R2358_U218 & P1_R2358_U217); 
assign P1_R2358_U234 = ~(P1_R2358_U225 & P1_R2358_U156); 
assign P1_R2358_U259 = ~(P1_R2358_U486 & P1_R2358_U485 & P1_R2358_U56); 
assign P1_R2358_U262 = ~(P1_R2358_U476 & P1_R2358_U475 & P1_R2358_U53); 
assign P1_R2358_U265 = ~(P1_R2358_U12 & P1_R2358_U52); 
assign P1_R2358_U266 = ~(P1_R2358_U233 & P1_R2358_U228 & P1_R2358_U263); 
assign P1_R2358_U270 = ~P1_R2358_U57; 
assign P1_R2358_U272 = ~(P1_R2358_U488 & P1_R2358_U487 & P1_R2358_U50); 
assign P1_R2358_U273 = ~P1_R2358_U51; 
assign P1_R2358_U278 = ~(P1_R2358_U507 & P1_R2358_U506 & P1_R2358_U46); 
assign P1_R2358_U333 = ~(P1_R2358_U229 & P1_R2358_U228); 
assign P1_R2358_U348 = ~(P1_R2358_U277 & P1_R2358_U276); 
assign P1_R2358_U349 = ~(P1_R2358_U275 & P1_R2358_U274); 
assign P1_R2358_U360 = ~(P1_R2358_U12 & P1_R2358_U52); 
assign P1_R2358_U455 = ~(P1_R2358_U335 & P1_R2358_U156); 
assign P1_R2358_U509 = ~(P1_U2662 & P1_R2358_U23); 
assign P1_R2358_U517 = ~(P1_U2662 & P1_R2358_U23); 
assign P1_R2358_U521 = ~(P1_R2358_U520 & P1_R2358_U519); 
assign P1_R2099_U74 = ~(P1_R2099_U315 & P1_R2099_U314); 
assign P1_R2099_U173 = ~P1_R2099_U18; 
assign P1_R2099_U313 = ~(P1_R2099_U51 & P1_R2099_U18); 
assign P1_R2337_U79 = ~(P1_R2337_U158 & P1_R2337_U157); 
assign P1_R2337_U114 = ~P1_R2337_U46; 
assign P1_R2337_U155 = ~(P1_R2337_U46 & P1_PHYADDRPOINTER_REG_23__SCAN_IN); 
assign P1_R2096_U79 = ~(P1_R2096_U158 & P1_R2096_U157); 
assign P1_R2096_U114 = ~P1_R2096_U46; 
assign P1_R2096_U155 = ~(P1_R2096_U46 & P1_REIP_REG_23__SCAN_IN); 
assign P1_ADD_405_U71 = ~(P1_ADD_405_U144 & P1_ADD_405_U143); 
assign P1_ADD_405_U117 = ~P1_ADD_405_U46; 
assign P1_ADD_405_U163 = ~(P1_ADD_405_U46 & P1_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P1_ADD_515_U71 = ~(P1_ADD_515_U142 & P1_ADD_515_U141); 
assign P1_ADD_515_U114 = ~P1_ADD_515_U46; 
assign P1_ADD_515_U161 = ~(P1_ADD_515_U46 & P1_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_U2812 = ~(P3_U6550 & P3_U6549 & P3_U6551 & P3_U6552 & P3_U3972); 
assign P3_U2846 = ~(P3_U6039 & P3_U6037 & P3_U6038); 
assign P3_U2848 = ~(P3_U3803 & P3_U5990); 
assign P3_U3833 = P3_U6094 & P3_U6093 & P3_U6095 & P3_U3834 & P3_U6089; 
assign P3_U3837 = P3_U3836 & P3_U3835 & P3_U6107; 
assign P3_U3973 = P3_U6564 & P3_U6561 & P3_U6562 & P3_U6563; 
assign P3_U4630 = ~P3_U3122; 
assign P3_U4632 = ~(P3_U3122 & P3_STATE2_REG_2__SCAN_IN); 
assign P3_U4635 = ~(P3_U4633 & P3_STATE2_REG_1__SCAN_IN); 
assign P3_U6014 = ~(P3_U4318 & P3_U6012); 
assign P3_U6062 = ~(P3_U4318 & P3_U6060); 
assign P3_U6084 = ~(P3_U6066 & P3_U3828 & P3_U6064 & P3_U3825 & P3_U3831); 
assign P3_U6131 = ~(P3_ADD_371_1212_U11 & P3_U2360); 
assign P3_U6138 = ~(P3_ADD_558_U83 & P3_U3220); 
assign P3_U6139 = ~(P3_ADD_553_U83 & P3_U4298); 
assign P3_U6140 = ~(P3_ADD_547_U83 & P3_U4299); 
assign P3_U6143 = ~(P3_ADD_531_U83 & P3_U2354); 
assign P3_U6151 = ~(P3_ADD_385_U83 & P3_U2358); 
assign P3_U6152 = ~(P3_ADD_380_U83 & P3_U2359); 
assign P3_U6153 = ~(P3_ADD_349_U83 & P3_U4306); 
assign P3_U6154 = ~(P3_ADD_344_U83 & P3_U2362); 
assign P3_U6165 = ~(P3_ADD_541_U79 & P3_U4300); 
assign P3_U6166 = ~(P3_ADD_536_U79 & P3_U4301); 
assign P3_U6169 = ~(P3_ADD_515_U79 & P3_U4302); 
assign P3_U6170 = ~(P3_ADD_494_U79 & P3_U2356); 
assign P3_U6171 = ~(P3_ADD_476_U79 & P3_U4303); 
assign P3_U6172 = ~(P3_ADD_441_U79 & P3_U4304); 
assign P3_U6173 = ~(P3_ADD_405_U78 & P3_U4305); 
assign P3_U6174 = ~(P3_ADD_394_U78 & P3_U2357); 
assign P3_U6257 = ~(P3_SUB_357_1258_U18 & P3_U2393); 
assign P3_U6571 = ~(P3_U2387 & P3_ADD_371_1212_U11); 
assign P3_U6581 = ~(P3_ADD_318_U79 & P3_U2398); 
assign P3_U6586 = ~(P3_ADD_339_U79 & P3_U2388); 
assign P3_U6590 = ~(P3_ADD_315_U75 & P3_U2397); 
assign P3_U6616 = ~(P3_U2394 & P3_SUB_357_1258_U18); 
assign P3_U7286 = ~(P3_ADD_467_U79 & P3_U2601); 
assign P3_U7288 = ~(P3_ADD_430_U79 & P3_U2405); 
assign P3_U7954 = ~(P3_U3122 & P3_STATE2_REG_3__SCAN_IN); 
assign P3_U7958 = ~(P3_U4638 & P3_STATE2_REG_0__SCAN_IN); 
assign P2_U2805 = P2_U3242 & P2_R2267_U81; 
assign P2_U2877 = ~(P2_U6502 & P2_U6503 & P2_U6501); 
assign P2_U3637 = ~(P2_U8328 & P2_U8327); 
assign P2_U3795 = P2_U5130 & P2_U5129 & P2_U5131; 
assign P2_U3796 = P2_U5135 & P2_U5134 & P2_U5136; 
assign P2_U3797 = P2_U5140 & P2_U5139 & P2_U5141; 
assign P2_U3798 = P2_U5145 & P2_U5144 & P2_U5146; 
assign P2_U3799 = P2_U5150 & P2_U5149 & P2_U5151; 
assign P2_U3800 = P2_U5155 & P2_U5154 & P2_U5156; 
assign P2_U3801 = P2_U5160 & P2_U5159 & P2_U5161; 
assign P2_U3802 = P2_U5165 & P2_U5164 & P2_U5166; 
assign P2_U3804 = P2_U5187 & P2_U5186 & P2_U5188; 
assign P2_U3805 = P2_U5192 & P2_U5191 & P2_U5193; 
assign P2_U3806 = P2_U5197 & P2_U5196 & P2_U5198; 
assign P2_U3807 = P2_U5202 & P2_U5201 & P2_U5203; 
assign P2_U3808 = P2_U5207 & P2_U5206 & P2_U5208; 
assign P2_U3809 = P2_U5212 & P2_U5211 & P2_U5213; 
assign P2_U3810 = P2_U5217 & P2_U5216 & P2_U5218; 
assign P2_U3811 = P2_U5222 & P2_U5221 & P2_U5223; 
assign P2_U3813 = P2_U5245 & P2_U5244 & P2_U5246; 
assign P2_U3814 = P2_U5250 & P2_U5249 & P2_U5251; 
assign P2_U3815 = P2_U5255 & P2_U5254 & P2_U5256; 
assign P2_U3816 = P2_U5260 & P2_U5259 & P2_U5261; 
assign P2_U3817 = P2_U5265 & P2_U5264 & P2_U5266; 
assign P2_U3818 = P2_U5270 & P2_U5269 & P2_U5271; 
assign P2_U3819 = P2_U5275 & P2_U5274 & P2_U5276; 
assign P2_U3820 = P2_U5280 & P2_U5279 & P2_U5281; 
assign P2_U3822 = P2_U5302 & P2_U5301 & P2_U5303; 
assign P2_U3823 = P2_U5307 & P2_U5306 & P2_U5308; 
assign P2_U3824 = P2_U5312 & P2_U5311 & P2_U5313; 
assign P2_U3825 = P2_U5317 & P2_U5316 & P2_U5318; 
assign P2_U3826 = P2_U5322 & P2_U5321 & P2_U5323; 
assign P2_U3827 = P2_U5327 & P2_U5326 & P2_U5328; 
assign P2_U3828 = P2_U5332 & P2_U5331 & P2_U5333; 
assign P2_U3829 = P2_U5337 & P2_U5336 & P2_U5338; 
assign P2_U3831 = P2_U5360 & P2_U5359 & P2_U5361; 
assign P2_U3832 = P2_U5365 & P2_U5364 & P2_U5366; 
assign P2_U3833 = P2_U5370 & P2_U5369 & P2_U5371; 
assign P2_U3834 = P2_U5375 & P2_U5374 & P2_U5376; 
assign P2_U3835 = P2_U5380 & P2_U5379 & P2_U5381; 
assign P2_U3836 = P2_U5385 & P2_U5384 & P2_U5386; 
assign P2_U3837 = P2_U5390 & P2_U5389 & P2_U5391; 
assign P2_U3838 = P2_U5395 & P2_U5394 & P2_U5396; 
assign P2_U3840 = P2_U5417 & P2_U5416 & P2_U5418; 
assign P2_U3841 = P2_U5422 & P2_U5421 & P2_U5423; 
assign P2_U3842 = P2_U5427 & P2_U5426 & P2_U5428; 
assign P2_U3843 = P2_U5432 & P2_U5431 & P2_U5433; 
assign P2_U3844 = P2_U5437 & P2_U5436 & P2_U5438; 
assign P2_U3845 = P2_U5442 & P2_U5441 & P2_U5443; 
assign P2_U3846 = P2_U5447 & P2_U5446 & P2_U5448; 
assign P2_U3847 = P2_U5452 & P2_U5451 & P2_U5453; 
assign P2_U3849 = P2_U5475 & P2_U5474 & P2_U5476; 
assign P2_U3850 = P2_U5480 & P2_U5479 & P2_U5481; 
assign P2_U3851 = P2_U5485 & P2_U5484 & P2_U5486; 
assign P2_U3852 = P2_U5490 & P2_U5489 & P2_U5491; 
assign P2_U3853 = P2_U5495 & P2_U5494 & P2_U5496; 
assign P2_U3854 = P2_U5500 & P2_U5499 & P2_U5501; 
assign P2_U3855 = P2_U5505 & P2_U5504 & P2_U5506; 
assign P2_U3856 = P2_U5510 & P2_U5509 & P2_U5511; 
assign P2_U3858 = P2_U5532 & P2_U5531 & P2_U5533; 
assign P2_U3859 = P2_U5537 & P2_U5536 & P2_U5538; 
assign P2_U3860 = P2_U5542 & P2_U5541 & P2_U5543; 
assign P2_U3861 = P2_U5547 & P2_U5546 & P2_U5548; 
assign P2_U3862 = P2_U5552 & P2_U5551 & P2_U5553; 
assign P2_U3863 = P2_U5557 & P2_U5556 & P2_U5558; 
assign P2_U3864 = P2_U5562 & P2_U5561 & P2_U5563; 
assign P2_U3865 = P2_U5567 & P2_U5566 & P2_U5568; 
assign P2_U4121 = P2_U6699 & P2_U4446; 
assign P2_U4444 = ~P2_LT_563_1260_U6; 
assign P2_U4660 = ~(P2_U4652 & P2_U4659); 
assign P2_U4666 = ~(P2_U4665 & P2_U3325); 
assign P2_U4718 = ~(P2_U4717 & P2_U3245); 
assign P2_U4724 = ~(P2_U4723 & P2_U4712); 
assign P2_U4777 = ~(P2_U4771 & P2_U4776); 
assign P2_U4783 = ~(P2_U4782 & P2_U3355); 
assign P2_U4834 = ~(P2_U4833 & P2_U3246); 
assign P2_U4840 = ~(P2_U4839 & P2_U4828); 
assign P2_U4892 = ~(P2_U4886 & P2_U4891); 
assign P2_U4898 = ~(P2_U4897 & P2_U3380); 
assign P2_U4949 = ~(P2_U4948 & P2_U3247); 
assign P2_U4955 = ~(P2_U4954 & P2_U4943); 
assign P2_U5007 = ~(P2_U5001 & P2_U5006); 
assign P2_U5013 = ~(P2_U5012 & P2_U3403); 
assign P2_U5064 = ~(P2_U5063 & P2_U3248); 
assign P2_U5070 = ~(P2_U5069 & P2_U5058); 
assign P2_U5119 = ~(P2_U4445 & P2_U5118); 
assign P2_U5125 = ~(P2_U4445 & P2_U5124); 
assign P2_U5176 = ~(P2_U4445 & P2_U5175); 
assign P2_U5182 = ~(P2_U4445 & P2_U5181); 
assign P2_U5234 = ~(P2_U4445 & P2_U5233); 
assign P2_U5240 = ~(P2_U4445 & P2_U5239); 
assign P2_U5291 = ~(P2_U4445 & P2_U5290); 
assign P2_U5297 = ~(P2_U4445 & P2_U5296); 
assign P2_U5349 = ~(P2_U4445 & P2_U5348); 
assign P2_U5355 = ~(P2_U4445 & P2_U5354); 
assign P2_U5406 = ~(P2_U4445 & P2_U5405); 
assign P2_U5412 = ~(P2_U4445 & P2_U5411); 
assign P2_U5464 = ~(P2_U4445 & P2_U5463); 
assign P2_U5470 = ~(P2_U4445 & P2_U5469); 
assign P2_U5521 = ~(P2_U4445 & P2_U5520); 
assign P2_U5527 = ~(P2_U4445 & P2_U5526); 
assign P2_U5651 = ~(P2_U3891 & P2_U5648); 
assign P2_U6348 = ~(P2_ADD_391_1196_U9 & P2_U2397); 
assign P2_U6404 = ~(P2_U2380 & P2_R2096_U89); 
assign P2_U6504 = ~(P2_R2182_U95 & P2_U2393); 
assign P2_U6707 = ~(P2_R2267_U81 & P2_U2587); 
assign P2_U6724 = ~(P2_U2588 & P2_R2096_U89); 
assign P2_U8325 = ~(P2_R2256_U22 & P2_U3572); 
assign P2_U8389 = ~(P2_R2337_U77 & P2_U3284); 
assign P1_U2500 = P1_U3359 & P1_U3357; 
assign P1_U2502 = P1_U3364 & P1_U5065; 
assign P1_U2504 = P1_U3367 & P1_U5123; 
assign P1_U2506 = P1_U3371 & P1_U5180; 
assign P1_U2511 = P1_U3374 & P1_U5238; 
assign P1_U2513 = P1_U3378 & P1_U5295; 
assign P1_U2515 = P1_U3381 & P1_U5353; 
assign P1_U2517 = P1_U3385 & P1_U5410; 
assign P1_U2661 = ~(P1_U6812 & P1_U4019); 
assign P1_U3295 = ~(P1_U7604 & P1_STATE2_REG_0__SCAN_IN); 
assign P1_U3772 = P1_U5587 & P1_U5586; 
assign P1_U4517 = ~(P1_U7604 & P1_U4246); 
assign P1_U4520 = ~(P1_U2368 & P1_U7604); 
assign P1_U4522 = ~(P1_U7604 & P1_U4245); 
assign P1_U4549 = ~(P1_U2480 & P1_U2358); 
assign P1_U4555 = ~(P1_U2480 & P1_U2388); 
assign P1_U4562 = ~(P1_U2412 & P1_U4532); 
assign P1_U4567 = ~(P1_U2410 & P1_U4532); 
assign P1_U4572 = ~(P1_U2408 & P1_U4532); 
assign P1_U4577 = ~(P1_U2406 & P1_U4532); 
assign P1_U4582 = ~(P1_U2404 & P1_U4532); 
assign P1_U4587 = ~(P1_U2402 & P1_U4532); 
assign P1_U4592 = ~(P1_U2400 & P1_U4532); 
assign P1_U4597 = ~(P1_U2398 & P1_U4532); 
assign P1_U4607 = ~(P1_U2482 & P1_U2358); 
assign P1_U4613 = ~(P1_U2482 & P1_U2388); 
assign P1_U4620 = ~(P1_U4601 & P1_U2412); 
assign P1_U4625 = ~(P1_U4601 & P1_U2410); 
assign P1_U4630 = ~(P1_U4601 & P1_U2408); 
assign P1_U4635 = ~(P1_U4601 & P1_U2406); 
assign P1_U4640 = ~(P1_U4601 & P1_U2404); 
assign P1_U4645 = ~(P1_U4601 & P1_U2402); 
assign P1_U4650 = ~(P1_U4601 & P1_U2400); 
assign P1_U4655 = ~(P1_U4601 & P1_U2398); 
assign P1_U4666 = ~(P1_U2484 & P1_U2358); 
assign P1_U4672 = ~(P1_U2484 & P1_U2388); 
assign P1_U4679 = ~(P1_U4659 & P1_U2412); 
assign P1_U4684 = ~(P1_U4659 & P1_U2410); 
assign P1_U4689 = ~(P1_U4659 & P1_U2408); 
assign P1_U4694 = ~(P1_U4659 & P1_U2406); 
assign P1_U4699 = ~(P1_U4659 & P1_U2404); 
assign P1_U4704 = ~(P1_U4659 & P1_U2402); 
assign P1_U4709 = ~(P1_U4659 & P1_U2400); 
assign P1_U4714 = ~(P1_U4659 & P1_U2398); 
assign P1_U4723 = ~(P1_U2489 & P1_U2358); 
assign P1_U4729 = ~(P1_U2489 & P1_U2388); 
assign P1_U4736 = ~(P1_U4717 & P1_U2412); 
assign P1_U4741 = ~(P1_U4717 & P1_U2410); 
assign P1_U4746 = ~(P1_U4717 & P1_U2408); 
assign P1_U4751 = ~(P1_U4717 & P1_U2406); 
assign P1_U4756 = ~(P1_U4717 & P1_U2404); 
assign P1_U4761 = ~(P1_U4717 & P1_U2402); 
assign P1_U4766 = ~(P1_U4717 & P1_U2400); 
assign P1_U4771 = ~(P1_U4717 & P1_U2398); 
assign P1_U4781 = ~(P1_U2492 & P1_U2358); 
assign P1_U4787 = ~(P1_U2492 & P1_U2388); 
assign P1_U4794 = ~(P1_U4774 & P1_U2412); 
assign P1_U4799 = ~(P1_U4774 & P1_U2410); 
assign P1_U4804 = ~(P1_U4774 & P1_U2408); 
assign P1_U4809 = ~(P1_U4774 & P1_U2406); 
assign P1_U4814 = ~(P1_U4774 & P1_U2404); 
assign P1_U4819 = ~(P1_U4774 & P1_U2402); 
assign P1_U4824 = ~(P1_U4774 & P1_U2400); 
assign P1_U4829 = ~(P1_U4774 & P1_U2398); 
assign P1_U4838 = ~(P1_U2494 & P1_U2358); 
assign P1_U4844 = ~(P1_U2494 & P1_U2388); 
assign P1_U4851 = ~(P1_U4832 & P1_U2412); 
assign P1_U4856 = ~(P1_U4832 & P1_U2410); 
assign P1_U4861 = ~(P1_U4832 & P1_U2408); 
assign P1_U4866 = ~(P1_U4832 & P1_U2406); 
assign P1_U4871 = ~(P1_U4832 & P1_U2404); 
assign P1_U4876 = ~(P1_U4832 & P1_U2402); 
assign P1_U4881 = ~(P1_U4832 & P1_U2400); 
assign P1_U4886 = ~(P1_U4832 & P1_U2398); 
assign P1_U4896 = ~(P1_U2496 & P1_U2358); 
assign P1_U4902 = ~(P1_U2496 & P1_U2388); 
assign P1_U4909 = ~(P1_U4889 & P1_U2412); 
assign P1_U4914 = ~(P1_U4889 & P1_U2410); 
assign P1_U4919 = ~(P1_U4889 & P1_U2408); 
assign P1_U4924 = ~(P1_U4889 & P1_U2406); 
assign P1_U4929 = ~(P1_U4889 & P1_U2404); 
assign P1_U4934 = ~(P1_U4889 & P1_U2402); 
assign P1_U4939 = ~(P1_U4889 & P1_U2400); 
assign P1_U4944 = ~(P1_U4889 & P1_U2398); 
assign P1_U4953 = ~(P1_U2498 & P1_U2358); 
assign P1_U4959 = ~(P1_U2498 & P1_U2388); 
assign P1_U4966 = ~(P1_U4947 & P1_U2412); 
assign P1_U4971 = ~(P1_U4947 & P1_U2410); 
assign P1_U4976 = ~(P1_U4947 & P1_U2408); 
assign P1_U4981 = ~(P1_U4947 & P1_U2406); 
assign P1_U4986 = ~(P1_U4947 & P1_U2404); 
assign P1_U4991 = ~(P1_U4947 & P1_U2402); 
assign P1_U4996 = ~(P1_U4947 & P1_U2400); 
assign P1_U5001 = ~(P1_U4947 & P1_U2398); 
assign P1_U5004 = ~P1_U3359; 
assign P1_U5060 = ~P1_U3364; 
assign P1_U5117 = ~P1_U3367; 
assign P1_U5175 = ~P1_U3371; 
assign P1_U5232 = ~P1_U3374; 
assign P1_U5290 = ~P1_U3378; 
assign P1_U5347 = ~P1_U3381; 
assign P1_U5405 = ~P1_U3385; 
assign P1_U5541 = ~(P1_U3359 & P1_U5540); 
assign P1_U5717 = ~(P1_R2099_U74 & P1_U2380); 
assign P1_U5727 = ~(P1_ADD_405_U71 & P1_U2375); 
assign P1_U5728 = ~(P1_ADD_515_U71 & P1_U2374); 
assign P1_U5812 = ~(P1_R2358_U18 & P1_U2364); 
assign P1_U5817 = ~(P1_R2358_U19 & P1_U2364); 
assign P1_U5909 = ~(P1_R2337_U79 & P1_U2376); 
assign P1_U6161 = ~(P1_U2386 & P1_R2358_U18); 
assign P1_U6164 = ~(P1_U2386 & P1_R2358_U19); 
assign P1_U6271 = ~(P1_U2383 & P1_R2358_U18); 
assign P1_U6274 = ~(P1_U2383 & P1_R2358_U19); 
assign P1_U6329 = ~(P1_U2371 & P1_R2099_U74); 
assign P1_U6521 = ~(P1_U2604 & P1_R2099_U74); 
assign P1_U6529 = ~(P1_R2096_U79 & P1_U7485); 
assign P1_U6811 = ~(P1_R2337_U79 & P1_U2352); 
assign P1_U7690 = ~(P1_U7604 & P1_U4521 & P1_U3294); 
assign P1_U7735 = ~(P1_U5549 & P1_U3404); 
assign P3_ADD_476_U48 = ~(P3_ADD_476_U114 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_476_U156 = ~(P3_ADD_476_U114 & P3_ADD_476_U47); 
assign P3_ADD_531_U49 = ~(P3_ADD_531_U118 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_531_U163 = ~(P3_ADD_531_U118 & P3_ADD_531_U48); 
assign P3_SUB_320_U43 = ~P3_ADD_318_U79; 
assign P3_SUB_320_U70 = P3_SUB_320_U147 & P3_SUB_320_U146; 
assign P3_SUB_320_U114 = ~(P3_ADD_318_U79 & P3_SUB_320_U113); 
assign P3_ADD_318_U48 = ~(P3_ADD_318_U114 & P3_PHYADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_318_U156 = ~(P3_ADD_318_U114 & P3_ADD_318_U47); 
assign P3_ADD_315_U48 = ~(P3_ADD_315_U111 & P3_PHYADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_315_U148 = ~(P3_ADD_315_U111 & P3_ADD_315_U47); 
assign P3_ADD_360_1242_U11 = P3_ADD_360_1242_U174 & P3_ADD_360_1242_U60; 
assign P3_ADD_360_1242_U160 = ~P3_ADD_360_1242_U60; 
assign P3_ADD_360_1242_U242 = ~(P3_ADD_360_1242_U60 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_467_U48 = ~(P3_ADD_467_U114 & P3_REIP_REG_23__SCAN_IN); 
assign P3_ADD_467_U156 = ~(P3_ADD_467_U114 & P3_ADD_467_U47); 
assign P3_ADD_430_U48 = ~(P3_ADD_430_U114 & P3_REIP_REG_23__SCAN_IN); 
assign P3_ADD_430_U156 = ~(P3_ADD_430_U114 & P3_ADD_430_U47); 
assign P3_ADD_380_U49 = ~(P3_ADD_380_U118 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_380_U163 = ~(P3_ADD_380_U118 & P3_ADD_380_U48); 
assign P3_ADD_344_U49 = ~(P3_ADD_344_U118 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_344_U163 = ~(P3_ADD_344_U118 & P3_ADD_344_U48); 
assign P3_ADD_339_U48 = ~(P3_ADD_339_U114 & P3_PHYADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_339_U156 = ~(P3_ADD_339_U114 & P3_ADD_339_U47); 
assign P3_ADD_541_U48 = ~(P3_ADD_541_U114 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_541_U156 = ~(P3_ADD_541_U114 & P3_ADD_541_U47); 
assign P3_SUB_357_1258_U80 = ~(P3_SUB_357_1258_U384 & P3_SUB_357_1258_U383); 
assign P3_SUB_357_1258_U151 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U129); 
assign P3_SUB_357_1258_U222 = ~(P3_SUB_357_1258_U129 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_SUB_357_1258_U227 = ~(P3_SUB_357_1258_U377 & P3_SUB_357_1258_U376 & P3_SUB_357_1258_U62); 
assign P3_SUB_357_1258_U238 = ~P3_SUB_357_1258_U139; 
assign P3_SUB_357_1258_U305 = ~P3_SUB_357_1258_U129; 
assign P3_SUB_357_1258_U372 = ~(P3_SUB_357_1258_U128 & P3_SUB_357_1258_U129); 
assign P3_SUB_357_1258_U375 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U226); 
assign P3_SUB_357_1258_U418 = ~(P3_SUB_357_1258_U138 & P3_SUB_357_1258_U139); 
assign P3_SUB_357_1258_U421 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U239); 
assign P3_ADD_515_U48 = ~(P3_ADD_515_U114 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_515_U156 = ~(P3_ADD_515_U114 & P3_ADD_515_U47); 
assign P3_ADD_394_U48 = ~(P3_ADD_394_U117 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_394_U158 = ~(P3_ADD_394_U117 & P3_ADD_394_U47); 
assign P3_ADD_441_U48 = ~(P3_ADD_441_U114 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_441_U156 = ~(P3_ADD_441_U114 & P3_ADD_441_U47); 
assign P3_ADD_349_U49 = ~(P3_ADD_349_U118 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_349_U163 = ~(P3_ADD_349_U118 & P3_ADD_349_U48); 
assign P3_ADD_405_U48 = ~(P3_ADD_405_U117 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_405_U158 = ~(P3_ADD_405_U117 & P3_ADD_405_U47); 
assign P3_ADD_553_U49 = ~(P3_ADD_553_U118 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_553_U163 = ~(P3_ADD_553_U118 & P3_ADD_553_U48); 
assign P3_ADD_558_U49 = ~(P3_ADD_558_U118 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_558_U163 = ~(P3_ADD_558_U118 & P3_ADD_558_U48); 
assign P3_ADD_385_U49 = ~(P3_ADD_385_U118 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_385_U163 = ~(P3_ADD_385_U118 & P3_ADD_385_U48); 
assign P3_ADD_547_U49 = ~(P3_ADD_547_U118 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_547_U163 = ~(P3_ADD_547_U118 & P3_ADD_547_U48); 
assign P3_ADD_371_1212_U12 = P3_ADD_371_1212_U184 & P3_ADD_371_1212_U62; 
assign P3_ADD_371_1212_U65 = ~(P3_ADD_371_1212_U105 & P3_ADD_371_1212_U169); 
assign P3_ADD_371_1212_U182 = ~(P3_ADD_371_1212_U169 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_371_1212_U250 = ~(P3_ADD_371_1212_U169 & P3_ADD_371_1212_U64); 
assign P3_ADD_494_U48 = ~(P3_ADD_494_U114 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_494_U156 = ~(P3_ADD_494_U114 & P3_ADD_494_U47); 
assign P3_ADD_536_U48 = ~(P3_ADD_536_U114 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_536_U156 = ~(P3_ADD_536_U114 & P3_ADD_536_U47); 
assign P2_R2099_U91 = ~(P2_R2099_U219 & P2_R2099_U218); 
assign P2_R2099_U128 = ~P2_R2099_U31; 
assign P2_R2099_U216 = ~(P2_U2734 & P2_R2099_U31); 
assign P2_ADD_391_1196_U37 = ~(P2_ADD_391_1196_U184 & P2_ADD_391_1196_U182 & P2_ADD_391_1196_U183); 
assign P2_ADD_391_1196_U46 = ~P2_R2182_U95; 
assign P2_ADD_391_1196_U59 = ~P2_R2096_U89; 
assign P2_ADD_391_1196_U89 = ~(P2_ADD_391_1196_U322 & P2_ADD_391_1196_U321); 
assign P2_ADD_391_1196_U110 = P2_ADD_391_1196_U308 & P2_ADD_391_1196_U307; 
assign P2_ADD_391_1196_U209 = P2_R2096_U96 | P2_R2182_U95; 
assign P2_ADD_391_1196_U212 = ~(P2_R2096_U96 & P2_R2182_U95); 
assign P2_ADD_391_1196_U300 = ~(P2_R2096_U96 & P2_R2182_U95); 
assign P2_ADD_391_1196_U305 = ~(P2_ADD_391_1196_U302 & P2_ADD_391_1196_U158); 
assign P2_ADD_391_1196_U471 = ~(P2_R2182_U95 & P2_ADD_391_1196_U47); 
assign P2_ADD_391_1196_U472 = ~(P2_R2096_U97 & P2_ADD_391_1196_U48); 
assign P2_R2182_U15 = P2_U2667 & P2_R2182_U14; 
assign P2_R2182_U94 = ~(P2_R2182_U299 & P2_R2182_U298); 
assign P2_R2182_U145 = ~P2_R2182_U14; 
assign P2_R2182_U294 = ~(P2_R2182_U26 & P2_R2182_U14); 
assign P2_R2182_U297 = ~(P2_R2182_U144 & P2_U2668); 
assign P2_R2027_U49 = ~(P2_R2027_U118 & P2_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P2_R2027_U163 = ~(P2_R2027_U118 & P2_R2027_U48); 
assign P2_R2337_U49 = ~(P2_R2337_U115 & P2_PHYADDRPOINTER_REG_24__SCAN_IN); 
assign P2_R2337_U154 = ~(P2_R2337_U115 & P2_R2337_U48); 
assign P2_R2096_U8 = P2_U2628 & P2_R2096_U7; 
assign P2_R2096_U88 = ~(P2_R2096_U245 & P2_R2096_U244); 
assign P2_R2096_U156 = ~P2_R2096_U7; 
assign P2_R2096_U235 = ~(P2_R2096_U46 & P2_R2096_U7); 
assign P2_R2096_U238 = ~(P2_R2096_U155 & P2_U2629); 
assign P2_LT_563_U23 = ~(P2_LT_563_U21 & P2_LT_563_U22 & P2_LT_563_U20); 
assign P2_R2256_U41 = ~P2_R2256_U10; 
assign P2_R2256_U53 = ~(P2_U3625 & P2_R2256_U10); 
assign P2_R2256_U56 = ~(P2_R2256_U40 & P2_R2256_U9); 
assign P2_R1957_U42 = ~P2_U3668; 
assign P2_R1957_U70 = P2_R1957_U147 & P2_R1957_U146; 
assign P2_R1957_U114 = ~(P2_U3668 & P2_R1957_U113); 
assign P2_R2278_U43 = ~P2_U2806; 
assign P2_R2278_U83 = ~(P2_R2278_U562 & P2_R2278_U561); 
assign P2_R2278_U124 = P2_R2278_U324 & P2_R2278_U250; 
assign P2_R2278_U197 = P2_R2278_U534 & P2_R2278_U533; 
assign P2_R2278_U254 = ~P2_R2278_U58; 
assign P2_R2278_U256 = P2_U2806 | P2_INSTADDRPOINTER_REG_15__SCAN_IN; 
assign P2_R2278_U257 = ~(P2_U2806 & P2_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P2_R2278_U310 = ~(P2_R2278_U208 & P2_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P2_R2278_U487 = ~(P2_R2278_U208 & P2_R2278_U17); 
assign P2_R2278_U520 = ~(P2_U2806 & P2_R2278_U44); 
assign P2_R2278_U522 = ~(P2_U2806 & P2_R2278_U44); 
assign P2_R2278_U526 = ~(P2_R2278_U56 & P2_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P2_R2278_U528 = ~(P2_R2278_U56 & P2_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P2_R2278_U537 = ~(P2_R2278_U536 & P2_R2278_U535); 
assign P2_ADD_394_U48 = ~(P2_ADD_394_U117 & P2_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P2_ADD_394_U164 = ~(P2_ADD_394_U117 & P2_ADD_394_U47); 
assign P2_R2267_U9 = P2_R2267_U127 & P2_R2267_U34; 
assign P2_R2267_U35 = ~(P2_R2267_U49 & P2_R2267_U105); 
assign P2_R2267_U124 = ~(P2_R2267_U105 & P2_R2267_U78); 
assign P2_R2267_U158 = ~(P2_R2267_U105 & P2_R2267_U78); 
assign P2_ADD_371_1212_U31 = ~P2_R2256_U22; 
assign P2_ADD_371_1212_U136 = ~P2_ADD_371_1212_U67; 
assign P2_ADD_371_1212_U138 = ~(P2_ADD_371_1212_U30 & P2_ADD_371_1212_U29); 
assign P2_ADD_371_1212_U141 = P2_R2256_U22 | P2_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P2_ADD_371_1212_U143 = ~(P2_R2256_U22 & P2_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P2_ADD_371_1212_U221 = ~(P2_R2256_U22 & P2_ADD_371_1212_U32); 
assign P2_ADD_371_1212_U223 = ~(P2_R2256_U22 & P2_ADD_371_1212_U32); 
assign P2_ADD_371_1212_U269 = ~(P2_ADD_371_1212_U267 & P2_ADD_371_1212_U30); 
assign P1_R2144_U37 = ~(P1_R2144_U248 & P1_R2144_U247); 
assign P1_R2278_U5 = P1_R2278_U466 & P1_R2278_U327; 
assign P1_R2278_U7 = P1_R2278_U6 & P1_R2278_U295; 
assign P1_R2278_U13 = P1_R2278_U9 & P1_R2278_U321; 
assign P1_R2278_U65 = ~P1_U2787; 
assign P1_R2278_U67 = ~P1_U2786; 
assign P1_R2278_U73 = ~(P1_R2278_U12 & P1_R2278_U8 & P1_R2278_U359 & P1_R2278_U308); 
assign P1_R2278_U80 = ~(P1_R2278_U144 & P1_R2278_U8); 
assign P1_R2278_U86 = ~(P1_R2278_U379 & P1_R2278_U322); 
assign P1_R2278_U92 = ~(P1_R2278_U143 & P1_R2278_U11); 
assign P1_R2278_U105 = ~(P1_R2278_U461 & P1_R2278_U460); 
assign P1_R2278_U129 = P1_R2278_U352 & P1_R2278_U259; 
assign P1_R2278_U136 = P1_R2278_U11 & P1_R2278_U135; 
assign P1_R2278_U150 = P1_R2278_U11 & P1_R2278_U149; 
assign P1_R2278_U152 = P1_R2278_U11 & P1_R2278_U324; 
assign P1_R2278_U157 = P1_R2278_U11 & P1_R2278_U324; 
assign P1_R2278_U175 = P1_R2278_U603 & P1_R2278_U602 & P1_R2278_U228; 
assign P1_R2278_U177 = P1_R2278_U433 & P1_R2278_U432; 
assign P1_R2278_U221 = P1_R2278_U582 & P1_R2278_U581; 
assign P1_R2278_U229 = ~(P1_U2787 & P1_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P1_R2278_U243 = ~P1_R2278_U182; 
assign P1_R2278_U245 = ~(P1_R2278_U244 & P1_R2278_U182); 
assign P1_R2278_U283 = P1_U2787 | P1_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P1_R2278_U284 = P1_U2786 | P1_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P1_R2278_U285 = ~(P1_U2786 & P1_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P1_R2278_U330 = P1_U2787 | P1_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P1_R2278_U333 = P1_U2786 | P1_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P1_R2278_U338 = P1_U2786 | P1_INSTADDRPOINTER_REG_14__SCAN_IN; 
assign P1_R2278_U339 = P1_U2787 | P1_INSTADDRPOINTER_REG_13__SCAN_IN; 
assign P1_R2278_U360 = ~(P1_R2278_U359 & P1_R2278_U292); 
assign P1_R2278_U362 = ~(P1_R2278_U12 & P1_R2278_U359); 
assign P1_R2278_U367 = ~(P1_R2278_U366 & P1_R2278_U305); 
assign P1_R2278_U371 = ~(P1_R2278_U381 & P1_R2278_U315); 
assign P1_R2278_U389 = ~(P1_R2278_U388 & P1_R2278_U228); 
assign P1_R2278_U436 = ~(P1_R2278_U435 & P1_R2278_U434); 
assign P1_R2278_U453 = ~(P1_R2278_U181 & P1_R2278_U182); 
assign P1_R2278_U469 = ~(P1_R2278_U14 & P1_R2278_U88 & P1_R2278_U89); 
assign P1_R2278_U470 = ~(P1_U2770 & P1_R2278_U466 & P1_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P1_R2278_U585 = ~(P1_R2278_U584 & P1_R2278_U583); 
assign P1_R2278_U590 = ~(P1_U2786 & P1_R2278_U66); 
assign P1_R2278_U595 = ~(P1_U2787 & P1_R2278_U64); 
assign P1_R2278_U606 = ~(P1_R2278_U605 & P1_R2278_U604); 
assign P1_R2358_U5 = P1_R2358_U274 & P1_R2358_U272; 
assign P1_R2358_U47 = ~(P1_U2631 & P1_R2358_U521); 
assign P1_R2358_U58 = ~P1_U2637; 
assign P1_R2358_U59 = ~(P1_U2637 & P1_R2358_U463); 
assign P1_R2358_U60 = ~P1_U2636; 
assign P1_R2358_U61 = ~(P1_U2636 & P1_R2358_U466); 
assign P1_R2358_U77 = P1_R2358_U233 & P1_R2358_U54; 
assign P1_R2358_U114 = P1_R2358_U51 & P1_R2358_U272; 
assign P1_R2358_U118 = P1_R2358_U57 & P1_R2358_U259; 
assign P1_R2358_U124 = P1_R2358_U229 & P1_R2358_U54; 
assign P1_R2358_U125 = P1_R2358_U265 & P1_R2358_U262; 
assign P1_R2358_U141 = P1_R2358_U265 & P1_R2358_U264; 
assign P1_R2358_U154 = ~(P1_R2358_U226 & P1_R2358_U216 & P1_R2358_U224); 
assign P1_R2358_U155 = ~(P1_R2358_U28 & P1_R2358_U234); 
assign P1_R2358_U232 = ~P1_R2358_U54; 
assign P1_R2358_U326 = ~(P1_R2358_U265 & P1_R2358_U264); 
assign P1_R2358_U328 = ~(P1_R2358_U263 & P1_R2358_U262); 
assign P1_R2358_U332 = ~(P1_R2358_U233 & P1_R2358_U54); 
assign P1_R2358_U350 = ~(P1_R2358_U51 & P1_R2358_U272); 
assign P1_R2358_U352 = ~(P1_R2358_U57 & P1_R2358_U259); 
assign P1_R2358_U358 = ~(P1_R2358_U273 & P1_R2358_U274); 
assign P1_R2358_U456 = ~(P1_R2358_U83 & P1_R2358_U214); 
assign P1_R2358_U508 = ~(P1_U2352 & P1_R2358_U169); 
assign P1_R2358_U516 = ~(P1_U2352 & P1_R2358_U169); 
assign P1_R2099_U19 = ~(P1_R2099_U173 & P1_R2099_U51); 
assign P1_R2099_U312 = ~(P1_R2099_U246 & P1_R2099_U173); 
assign P1_R2337_U48 = ~(P1_R2337_U114 & P1_PHYADDRPOINTER_REG_23__SCAN_IN); 
assign P1_R2337_U156 = ~(P1_R2337_U114 & P1_R2337_U47); 
assign P1_R2096_U48 = ~(P1_R2096_U114 & P1_REIP_REG_23__SCAN_IN); 
assign P1_R2096_U156 = ~(P1_R2096_U114 & P1_R2096_U47); 
assign P1_ADD_405_U48 = ~(P1_ADD_405_U117 & P1_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P1_ADD_405_U164 = ~(P1_ADD_405_U117 & P1_ADD_405_U47); 
assign P1_ADD_515_U48 = ~(P1_ADD_515_U114 & P1_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P1_ADD_515_U162 = ~(P1_ADD_515_U114 & P1_ADD_515_U47); 
assign P3_U2811 = ~(P3_U6558 & P3_U6557 & P3_U6559 & P3_U6560 & P3_U3973); 
assign P3_U2845 = ~(P3_U6063 & P3_U6061 & P3_U6062); 
assign P3_U2847 = ~(P3_U3811 & P3_U6014); 
assign P3_U2996 = ~(P3_U7959 & P3_U7958 & P3_U3367); 
assign P3_U2998 = ~(P3_U3363 & P3_U4632); 
assign P3_U3844 = P3_U3843 & P3_U3842 & P3_U6131; 
assign P3_U3846 = P3_U6140 & P3_U6139; 
assign P3_U3848 = P3_U6142 & P3_U6141 & P3_U6143 & P3_U3847; 
assign P3_U3851 = P3_U6154 & P3_U6153 & P3_U6152 & P3_U6151; 
assign P3_U3855 = P3_U6169 & P3_U6168; 
assign P3_U3858 = P3_U6171 & P3_U6170 & P3_U6172; 
assign P3_U3859 = P3_U6174 & P3_U6173; 
assign P3_U3974 = P3_U6572 & P3_U6569 & P3_U6570 & P3_U6571; 
assign P3_U4105 = P3_U7286 & P3_U7285; 
assign P3_U4634 = ~(P3_U3364 & P3_U4630); 
assign P3_U6086 = ~(P3_U4318 & P3_U6084); 
assign P3_U6108 = ~(P3_U6090 & P3_U3832 & P3_U6088 & P3_U3837 & P3_U3833); 
assign P3_U6136 = ~(P3_ADD_360_1242_U11 & P3_U2395); 
assign P3_U6155 = ~(P3_ADD_371_1212_U12 & P3_U2360); 
assign P3_U6281 = ~(P3_SUB_357_1258_U80 & P3_U2393); 
assign P3_U6575 = ~(P3_U2396 & P3_ADD_360_1242_U11); 
assign P3_U6579 = ~(P3_U2387 & P3_ADD_371_1212_U12); 
assign P3_U6624 = ~(P3_U2394 & P3_SUB_357_1258_U80); 
assign P3_U7955 = ~(P3_U2453 & P3_U4630); 
assign P2_U2804 = P2_U3242 & P2_R2267_U9; 
assign P2_U2876 = ~(P2_U6505 & P2_U6506 & P2_U6504); 
assign P2_U2914 = ~(P2_U6348 & P2_U6347 & P2_U4064); 
assign P2_U3636 = ~(P2_U8326 & P2_U8325); 
assign P2_U3667 = ~(P2_U8390 & P2_U8389); 
assign P2_U4125 = P2_U6707 & P2_U4446; 
assign P2_U4663 = ~(P2_U4660 & P2_U3722); 
assign P2_U4668 = ~(P2_U4667 & P2_U4666); 
assign P2_U4721 = ~(P2_U4718 & P2_U3731); 
assign P2_U4726 = ~(P2_U4725 & P2_U4724); 
assign P2_U4780 = ~(P2_U4777 & P2_U3740); 
assign P2_U4785 = ~(P2_U4784 & P2_U4783); 
assign P2_U4837 = ~(P2_U4834 & P2_U3749); 
assign P2_U4842 = ~(P2_U4841 & P2_U4840); 
assign P2_U4895 = ~(P2_U4892 & P2_U3758); 
assign P2_U4900 = ~(P2_U4899 & P2_U4898); 
assign P2_U4952 = ~(P2_U4949 & P2_U3767); 
assign P2_U4957 = ~(P2_U4956 & P2_U4955); 
assign P2_U5010 = ~(P2_U5007 & P2_U3776); 
assign P2_U5015 = ~(P2_U5014 & P2_U5013); 
assign P2_U5067 = ~(P2_U5064 & P2_U3785); 
assign P2_U5072 = ~(P2_U5071 & P2_U5070); 
assign P2_U5120 = ~(P2_U5115 & P2_U5119); 
assign P2_U5126 = ~(P2_U5125 & P2_U3429); 
assign P2_U5177 = ~(P2_U5176 & P2_U3249); 
assign P2_U5183 = ~(P2_U5182 & P2_U5171); 
assign P2_U5235 = ~(P2_U5229 & P2_U5234); 
assign P2_U5241 = ~(P2_U5240 & P2_U3452); 
assign P2_U5292 = ~(P2_U5291 & P2_U3250); 
assign P2_U5298 = ~(P2_U5297 & P2_U5286); 
assign P2_U5350 = ~(P2_U5344 & P2_U5349); 
assign P2_U5356 = ~(P2_U5355 & P2_U3475); 
assign P2_U5407 = ~(P2_U5406 & P2_U3251); 
assign P2_U5413 = ~(P2_U5412 & P2_U5401); 
assign P2_U5465 = ~(P2_U5459 & P2_U5464); 
assign P2_U5471 = ~(P2_U5470 & P2_U3498); 
assign P2_U5522 = ~(P2_U5521 & P2_U3252); 
assign P2_U5528 = ~(P2_U5527 & P2_U5516); 
assign P2_U6352 = ~(P2_ADD_391_1196_U89 & P2_U2397); 
assign P2_U6409 = ~(P2_U2380 & P2_R2096_U88); 
assign P2_U6507 = ~(P2_R2182_U94 & P2_U2393); 
assign P2_U6508 = ~(P2_U2379 & P2_R2099_U91); 
assign P2_U6678 = ~(P2_U2392 & P2_R2099_U91); 
assign P2_U6715 = ~(P2_R2267_U9 & P2_U2587); 
assign P2_U6732 = ~(P2_U2588 & P2_R2096_U88); 
assign P1_U2635 = P1_R2144_U37 & P1_U6746; 
assign P1_U2785 = P1_U4159 & P1_R2144_U37; 
assign P1_U2869 = ~(P1_U6275 & P1_U6276 & P1_U6274); 
assign P1_U2870 = ~(P1_U6272 & P1_U6273 & P1_U6271); 
assign P1_U2901 = ~(P1_U6165 & P1_U6163 & P1_U6164); 
assign P1_U2902 = ~(P1_U6162 & P1_U6160 & P1_U6161); 
assign P1_U2997 = ~(P1_U5811 & P1_U5809 & P1_U5810 & P1_U5813 & P1_U5812); 
assign P1_U3029 = ~(P1_U3772 & P1_U3771 & P1_U3774); 
assign P1_U3476 = ~(P1_U7735 & P1_U7734); 
assign P1_U3588 = P1_U4561 & P1_U4560 & P1_U4562; 
assign P1_U3589 = P1_U4566 & P1_U4565 & P1_U4567; 
assign P1_U3590 = P1_U4571 & P1_U4570 & P1_U4572; 
assign P1_U3591 = P1_U4576 & P1_U4575 & P1_U4577; 
assign P1_U3592 = P1_U4581 & P1_U4580 & P1_U4582; 
assign P1_U3593 = P1_U4586 & P1_U4585 & P1_U4587; 
assign P1_U3594 = P1_U4591 & P1_U4590 & P1_U4592; 
assign P1_U3595 = P1_U4596 & P1_U4595 & P1_U4597; 
assign P1_U3597 = P1_U4619 & P1_U4618 & P1_U4620; 
assign P1_U3598 = P1_U4624 & P1_U4623 & P1_U4625; 
assign P1_U3599 = P1_U4629 & P1_U4628 & P1_U4630; 
assign P1_U3600 = P1_U4634 & P1_U4633 & P1_U4635; 
assign P1_U3601 = P1_U4639 & P1_U4638 & P1_U4640; 
assign P1_U3602 = P1_U4644 & P1_U4643 & P1_U4645; 
assign P1_U3603 = P1_U4649 & P1_U4648 & P1_U4650; 
assign P1_U3604 = P1_U4654 & P1_U4653 & P1_U4655; 
assign P1_U3606 = P1_U4678 & P1_U4677 & P1_U4679; 
assign P1_U3607 = P1_U4683 & P1_U4682 & P1_U4684; 
assign P1_U3608 = P1_U4688 & P1_U4687 & P1_U4689; 
assign P1_U3609 = P1_U4693 & P1_U4692 & P1_U4694; 
assign P1_U3610 = P1_U4698 & P1_U4697 & P1_U4699; 
assign P1_U3611 = P1_U4703 & P1_U4702 & P1_U4704; 
assign P1_U3612 = P1_U4708 & P1_U4707 & P1_U4709; 
assign P1_U3613 = P1_U4713 & P1_U4712 & P1_U4714; 
assign P1_U3615 = P1_U4735 & P1_U4734 & P1_U4736; 
assign P1_U3616 = P1_U4740 & P1_U4739 & P1_U4741; 
assign P1_U3617 = P1_U4745 & P1_U4744 & P1_U4746; 
assign P1_U3618 = P1_U4750 & P1_U4749 & P1_U4751; 
assign P1_U3619 = P1_U4755 & P1_U4754 & P1_U4756; 
assign P1_U3620 = P1_U4760 & P1_U4759 & P1_U4761; 
assign P1_U3621 = P1_U4765 & P1_U4764 & P1_U4766; 
assign P1_U3622 = P1_U4770 & P1_U4769 & P1_U4771; 
assign P1_U3624 = P1_U4793 & P1_U4792 & P1_U4794; 
assign P1_U3625 = P1_U4798 & P1_U4797 & P1_U4799; 
assign P1_U3626 = P1_U4803 & P1_U4802 & P1_U4804; 
assign P1_U3627 = P1_U4808 & P1_U4807 & P1_U4809; 
assign P1_U3628 = P1_U4813 & P1_U4812 & P1_U4814; 
assign P1_U3629 = P1_U4818 & P1_U4817 & P1_U4819; 
assign P1_U3630 = P1_U4823 & P1_U4822 & P1_U4824; 
assign P1_U3631 = P1_U4828 & P1_U4827 & P1_U4829; 
assign P1_U3633 = P1_U4850 & P1_U4849 & P1_U4851; 
assign P1_U3634 = P1_U4855 & P1_U4854 & P1_U4856; 
assign P1_U3635 = P1_U4860 & P1_U4859 & P1_U4861; 
assign P1_U3636 = P1_U4865 & P1_U4864 & P1_U4866; 
assign P1_U3637 = P1_U4870 & P1_U4869 & P1_U4871; 
assign P1_U3638 = P1_U4875 & P1_U4874 & P1_U4876; 
assign P1_U3639 = P1_U4880 & P1_U4879 & P1_U4881; 
assign P1_U3640 = P1_U4885 & P1_U4884 & P1_U4886; 
assign P1_U3642 = P1_U4908 & P1_U4907 & P1_U4909; 
assign P1_U3643 = P1_U4913 & P1_U4912 & P1_U4914; 
assign P1_U3644 = P1_U4918 & P1_U4917 & P1_U4919; 
assign P1_U3645 = P1_U4923 & P1_U4922 & P1_U4924; 
assign P1_U3646 = P1_U4928 & P1_U4927 & P1_U4929; 
assign P1_U3647 = P1_U4933 & P1_U4932 & P1_U4934; 
assign P1_U3648 = P1_U4938 & P1_U4937 & P1_U4939; 
assign P1_U3649 = P1_U4943 & P1_U4942 & P1_U4944; 
assign P1_U3651 = P1_U4965 & P1_U4964 & P1_U4966; 
assign P1_U3652 = P1_U4970 & P1_U4969 & P1_U4971; 
assign P1_U3653 = P1_U4975 & P1_U4974 & P1_U4976; 
assign P1_U3654 = P1_U4980 & P1_U4979 & P1_U4981; 
assign P1_U3655 = P1_U4985 & P1_U4984 & P1_U4986; 
assign P1_U3656 = P1_U4990 & P1_U4989 & P1_U4991; 
assign P1_U3657 = P1_U4995 & P1_U4994 & P1_U4996; 
assign P1_U3658 = P1_U5000 & P1_U4999 & P1_U5001; 
assign P1_U3832 = P1_U5725 & P1_U5727; 
assign P1_U3834 = P1_U3833 & P1_U5728; 
assign P1_U3930 = P1_U6531 & P1_U6529; 
assign P1_U4018 = P1_U6809 & P1_U6810 & P1_U6811; 
assign P1_U4514 = ~P1_U3295; 
assign P1_U4516 = ~(P1_U3295 & P1_STATE2_REG_2__SCAN_IN); 
assign P1_U4519 = ~(P1_U4517 & P1_STATE2_REG_1__SCAN_IN); 
assign P1_U4550 = ~(P1_U3320 & P1_U4549); 
assign P1_U4556 = ~(P1_U3320 & P1_U4555); 
assign P1_U4608 = ~(P1_U3320 & P1_U4607); 
assign P1_U4614 = ~(P1_U3320 & P1_U4613); 
assign P1_U4667 = ~(P1_U3320 & P1_U4666); 
assign P1_U4673 = ~(P1_U3320 & P1_U4672); 
assign P1_U4724 = ~(P1_U3320 & P1_U4723); 
assign P1_U4730 = ~(P1_U3320 & P1_U4729); 
assign P1_U4782 = ~(P1_U3320 & P1_U4781); 
assign P1_U4788 = ~(P1_U3320 & P1_U4787); 
assign P1_U4839 = ~(P1_U3320 & P1_U4838); 
assign P1_U4845 = ~(P1_U3320 & P1_U4844); 
assign P1_U4897 = ~(P1_U3320 & P1_U4896); 
assign P1_U4903 = ~(P1_U3320 & P1_U4902); 
assign P1_U4954 = ~(P1_U3320 & P1_U4953); 
assign P1_U4960 = ~(P1_U3320 & P1_U4959); 
assign P1_U5009 = ~(P1_U2500 & P1_U2358); 
assign P1_U5015 = ~(P1_U2500 & P1_U2388); 
assign P1_U5022 = ~(P1_U5004 & P1_U2412); 
assign P1_U5027 = ~(P1_U5004 & P1_U2410); 
assign P1_U5032 = ~(P1_U5004 & P1_U2408); 
assign P1_U5037 = ~(P1_U5004 & P1_U2406); 
assign P1_U5042 = ~(P1_U5004 & P1_U2404); 
assign P1_U5047 = ~(P1_U5004 & P1_U2402); 
assign P1_U5052 = ~(P1_U5004 & P1_U2400); 
assign P1_U5057 = ~(P1_U5004 & P1_U2398); 
assign P1_U5066 = ~(P1_U2502 & P1_U2358); 
assign P1_U5072 = ~(P1_U2502 & P1_U2388); 
assign P1_U5079 = ~(P1_U5060 & P1_U2412); 
assign P1_U5084 = ~(P1_U5060 & P1_U2410); 
assign P1_U5089 = ~(P1_U5060 & P1_U2408); 
assign P1_U5094 = ~(P1_U5060 & P1_U2406); 
assign P1_U5099 = ~(P1_U5060 & P1_U2404); 
assign P1_U5104 = ~(P1_U5060 & P1_U2402); 
assign P1_U5109 = ~(P1_U5060 & P1_U2400); 
assign P1_U5114 = ~(P1_U5060 & P1_U2398); 
assign P1_U5124 = ~(P1_U2504 & P1_U2358); 
assign P1_U5130 = ~(P1_U2504 & P1_U2388); 
assign P1_U5137 = ~(P1_U5117 & P1_U2412); 
assign P1_U5142 = ~(P1_U5117 & P1_U2410); 
assign P1_U5147 = ~(P1_U5117 & P1_U2408); 
assign P1_U5152 = ~(P1_U5117 & P1_U2406); 
assign P1_U5157 = ~(P1_U5117 & P1_U2404); 
assign P1_U5162 = ~(P1_U5117 & P1_U2402); 
assign P1_U5167 = ~(P1_U5117 & P1_U2400); 
assign P1_U5172 = ~(P1_U5117 & P1_U2398); 
assign P1_U5181 = ~(P1_U2506 & P1_U2358); 
assign P1_U5187 = ~(P1_U2506 & P1_U2388); 
assign P1_U5194 = ~(P1_U5175 & P1_U2412); 
assign P1_U5199 = ~(P1_U5175 & P1_U2410); 
assign P1_U5204 = ~(P1_U5175 & P1_U2408); 
assign P1_U5209 = ~(P1_U5175 & P1_U2406); 
assign P1_U5214 = ~(P1_U5175 & P1_U2404); 
assign P1_U5219 = ~(P1_U5175 & P1_U2402); 
assign P1_U5224 = ~(P1_U5175 & P1_U2400); 
assign P1_U5229 = ~(P1_U5175 & P1_U2398); 
assign P1_U5239 = ~(P1_U2511 & P1_U2358); 
assign P1_U5245 = ~(P1_U2511 & P1_U2388); 
assign P1_U5252 = ~(P1_U5232 & P1_U2412); 
assign P1_U5257 = ~(P1_U5232 & P1_U2410); 
assign P1_U5262 = ~(P1_U5232 & P1_U2408); 
assign P1_U5267 = ~(P1_U5232 & P1_U2406); 
assign P1_U5272 = ~(P1_U5232 & P1_U2404); 
assign P1_U5277 = ~(P1_U5232 & P1_U2402); 
assign P1_U5282 = ~(P1_U5232 & P1_U2400); 
assign P1_U5287 = ~(P1_U5232 & P1_U2398); 
assign P1_U5296 = ~(P1_U2513 & P1_U2358); 
assign P1_U5302 = ~(P1_U2513 & P1_U2388); 
assign P1_U5309 = ~(P1_U5290 & P1_U2412); 
assign P1_U5314 = ~(P1_U5290 & P1_U2410); 
assign P1_U5319 = ~(P1_U5290 & P1_U2408); 
assign P1_U5324 = ~(P1_U5290 & P1_U2406); 
assign P1_U5329 = ~(P1_U5290 & P1_U2404); 
assign P1_U5334 = ~(P1_U5290 & P1_U2402); 
assign P1_U5339 = ~(P1_U5290 & P1_U2400); 
assign P1_U5344 = ~(P1_U5290 & P1_U2398); 
assign P1_U5354 = ~(P1_U2515 & P1_U2358); 
assign P1_U5360 = ~(P1_U2515 & P1_U2388); 
assign P1_U5367 = ~(P1_U5347 & P1_U2412); 
assign P1_U5372 = ~(P1_U5347 & P1_U2410); 
assign P1_U5377 = ~(P1_U5347 & P1_U2408); 
assign P1_U5382 = ~(P1_U5347 & P1_U2406); 
assign P1_U5387 = ~(P1_U5347 & P1_U2404); 
assign P1_U5392 = ~(P1_U5347 & P1_U2402); 
assign P1_U5397 = ~(P1_U5347 & P1_U2400); 
assign P1_U5402 = ~(P1_U5347 & P1_U2398); 
assign P1_U5411 = ~(P1_U2517 & P1_U2358); 
assign P1_U5417 = ~(P1_U2517 & P1_U2388); 
assign P1_U5424 = ~(P1_U5405 & P1_U2412); 
assign P1_U5429 = ~(P1_U5405 & P1_U2410); 
assign P1_U5434 = ~(P1_U5405 & P1_U2408); 
assign P1_U5439 = ~(P1_U5405 & P1_U2406); 
assign P1_U5443 = ~(P1_U5405 & P1_U2404); 
assign P1_U5448 = ~(P1_U5405 & P1_U2402); 
assign P1_U5453 = ~(P1_U5405 & P1_U2400); 
assign P1_U5458 = ~(P1_U5405 & P1_U2398); 
assign P1_U5542 = ~(P1_U2388 & P1_U5541); 
assign P1_U5593 = ~(P1_R2278_U105 & P1_U2377); 
assign P1_U5815 = ~(P1_U2372 & P1_R2278_U105); 
assign P1_U7685 = ~(P1_U3295 & P1_STATE2_REG_3__SCAN_IN); 
assign P1_U7689 = ~(P1_U4522 & P1_STATE2_REG_0__SCAN_IN); 
assign P3_ADD_476_U78 = ~(P3_ADD_476_U156 & P3_ADD_476_U155); 
assign P3_ADD_476_U115 = ~P3_ADD_476_U48; 
assign P3_ADD_476_U153 = ~(P3_ADD_476_U48 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_531_U82 = ~(P3_ADD_531_U163 & P3_ADD_531_U162); 
assign P3_ADD_531_U119 = ~P3_ADD_531_U49; 
assign P3_ADD_531_U160 = ~(P3_ADD_531_U49 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_SUB_320_U34 = ~(P3_SUB_320_U43 & P3_SUB_320_U69 & P3_SUB_320_U98); 
assign P3_ADD_318_U78 = ~(P3_ADD_318_U156 & P3_ADD_318_U155); 
assign P3_ADD_318_U115 = ~P3_ADD_318_U48; 
assign P3_ADD_318_U153 = ~(P3_ADD_318_U48 & P3_PHYADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_315_U74 = ~(P3_ADD_315_U148 & P3_ADD_315_U147); 
assign P3_ADD_315_U112 = ~P3_ADD_315_U48; 
assign P3_ADD_315_U145 = ~(P3_ADD_315_U48 & P3_PHYADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_360_1242_U63 = ~(P3_ADD_360_1242_U102 & P3_ADD_360_1242_U160); 
assign P3_ADD_360_1242_U172 = ~(P3_ADD_360_1242_U160 & P3_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P3_ADD_360_1242_U243 = ~(P3_ADD_360_1242_U160 & P3_ADD_360_1242_U62); 
assign P3_ADD_467_U78 = ~(P3_ADD_467_U156 & P3_ADD_467_U155); 
assign P3_ADD_467_U115 = ~P3_ADD_467_U48; 
assign P3_ADD_467_U153 = ~(P3_ADD_467_U48 & P3_REIP_REG_24__SCAN_IN); 
assign P3_ADD_430_U78 = ~(P3_ADD_430_U156 & P3_ADD_430_U155); 
assign P3_ADD_430_U115 = ~P3_ADD_430_U48; 
assign P3_ADD_430_U153 = ~(P3_ADD_430_U48 & P3_REIP_REG_24__SCAN_IN); 
assign P3_ADD_380_U82 = ~(P3_ADD_380_U163 & P3_ADD_380_U162); 
assign P3_ADD_380_U119 = ~P3_ADD_380_U49; 
assign P3_ADD_380_U160 = ~(P3_ADD_380_U49 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_344_U82 = ~(P3_ADD_344_U163 & P3_ADD_344_U162); 
assign P3_ADD_344_U119 = ~P3_ADD_344_U49; 
assign P3_ADD_344_U160 = ~(P3_ADD_344_U49 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_339_U78 = ~(P3_ADD_339_U156 & P3_ADD_339_U155); 
assign P3_ADD_339_U115 = ~P3_ADD_339_U48; 
assign P3_ADD_339_U153 = ~(P3_ADD_339_U48 & P3_PHYADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_541_U78 = ~(P3_ADD_541_U156 & P3_ADD_541_U155); 
assign P3_ADD_541_U115 = ~P3_ADD_541_U48; 
assign P3_ADD_541_U153 = ~(P3_ADD_541_U48 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_SUB_357_1258_U61 = ~(P3_SUB_357_1258_U222 & P3_SUB_357_1258_U151 & P3_SUB_357_1258_U269); 
assign P3_SUB_357_1258_U224 = ~(P3_SUB_357_1258_U151 & P3_SUB_357_1258_U107); 
assign P3_SUB_357_1258_U241 = ~(P3_SUB_357_1258_U421 & P3_SUB_357_1258_U420 & P3_SUB_357_1258_U240); 
assign P3_SUB_357_1258_U303 = ~(P3_SUB_357_1258_U375 & P3_SUB_357_1258_U374 & P3_SUB_357_1258_U302); 
assign P3_SUB_357_1258_U373 = ~(P3_SUB_357_1258_U305 & P3_SUB_357_1258_U371); 
assign P3_SUB_357_1258_U419 = ~(P3_SUB_357_1258_U238 & P3_SUB_357_1258_U417); 
assign P3_ADD_515_U78 = ~(P3_ADD_515_U156 & P3_ADD_515_U155); 
assign P3_ADD_515_U115 = ~P3_ADD_515_U48; 
assign P3_ADD_515_U153 = ~(P3_ADD_515_U48 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_394_U77 = ~(P3_ADD_394_U158 & P3_ADD_394_U157); 
assign P3_ADD_394_U118 = ~P3_ADD_394_U48; 
assign P3_ADD_394_U155 = ~(P3_ADD_394_U48 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_441_U78 = ~(P3_ADD_441_U156 & P3_ADD_441_U155); 
assign P3_ADD_441_U115 = ~P3_ADD_441_U48; 
assign P3_ADD_441_U153 = ~(P3_ADD_441_U48 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_349_U82 = ~(P3_ADD_349_U163 & P3_ADD_349_U162); 
assign P3_ADD_349_U119 = ~P3_ADD_349_U49; 
assign P3_ADD_349_U160 = ~(P3_ADD_349_U49 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_405_U77 = ~(P3_ADD_405_U158 & P3_ADD_405_U157); 
assign P3_ADD_405_U118 = ~P3_ADD_405_U48; 
assign P3_ADD_405_U155 = ~(P3_ADD_405_U48 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_553_U82 = ~(P3_ADD_553_U163 & P3_ADD_553_U162); 
assign P3_ADD_553_U119 = ~P3_ADD_553_U49; 
assign P3_ADD_553_U160 = ~(P3_ADD_553_U49 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_558_U82 = ~(P3_ADD_558_U163 & P3_ADD_558_U162); 
assign P3_ADD_558_U119 = ~P3_ADD_558_U49; 
assign P3_ADD_558_U160 = ~(P3_ADD_558_U49 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_385_U82 = ~(P3_ADD_385_U163 & P3_ADD_385_U162); 
assign P3_ADD_385_U119 = ~P3_ADD_385_U49; 
assign P3_ADD_385_U160 = ~(P3_ADD_385_U49 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_547_U82 = ~(P3_ADD_547_U163 & P3_ADD_547_U162); 
assign P3_ADD_547_U119 = ~P3_ADD_547_U49; 
assign P3_ADD_547_U160 = ~(P3_ADD_547_U49 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_371_1212_U82 = ~(P3_ADD_371_1212_U250 & P3_ADD_371_1212_U249); 
assign P3_ADD_371_1212_U170 = ~P3_ADD_371_1212_U65; 
assign P3_ADD_371_1212_U183 = ~(P3_ADD_371_1212_U63 & P3_ADD_371_1212_U182); 
assign P3_ADD_371_1212_U247 = ~(P3_ADD_371_1212_U65 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_494_U78 = ~(P3_ADD_494_U156 & P3_ADD_494_U155); 
assign P3_ADD_494_U115 = ~P3_ADD_494_U48; 
assign P3_ADD_494_U153 = ~(P3_ADD_494_U48 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_536_U78 = ~(P3_ADD_536_U156 & P3_ADD_536_U155); 
assign P3_ADD_536_U115 = ~P3_ADD_536_U48; 
assign P3_ADD_536_U153 = ~(P3_ADD_536_U48 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P2_R2099_U33 = ~(P2_U2734 & P2_R2099_U128); 
assign P2_R2099_U217 = ~(P2_R2099_U128 & P2_R2099_U32); 
assign P2_ADD_391_1196_U51 = ~P2_R2182_U94; 
assign P2_ADD_391_1196_U61 = ~P2_R2096_U88; 
assign P2_ADD_391_1196_U112 = ~(P2_ADD_391_1196_U37 & P2_ADD_391_1196_U186); 
assign P2_ADD_391_1196_U185 = ~P2_ADD_391_1196_U37; 
assign P2_ADD_391_1196_U214 = P2_R2182_U94 | P2_R2096_U95; 
assign P2_ADD_391_1196_U216 = ~(P2_R2096_U95 & P2_R2182_U94); 
assign P2_ADD_391_1196_U464 = ~(P2_R2182_U94 & P2_ADD_391_1196_U52); 
assign P2_ADD_391_1196_U466 = ~(P2_R2182_U94 & P2_ADD_391_1196_U52); 
assign P2_ADD_391_1196_U470 = ~(P2_R2096_U96 & P2_ADD_391_1196_U46); 
assign P2_ADD_391_1196_U474 = ~(P2_ADD_391_1196_U473 & P2_ADD_391_1196_U472); 
assign P2_R2182_U16 = P2_U2666 & P2_R2182_U15; 
assign P2_R2182_U93 = ~(P2_R2182_U297 & P2_R2182_U296); 
assign P2_R2182_U146 = ~P2_R2182_U15; 
assign P2_R2182_U292 = ~(P2_R2182_U25 & P2_R2182_U15); 
assign P2_R2182_U295 = ~(P2_R2182_U145 & P2_U2667); 
assign P2_R2027_U82 = ~(P2_R2027_U163 & P2_R2027_U162); 
assign P2_R2027_U119 = ~P2_R2027_U49; 
assign P2_R2027_U160 = ~(P2_R2027_U49 & P2_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P2_R2337_U76 = ~(P2_R2337_U154 & P2_R2337_U153); 
assign P2_R2337_U116 = ~P2_R2337_U49; 
assign P2_R2337_U151 = ~(P2_R2337_U49 & P2_PHYADDRPOINTER_REG_25__SCAN_IN); 
assign P2_R2096_U9 = P2_U2627 & P2_R2096_U8; 
assign P2_R2096_U87 = ~(P2_R2096_U238 & P2_R2096_U237); 
assign P2_R2096_U157 = ~P2_R2096_U8; 
assign P2_R2096_U233 = ~(P2_R2096_U39 & P2_R2096_U8); 
assign P2_R2096_U236 = ~(P2_R2096_U156 & P2_U2628); 
assign P2_LT_563_U26 = ~(P2_LT_563_U24 & P2_LT_563_U25 & P2_LT_563_U23); 
assign P2_R2256_U12 = ~(P2_U3625 & P2_R2256_U41); 
assign P2_R2256_U26 = P2_R2256_U56 & P2_R2256_U55; 
assign P2_R2256_U54 = ~(P2_R2256_U41 & P2_R2256_U11); 
assign P2_R1957_U33 = ~(P2_R1957_U98 & P2_R1957_U69 & P2_R1957_U42); 
assign P2_R2278_U16 = ~P2_U3637; 
assign P2_R2278_U59 = ~P2_U2805; 
assign P2_R2278_U61 = ~(P2_U2805 & P2_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P2_R2278_U82 = ~(P2_U3637 & P2_R2278_U208); 
assign P2_R2278_U125 = P2_R2278_U252 & P2_R2278_U256; 
assign P2_R2278_U195 = P2_R2278_U527 & P2_R2278_U526; 
assign P2_R2278_U259 = P2_U2805 | P2_INSTADDRPOINTER_REG_16__SCAN_IN; 
assign P2_R2278_U311 = ~(P2_U3637 & P2_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P2_R2278_U326 = ~(P2_R2278_U254 & P2_R2278_U256); 
assign P2_R2278_U488 = ~(P2_R2278_U487 & P2_R2278_U486); 
assign P2_R2278_U489 = ~(P2_R2278_U15 & P2_R2278_U17 & P2_U3637); 
assign P2_R2278_U513 = ~(P2_U2805 & P2_R2278_U60); 
assign P2_R2278_U515 = ~(P2_U2805 & P2_R2278_U60); 
assign P2_R2278_U519 = ~(P2_R2278_U43 & P2_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P2_R2278_U521 = ~(P2_R2278_U43 & P2_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P2_R2278_U530 = ~(P2_R2278_U529 & P2_R2278_U528); 
assign P2_ADD_394_U81 = ~(P2_ADD_394_U164 & P2_ADD_394_U163); 
assign P2_ADD_394_U118 = ~P2_ADD_394_U48; 
assign P2_ADD_394_U133 = ~(P2_ADD_394_U48 & P2_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P2_R2267_U79 = P2_R2267_U158 & P2_R2267_U157; 
assign P2_R2267_U106 = ~P2_R2267_U35; 
assign P2_R2267_U125 = ~(P2_U2778 & P2_R2267_U124); 
assign P2_R2267_U153 = ~(P2_U2777 & P2_R2267_U35); 
assign P2_ADD_371_1212_U139 = ~(P2_ADD_371_1212_U138 & P2_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P2_ADD_371_1212_U204 = ~(P2_ADD_371_1212_U136 & P2_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P2_ADD_371_1212_U220 = ~(P2_ADD_371_1212_U31 & P2_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P2_ADD_371_1212_U222 = ~(P2_ADD_371_1212_U31 & P2_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P1_R2278_U42 = ~(P1_R2278_U246 & P1_R2278_U245); 
assign P1_R2278_U138 = P1_R2278_U389 & P1_R2278_U276; 
assign P1_R2278_U140 = P1_R2278_U281 & P1_R2278_U283 & P1_R2278_U284; 
assign P1_R2278_U142 = P1_R2278_U7 & P1_R2278_U13; 
assign P1_R2278_U147 = P1_R2278_U324 & P1_R2278_U5; 
assign P1_R2278_U153 = P1_R2278_U7 & P1_R2278_U13; 
assign P1_R2278_U158 = P1_R2278_U7 & P1_R2278_U13; 
assign P1_R2278_U161 = P1_R2278_U9 & P1_R2278_U7; 
assign P1_R2278_U163 = P1_R2278_U73 & P1_R2278_U80; 
assign P1_R2278_U165 = P1_R2278_U371 & P1_R2278_U316; 
assign P1_R2278_U169 = P1_R2278_U362 & P1_R2278_U79; 
assign P1_R2278_U170 = P1_R2278_U367 & P1_R2278_U306; 
assign P1_R2278_U188 = P1_R2278_U470 & P1_R2278_U469; 
assign P1_R2278_U348 = ~(P1_R2278_U338 & P1_R2278_U285); 
assign P1_R2278_U349 = ~(P1_R2278_U339 & P1_R2278_U229); 
assign P1_R2278_U356 = ~(P1_R2278_U284 & P1_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P1_R2278_U368 = ~(P1_R2278_U367 & P1_R2278_U306); 
assign P1_R2278_U372 = ~(P1_R2278_U131 & P1_R2278_U371); 
assign P1_R2278_U377 = ~P1_R2278_U80; 
assign P1_R2278_U378 = ~P1_R2278_U73; 
assign P1_R2278_U383 = ~P1_R2278_U92; 
assign P1_R2278_U391 = ~(P1_R2278_U282 & P1_R2278_U283); 
assign P1_R2278_U392 = ~P1_R2278_U86; 
assign P1_R2278_U400 = ~(P1_R2278_U86 & P1_R2278_U324); 
assign P1_R2278_U454 = ~(P1_R2278_U243 & P1_R2278_U452); 
assign P1_R2278_U468 = ~(P1_R2278_U325 & P1_R2278_U5); 
assign P1_R2278_U591 = ~(P1_R2278_U67 & P1_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P1_R2278_U596 = ~(P1_R2278_U65 & P1_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P1_R2358_U70 = ~(P1_R2358_U358 & P1_R2358_U275); 
assign P1_R2358_U84 = ~(P1_R2358_U456 & P1_R2358_U455); 
assign P1_R2358_U108 = P1_R2358_U47 & P1_R2358_U278; 
assign P1_R2358_U128 = P1_R2358_U276 & P1_R2358_U5; 
assign P1_R2358_U142 = P1_R2358_U326 & P1_R2358_U263; 
assign P1_R2358_U167 = ~P1_U2661; 
assign P1_R2358_U227 = ~P1_R2358_U154; 
assign P1_R2358_U230 = ~(P1_R2358_U229 & P1_R2358_U154); 
assign P1_R2358_U235 = ~P1_R2358_U155; 
assign P1_R2358_U236 = ~(P1_R2358_U155 & P1_R2358_U219); 
assign P1_R2358_U255 = ~(P1_R2358_U460 & P1_R2358_U459 & P1_R2358_U60); 
assign P1_R2358_U258 = ~(P1_R2358_U468 & P1_R2358_U467 & P1_R2358_U58); 
assign P1_R2358_U260 = ~P1_R2358_U59; 
assign P1_R2358_U261 = ~P1_R2358_U61; 
assign P1_R2358_U268 = ~(P1_R2358_U124 & P1_R2358_U154 & P1_R2358_U125); 
assign P1_R2358_U279 = ~P1_R2358_U47; 
assign P1_R2358_U280 = ~(P1_R2358_U509 & P1_R2358_U508 & P1_R2358_U45); 
assign P1_R2358_U347 = ~(P1_R2358_U47 & P1_R2358_U278); 
assign P1_R2358_U357 = ~(P1_R2358_U232 & P1_R2358_U263); 
assign P1_R2358_U451 = ~(P1_R2358_U333 & P1_R2358_U154); 
assign P1_R2358_U453 = ~(P1_R2358_U334 & P1_R2358_U155); 
assign P1_R2358_U505 = ~(P1_U2661 & P1_R2358_U23); 
assign P1_R2358_U514 = ~(P1_U2661 & P1_R2358_U23); 
assign P1_R2358_U518 = ~(P1_R2358_U517 & P1_R2358_U516); 
assign P1_R2099_U73 = ~(P1_R2099_U313 & P1_R2099_U312); 
assign P1_R2099_U174 = ~P1_R2099_U19; 
assign P1_R2099_U311 = ~(P1_R2099_U50 & P1_R2099_U19); 
assign P1_R2337_U78 = ~(P1_R2337_U156 & P1_R2337_U155); 
assign P1_R2337_U115 = ~P1_R2337_U48; 
assign P1_R2337_U153 = ~(P1_R2337_U48 & P1_PHYADDRPOINTER_REG_24__SCAN_IN); 
assign P1_R2096_U78 = ~(P1_R2096_U156 & P1_R2096_U155); 
assign P1_R2096_U115 = ~P1_R2096_U48; 
assign P1_R2096_U153 = ~(P1_R2096_U48 & P1_REIP_REG_24__SCAN_IN); 
assign P1_ADD_405_U81 = ~(P1_ADD_405_U164 & P1_ADD_405_U163); 
assign P1_ADD_405_U118 = ~P1_ADD_405_U48; 
assign P1_ADD_405_U133 = ~(P1_ADD_405_U48 & P1_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P1_ADD_515_U81 = ~(P1_ADD_515_U162 & P1_ADD_515_U161); 
assign P1_ADD_515_U115 = ~P1_ADD_515_U48; 
assign P1_ADD_515_U129 = ~(P1_ADD_515_U48 & P1_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_U2844 = ~(P3_U6087 & P3_U6085 & P3_U6086); 
assign P3_U2997 = ~(P3_U4636 & P3_U4635 & P3_U4634 & P3_U4329); 
assign P3_U3282 = ~(P3_U7955 & P3_U7954); 
assign P3_U3841 = P3_U6114 & P3_U3838 & P3_U3840 & P3_U6112 & P3_U3844; 
assign P3_U3852 = P3_U3850 & P3_U3851 & P3_U6155; 
assign P3_U3975 = P3_U6580 & P3_U6577 & P3_U6578 & P3_U6579; 
assign P3_U6110 = ~(P3_U4318 & P3_U6108); 
assign P3_U6162 = ~(P3_ADD_558_U82 & P3_U3220); 
assign P3_U6163 = ~(P3_ADD_553_U82 & P3_U4298); 
assign P3_U6164 = ~(P3_ADD_547_U82 & P3_U4299); 
assign P3_U6167 = ~(P3_ADD_531_U82 & P3_U2354); 
assign P3_U6175 = ~(P3_ADD_385_U82 & P3_U2358); 
assign P3_U6176 = ~(P3_ADD_380_U82 & P3_U2359); 
assign P3_U6177 = ~(P3_ADD_349_U82 & P3_U4306); 
assign P3_U6178 = ~(P3_ADD_344_U82 & P3_U2362); 
assign P3_U6179 = ~(P3_ADD_371_1212_U82 & P3_U2360); 
assign P3_U6189 = ~(P3_ADD_541_U78 & P3_U4300); 
assign P3_U6190 = ~(P3_ADD_536_U78 & P3_U4301); 
assign P3_U6193 = ~(P3_ADD_515_U78 & P3_U4302); 
assign P3_U6194 = ~(P3_ADD_494_U78 & P3_U2356); 
assign P3_U6195 = ~(P3_ADD_476_U78 & P3_U4303); 
assign P3_U6196 = ~(P3_ADD_441_U78 & P3_U4304); 
assign P3_U6197 = ~(P3_ADD_405_U77 & P3_U4305); 
assign P3_U6198 = ~(P3_ADD_394_U77 & P3_U2357); 
assign P3_U6587 = ~(P3_U2387 & P3_ADD_371_1212_U82); 
assign P3_U6589 = ~(P3_ADD_318_U78 & P3_U2398); 
assign P3_U6594 = ~(P3_ADD_339_U78 & P3_U2388); 
assign P3_U6598 = ~(P3_ADD_315_U74 & P3_U2397); 
assign P3_U7294 = ~(P3_ADD_467_U78 & P3_U2601); 
assign P3_U7296 = ~(P3_ADD_430_U78 & P3_U2405); 
assign P2_U2803 = P2_U3242 & P2_R2267_U79; 
assign P2_U2875 = ~(P2_U6508 & P2_U6509 & P2_U6507); 
assign P2_U2913 = ~(P2_U6352 & P2_U6351 & P2_U4065); 
assign P2_U4112 = P2_U6675 & P2_U4446 & P2_U6678; 
assign P2_U4129 = P2_U6715 & P2_U4446; 
assign P2_U4672 = ~(P2_U2406 & P2_U4668); 
assign P2_U4673 = ~(P2_U4663 & P2_INSTQUEUE_REG_15__7__SCAN_IN); 
assign P2_U4677 = ~(P2_U2405 & P2_U4668); 
assign P2_U4678 = ~(P2_U4663 & P2_INSTQUEUE_REG_15__6__SCAN_IN); 
assign P2_U4682 = ~(P2_U2404 & P2_U4668); 
assign P2_U4683 = ~(P2_U4663 & P2_INSTQUEUE_REG_15__5__SCAN_IN); 
assign P2_U4687 = ~(P2_U2403 & P2_U4668); 
assign P2_U4688 = ~(P2_U4663 & P2_INSTQUEUE_REG_15__4__SCAN_IN); 
assign P2_U4692 = ~(P2_U2402 & P2_U4668); 
assign P2_U4693 = ~(P2_U4663 & P2_INSTQUEUE_REG_15__3__SCAN_IN); 
assign P2_U4697 = ~(P2_U2401 & P2_U4668); 
assign P2_U4698 = ~(P2_U4663 & P2_INSTQUEUE_REG_15__2__SCAN_IN); 
assign P2_U4702 = ~(P2_U2400 & P2_U4668); 
assign P2_U4703 = ~(P2_U4663 & P2_INSTQUEUE_REG_15__1__SCAN_IN); 
assign P2_U4707 = ~(P2_U2399 & P2_U4668); 
assign P2_U4708 = ~(P2_U4663 & P2_INSTQUEUE_REG_15__0__SCAN_IN); 
assign P2_U4730 = ~(P2_U2406 & P2_U4726); 
assign P2_U4731 = ~(P2_U4721 & P2_INSTQUEUE_REG_14__7__SCAN_IN); 
assign P2_U4735 = ~(P2_U2405 & P2_U4726); 
assign P2_U4736 = ~(P2_U4721 & P2_INSTQUEUE_REG_14__6__SCAN_IN); 
assign P2_U4740 = ~(P2_U2404 & P2_U4726); 
assign P2_U4741 = ~(P2_U4721 & P2_INSTQUEUE_REG_14__5__SCAN_IN); 
assign P2_U4745 = ~(P2_U2403 & P2_U4726); 
assign P2_U4746 = ~(P2_U4721 & P2_INSTQUEUE_REG_14__4__SCAN_IN); 
assign P2_U4750 = ~(P2_U2402 & P2_U4726); 
assign P2_U4751 = ~(P2_U4721 & P2_INSTQUEUE_REG_14__3__SCAN_IN); 
assign P2_U4755 = ~(P2_U2401 & P2_U4726); 
assign P2_U4756 = ~(P2_U4721 & P2_INSTQUEUE_REG_14__2__SCAN_IN); 
assign P2_U4760 = ~(P2_U2400 & P2_U4726); 
assign P2_U4761 = ~(P2_U4721 & P2_INSTQUEUE_REG_14__1__SCAN_IN); 
assign P2_U4765 = ~(P2_U2399 & P2_U4726); 
assign P2_U4766 = ~(P2_U4721 & P2_INSTQUEUE_REG_14__0__SCAN_IN); 
assign P2_U4789 = ~(P2_U2406 & P2_U4785); 
assign P2_U4790 = ~(P2_U4780 & P2_INSTQUEUE_REG_13__7__SCAN_IN); 
assign P2_U4794 = ~(P2_U2405 & P2_U4785); 
assign P2_U4795 = ~(P2_U4780 & P2_INSTQUEUE_REG_13__6__SCAN_IN); 
assign P2_U4799 = ~(P2_U2404 & P2_U4785); 
assign P2_U4800 = ~(P2_U4780 & P2_INSTQUEUE_REG_13__5__SCAN_IN); 
assign P2_U4804 = ~(P2_U2403 & P2_U4785); 
assign P2_U4805 = ~(P2_U4780 & P2_INSTQUEUE_REG_13__4__SCAN_IN); 
assign P2_U4809 = ~(P2_U2402 & P2_U4785); 
assign P2_U4810 = ~(P2_U4780 & P2_INSTQUEUE_REG_13__3__SCAN_IN); 
assign P2_U4814 = ~(P2_U2401 & P2_U4785); 
assign P2_U4815 = ~(P2_U4780 & P2_INSTQUEUE_REG_13__2__SCAN_IN); 
assign P2_U4819 = ~(P2_U2400 & P2_U4785); 
assign P2_U4820 = ~(P2_U4780 & P2_INSTQUEUE_REG_13__1__SCAN_IN); 
assign P2_U4824 = ~(P2_U2399 & P2_U4785); 
assign P2_U4825 = ~(P2_U4780 & P2_INSTQUEUE_REG_13__0__SCAN_IN); 
assign P2_U4846 = ~(P2_U2406 & P2_U4842); 
assign P2_U4847 = ~(P2_U4837 & P2_INSTQUEUE_REG_12__7__SCAN_IN); 
assign P2_U4851 = ~(P2_U2405 & P2_U4842); 
assign P2_U4852 = ~(P2_U4837 & P2_INSTQUEUE_REG_12__6__SCAN_IN); 
assign P2_U4856 = ~(P2_U2404 & P2_U4842); 
assign P2_U4857 = ~(P2_U4837 & P2_INSTQUEUE_REG_12__5__SCAN_IN); 
assign P2_U4861 = ~(P2_U2403 & P2_U4842); 
assign P2_U4862 = ~(P2_U4837 & P2_INSTQUEUE_REG_12__4__SCAN_IN); 
assign P2_U4866 = ~(P2_U2402 & P2_U4842); 
assign P2_U4867 = ~(P2_U4837 & P2_INSTQUEUE_REG_12__3__SCAN_IN); 
assign P2_U4871 = ~(P2_U2401 & P2_U4842); 
assign P2_U4872 = ~(P2_U4837 & P2_INSTQUEUE_REG_12__2__SCAN_IN); 
assign P2_U4876 = ~(P2_U2400 & P2_U4842); 
assign P2_U4877 = ~(P2_U4837 & P2_INSTQUEUE_REG_12__1__SCAN_IN); 
assign P2_U4881 = ~(P2_U2399 & P2_U4842); 
assign P2_U4882 = ~(P2_U4837 & P2_INSTQUEUE_REG_12__0__SCAN_IN); 
assign P2_U4904 = ~(P2_U2406 & P2_U4900); 
assign P2_U4905 = ~(P2_U4895 & P2_INSTQUEUE_REG_11__7__SCAN_IN); 
assign P2_U4909 = ~(P2_U2405 & P2_U4900); 
assign P2_U4910 = ~(P2_U4895 & P2_INSTQUEUE_REG_11__6__SCAN_IN); 
assign P2_U4914 = ~(P2_U2404 & P2_U4900); 
assign P2_U4915 = ~(P2_U4895 & P2_INSTQUEUE_REG_11__5__SCAN_IN); 
assign P2_U4919 = ~(P2_U2403 & P2_U4900); 
assign P2_U4920 = ~(P2_U4895 & P2_INSTQUEUE_REG_11__4__SCAN_IN); 
assign P2_U4924 = ~(P2_U2402 & P2_U4900); 
assign P2_U4925 = ~(P2_U4895 & P2_INSTQUEUE_REG_11__3__SCAN_IN); 
assign P2_U4929 = ~(P2_U2401 & P2_U4900); 
assign P2_U4930 = ~(P2_U4895 & P2_INSTQUEUE_REG_11__2__SCAN_IN); 
assign P2_U4934 = ~(P2_U2400 & P2_U4900); 
assign P2_U4935 = ~(P2_U4895 & P2_INSTQUEUE_REG_11__1__SCAN_IN); 
assign P2_U4939 = ~(P2_U2399 & P2_U4900); 
assign P2_U4940 = ~(P2_U4895 & P2_INSTQUEUE_REG_11__0__SCAN_IN); 
assign P2_U4961 = ~(P2_U2406 & P2_U4957); 
assign P2_U4962 = ~(P2_U4952 & P2_INSTQUEUE_REG_10__7__SCAN_IN); 
assign P2_U4966 = ~(P2_U2405 & P2_U4957); 
assign P2_U4967 = ~(P2_U4952 & P2_INSTQUEUE_REG_10__6__SCAN_IN); 
assign P2_U4971 = ~(P2_U2404 & P2_U4957); 
assign P2_U4972 = ~(P2_U4952 & P2_INSTQUEUE_REG_10__5__SCAN_IN); 
assign P2_U4976 = ~(P2_U2403 & P2_U4957); 
assign P2_U4977 = ~(P2_U4952 & P2_INSTQUEUE_REG_10__4__SCAN_IN); 
assign P2_U4981 = ~(P2_U2402 & P2_U4957); 
assign P2_U4982 = ~(P2_U4952 & P2_INSTQUEUE_REG_10__3__SCAN_IN); 
assign P2_U4986 = ~(P2_U2401 & P2_U4957); 
assign P2_U4987 = ~(P2_U4952 & P2_INSTQUEUE_REG_10__2__SCAN_IN); 
assign P2_U4991 = ~(P2_U2400 & P2_U4957); 
assign P2_U4992 = ~(P2_U4952 & P2_INSTQUEUE_REG_10__1__SCAN_IN); 
assign P2_U4996 = ~(P2_U2399 & P2_U4957); 
assign P2_U4997 = ~(P2_U4952 & P2_INSTQUEUE_REG_10__0__SCAN_IN); 
assign P2_U5019 = ~(P2_U2406 & P2_U5015); 
assign P2_U5020 = ~(P2_U5010 & P2_INSTQUEUE_REG_9__7__SCAN_IN); 
assign P2_U5024 = ~(P2_U2405 & P2_U5015); 
assign P2_U5025 = ~(P2_U5010 & P2_INSTQUEUE_REG_9__6__SCAN_IN); 
assign P2_U5029 = ~(P2_U2404 & P2_U5015); 
assign P2_U5030 = ~(P2_U5010 & P2_INSTQUEUE_REG_9__5__SCAN_IN); 
assign P2_U5034 = ~(P2_U2403 & P2_U5015); 
assign P2_U5035 = ~(P2_U5010 & P2_INSTQUEUE_REG_9__4__SCAN_IN); 
assign P2_U5039 = ~(P2_U2402 & P2_U5015); 
assign P2_U5040 = ~(P2_U5010 & P2_INSTQUEUE_REG_9__3__SCAN_IN); 
assign P2_U5044 = ~(P2_U2401 & P2_U5015); 
assign P2_U5045 = ~(P2_U5010 & P2_INSTQUEUE_REG_9__2__SCAN_IN); 
assign P2_U5049 = ~(P2_U2400 & P2_U5015); 
assign P2_U5050 = ~(P2_U5010 & P2_INSTQUEUE_REG_9__1__SCAN_IN); 
assign P2_U5054 = ~(P2_U2399 & P2_U5015); 
assign P2_U5055 = ~(P2_U5010 & P2_INSTQUEUE_REG_9__0__SCAN_IN); 
assign P2_U5076 = ~(P2_U2406 & P2_U5072); 
assign P2_U5077 = ~(P2_U5067 & P2_INSTQUEUE_REG_8__7__SCAN_IN); 
assign P2_U5081 = ~(P2_U2405 & P2_U5072); 
assign P2_U5082 = ~(P2_U5067 & P2_INSTQUEUE_REG_8__6__SCAN_IN); 
assign P2_U5086 = ~(P2_U2404 & P2_U5072); 
assign P2_U5087 = ~(P2_U5067 & P2_INSTQUEUE_REG_8__5__SCAN_IN); 
assign P2_U5091 = ~(P2_U2403 & P2_U5072); 
assign P2_U5092 = ~(P2_U5067 & P2_INSTQUEUE_REG_8__4__SCAN_IN); 
assign P2_U5096 = ~(P2_U2402 & P2_U5072); 
assign P2_U5097 = ~(P2_U5067 & P2_INSTQUEUE_REG_8__3__SCAN_IN); 
assign P2_U5101 = ~(P2_U2401 & P2_U5072); 
assign P2_U5102 = ~(P2_U5067 & P2_INSTQUEUE_REG_8__2__SCAN_IN); 
assign P2_U5106 = ~(P2_U2400 & P2_U5072); 
assign P2_U5107 = ~(P2_U5067 & P2_INSTQUEUE_REG_8__1__SCAN_IN); 
assign P2_U5111 = ~(P2_U2399 & P2_U5072); 
assign P2_U5112 = ~(P2_U5067 & P2_INSTQUEUE_REG_8__0__SCAN_IN); 
assign P2_U5123 = ~(P2_U5120 & P2_U3794); 
assign P2_U5128 = ~(P2_U5127 & P2_U5126); 
assign P2_U5180 = ~(P2_U5177 & P2_U3803); 
assign P2_U5185 = ~(P2_U5184 & P2_U5183); 
assign P2_U5238 = ~(P2_U5235 & P2_U3812); 
assign P2_U5243 = ~(P2_U5242 & P2_U5241); 
assign P2_U5295 = ~(P2_U5292 & P2_U3821); 
assign P2_U5300 = ~(P2_U5299 & P2_U5298); 
assign P2_U5353 = ~(P2_U5350 & P2_U3830); 
assign P2_U5358 = ~(P2_U5357 & P2_U5356); 
assign P2_U5410 = ~(P2_U5407 & P2_U3839); 
assign P2_U5415 = ~(P2_U5414 & P2_U5413); 
assign P2_U5468 = ~(P2_U5465 & P2_U3848); 
assign P2_U5473 = ~(P2_U5472 & P2_U5471); 
assign P2_U5525 = ~(P2_U5522 & P2_U3857); 
assign P2_U5530 = ~(P2_U5529 & P2_U5528); 
assign P2_U6414 = ~(P2_U2380 & P2_R2096_U87); 
assign P2_U6510 = ~(P2_R2182_U93 & P2_U2393); 
assign P2_U6723 = ~(P2_R2267_U79 & P2_U2587); 
assign P2_U6740 = ~(P2_U2588 & P2_R2096_U87); 
assign P2_U8323 = ~(P2_R2256_U26 & P2_U3572); 
assign P2_U8387 = ~(P2_R2337_U76 & P2_U3284); 
assign P1_U2660 = ~(P1_U6808 & P1_U4018); 
assign P1_U2996 = ~(P1_U5816 & P1_U5814 & P1_U5815 & P1_U5818 & P1_U5817); 
assign P1_U3161 = ~(P1_U7690 & P1_U7689 & P1_U3586); 
assign P1_U3163 = ~(P1_U3582 & P1_U4516); 
assign P1_U3660 = P1_U5021 & P1_U5020 & P1_U5022; 
assign P1_U3661 = P1_U5026 & P1_U5025 & P1_U5027; 
assign P1_U3662 = P1_U5031 & P1_U5030 & P1_U5032; 
assign P1_U3663 = P1_U5036 & P1_U5035 & P1_U5037; 
assign P1_U3664 = P1_U5041 & P1_U5040 & P1_U5042; 
assign P1_U3665 = P1_U5046 & P1_U5045 & P1_U5047; 
assign P1_U3666 = P1_U5051 & P1_U5050 & P1_U5052; 
assign P1_U3667 = P1_U5056 & P1_U5055 & P1_U5057; 
assign P1_U3669 = P1_U5078 & P1_U5077 & P1_U5079; 
assign P1_U3670 = P1_U5083 & P1_U5082 & P1_U5084; 
assign P1_U3671 = P1_U5088 & P1_U5087 & P1_U5089; 
assign P1_U3672 = P1_U5093 & P1_U5092 & P1_U5094; 
assign P1_U3673 = P1_U5098 & P1_U5097 & P1_U5099; 
assign P1_U3674 = P1_U5103 & P1_U5102 & P1_U5104; 
assign P1_U3675 = P1_U5108 & P1_U5107 & P1_U5109; 
assign P1_U3676 = P1_U5113 & P1_U5112 & P1_U5114; 
assign P1_U3678 = P1_U5136 & P1_U5135 & P1_U5137; 
assign P1_U3679 = P1_U5141 & P1_U5140 & P1_U5142; 
assign P1_U3680 = P1_U5146 & P1_U5145 & P1_U5147; 
assign P1_U3681 = P1_U5151 & P1_U5150 & P1_U5152; 
assign P1_U3682 = P1_U5156 & P1_U5155 & P1_U5157; 
assign P1_U3683 = P1_U5161 & P1_U5160 & P1_U5162; 
assign P1_U3684 = P1_U5166 & P1_U5165 & P1_U5167; 
assign P1_U3685 = P1_U5171 & P1_U5170 & P1_U5172; 
assign P1_U3687 = P1_U5193 & P1_U5192 & P1_U5194; 
assign P1_U3688 = P1_U5198 & P1_U5197 & P1_U5199; 
assign P1_U3689 = P1_U5203 & P1_U5202 & P1_U5204; 
assign P1_U3690 = P1_U5208 & P1_U5207 & P1_U5209; 
assign P1_U3691 = P1_U5213 & P1_U5212 & P1_U5214; 
assign P1_U3692 = P1_U5218 & P1_U5217 & P1_U5219; 
assign P1_U3693 = P1_U5223 & P1_U5222 & P1_U5224; 
assign P1_U3694 = P1_U5228 & P1_U5227 & P1_U5229; 
assign P1_U3696 = P1_U5251 & P1_U5250 & P1_U5252; 
assign P1_U3697 = P1_U5256 & P1_U5255 & P1_U5257; 
assign P1_U3698 = P1_U5261 & P1_U5260 & P1_U5262; 
assign P1_U3699 = P1_U5266 & P1_U5265 & P1_U5267; 
assign P1_U3700 = P1_U5271 & P1_U5270 & P1_U5272; 
assign P1_U3701 = P1_U5276 & P1_U5275 & P1_U5277; 
assign P1_U3702 = P1_U5281 & P1_U5280 & P1_U5282; 
assign P1_U3703 = P1_U5286 & P1_U5285 & P1_U5287; 
assign P1_U3705 = P1_U5308 & P1_U5307 & P1_U5309; 
assign P1_U3706 = P1_U5313 & P1_U5312 & P1_U5314; 
assign P1_U3707 = P1_U5318 & P1_U5317 & P1_U5319; 
assign P1_U3708 = P1_U5323 & P1_U5322 & P1_U5324; 
assign P1_U3709 = P1_U5328 & P1_U5327 & P1_U5329; 
assign P1_U3710 = P1_U5333 & P1_U5332 & P1_U5334; 
assign P1_U3711 = P1_U5338 & P1_U5337 & P1_U5339; 
assign P1_U3712 = P1_U5343 & P1_U5342 & P1_U5344; 
assign P1_U3714 = P1_U5366 & P1_U5365 & P1_U5367; 
assign P1_U3715 = P1_U5371 & P1_U5370 & P1_U5372; 
assign P1_U3716 = P1_U5376 & P1_U5375 & P1_U5377; 
assign P1_U3717 = P1_U5381 & P1_U5380 & P1_U5382; 
assign P1_U3718 = P1_U5386 & P1_U5385 & P1_U5387; 
assign P1_U3719 = P1_U5391 & P1_U5390 & P1_U5392; 
assign P1_U3720 = P1_U5396 & P1_U5395 & P1_U5397; 
assign P1_U3721 = P1_U5401 & P1_U5400 & P1_U5402; 
assign P1_U3723 = P1_U5423 & P1_U5422 & P1_U5424; 
assign P1_U3724 = P1_U5428 & P1_U5427 & P1_U5429; 
assign P1_U3725 = P1_U5433 & P1_U5432 & P1_U5434; 
assign P1_U3726 = P1_U5438 & P1_U5437 & P1_U5439; 
assign P1_U3727 = P1_U5442 & P1_U5441 & P1_U5443; 
assign P1_U3728 = P1_U5447 & P1_U5446 & P1_U5448; 
assign P1_U3729 = P1_U5452 & P1_U5451 & P1_U5453; 
assign P1_U3730 = P1_U5457 & P1_U5456 & P1_U5458; 
assign P1_U3776 = P1_U3777 & P1_U5595 & P1_U5593; 
assign P1_U4518 = ~(P1_U3583 & P1_U4514); 
assign P1_U4551 = ~(P1_U4536 & P1_U4550); 
assign P1_U4557 = ~(P1_U4556 & P1_U3321); 
assign P1_U4609 = ~(P1_U4604 & P1_U4608); 
assign P1_U4615 = ~(P1_U4614 & P1_U3328); 
assign P1_U4668 = ~(P1_U4662 & P1_U4667); 
assign P1_U4674 = ~(P1_U4673 & P1_U3335); 
assign P1_U4725 = ~(P1_U4720 & P1_U4724); 
assign P1_U4731 = ~(P1_U4730 & P1_U3339); 
assign P1_U4783 = ~(P1_U4777 & P1_U4782); 
assign P1_U4789 = ~(P1_U4788 & P1_U3344); 
assign P1_U4840 = ~(P1_U4835 & P1_U4839); 
assign P1_U4846 = ~(P1_U4845 & P1_U3348); 
assign P1_U4898 = ~(P1_U4892 & P1_U4897); 
assign P1_U4904 = ~(P1_U4903 & P1_U3351); 
assign P1_U4955 = ~(P1_U4950 & P1_U4954); 
assign P1_U4961 = ~(P1_U4960 & P1_U3355); 
assign P1_U5010 = ~(P1_U3320 & P1_U5009); 
assign P1_U5016 = ~(P1_U3320 & P1_U5015); 
assign P1_U5067 = ~(P1_U3320 & P1_U5066); 
assign P1_U5073 = ~(P1_U3320 & P1_U5072); 
assign P1_U5125 = ~(P1_U3320 & P1_U5124); 
assign P1_U5131 = ~(P1_U3320 & P1_U5130); 
assign P1_U5182 = ~(P1_U3320 & P1_U5181); 
assign P1_U5188 = ~(P1_U3320 & P1_U5187); 
assign P1_U5240 = ~(P1_U3320 & P1_U5239); 
assign P1_U5246 = ~(P1_U3320 & P1_U5245); 
assign P1_U5297 = ~(P1_U3320 & P1_U5296); 
assign P1_U5303 = ~(P1_U3320 & P1_U5302); 
assign P1_U5355 = ~(P1_U3320 & P1_U5354); 
assign P1_U5361 = ~(P1_U3320 & P1_U5360); 
assign P1_U5412 = ~(P1_U3320 & P1_U5411); 
assign P1_U5418 = ~(P1_U3320 & P1_U5417); 
assign P1_U5545 = ~(P1_U3751 & P1_U5542); 
assign P1_U5724 = ~(P1_R2099_U73 & P1_U2380); 
assign P1_U5734 = ~(P1_ADD_405_U81 & P1_U2375); 
assign P1_U5735 = ~(P1_ADD_515_U81 & P1_U2374); 
assign P1_U5822 = ~(P1_R2358_U84 & P1_U2364); 
assign P1_U5914 = ~(P1_R2337_U78 & P1_U2376); 
assign P1_U6167 = ~(P1_U2386 & P1_R2358_U84); 
assign P1_U6277 = ~(P1_U2383 & P1_R2358_U84); 
assign P1_U6332 = ~(P1_U2371 & P1_R2099_U73); 
assign P1_U6528 = ~(P1_U2604 & P1_R2099_U73); 
assign P1_U6536 = ~(P1_R2096_U78 & P1_U7485); 
assign P1_U6807 = ~(P1_R2337_U78 & P1_U2352); 
assign P1_U7686 = ~(P1_U2428 & P1_U4514); 
assign P3_ADD_476_U50 = ~(P3_ADD_476_U115 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_476_U154 = ~(P3_ADD_476_U115 & P3_ADD_476_U49); 
assign P3_ADD_531_U51 = ~(P3_ADD_531_U119 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_531_U161 = ~(P3_ADD_531_U119 & P3_ADD_531_U50); 
assign P3_SUB_320_U12 = P3_SUB_320_U114 & P3_SUB_320_U34; 
assign P3_SUB_320_U67 = ~P3_ADD_318_U78; 
assign P3_SUB_320_U99 = ~P3_SUB_320_U34; 
assign P3_SUB_320_U144 = ~(P3_ADD_318_U78 & P3_SUB_320_U34); 
assign P3_ADD_318_U50 = ~(P3_ADD_318_U115 & P3_PHYADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_318_U154 = ~(P3_ADD_318_U115 & P3_ADD_318_U49); 
assign P3_ADD_315_U50 = ~(P3_ADD_315_U112 & P3_PHYADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_315_U146 = ~(P3_ADD_315_U112 & P3_ADD_315_U49); 
assign P3_ADD_360_1242_U80 = ~(P3_ADD_360_1242_U243 & P3_ADD_360_1242_U242); 
assign P3_ADD_360_1242_U161 = ~P3_ADD_360_1242_U63; 
assign P3_ADD_360_1242_U173 = ~(P3_ADD_360_1242_U61 & P3_ADD_360_1242_U172); 
assign P3_ADD_360_1242_U240 = ~(P3_ADD_360_1242_U63 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_467_U50 = ~(P3_ADD_467_U115 & P3_REIP_REG_24__SCAN_IN); 
assign P3_ADD_467_U154 = ~(P3_ADD_467_U115 & P3_ADD_467_U49); 
assign P3_ADD_430_U50 = ~(P3_ADD_430_U115 & P3_REIP_REG_24__SCAN_IN); 
assign P3_ADD_430_U154 = ~(P3_ADD_430_U115 & P3_ADD_430_U49); 
assign P3_ADD_380_U51 = ~(P3_ADD_380_U119 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_380_U161 = ~(P3_ADD_380_U119 & P3_ADD_380_U50); 
assign P3_ADD_344_U51 = ~(P3_ADD_344_U119 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_344_U161 = ~(P3_ADD_344_U119 & P3_ADD_344_U50); 
assign P3_ADD_339_U50 = ~(P3_ADD_339_U115 & P3_PHYADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_339_U154 = ~(P3_ADD_339_U115 & P3_ADD_339_U49); 
assign P3_ADD_541_U50 = ~(P3_ADD_541_U115 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_541_U154 = ~(P3_ADD_541_U115 & P3_ADD_541_U49); 
assign P3_SUB_357_1258_U17 = P3_SUB_357_1258_U244 & P3_SUB_357_1258_U241; 
assign P3_SUB_357_1258_U19 = P3_SUB_357_1258_U227 & P3_SUB_357_1258_U303; 
assign P3_SUB_357_1258_U79 = ~(P3_SUB_357_1258_U373 & P3_SUB_357_1258_U372); 
assign P3_SUB_357_1258_U85 = ~(P3_SUB_357_1258_U419 & P3_SUB_357_1258_U418); 
assign P3_SUB_357_1258_U223 = ~P3_SUB_357_1258_U61; 
assign P3_SUB_357_1258_U295 = ~(P3_SUB_357_1258_U61 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_SUB_357_1258_U297 = ~(P3_SUB_357_1258_U108 & P3_SUB_357_1258_U61); 
assign P3_SUB_357_1258_U352 = ~(P3_ADD_357_U6 & P3_SUB_357_1258_U224); 
assign P3_SUB_357_1258_U360 = ~(P3_SUB_357_1258_U126 & P3_SUB_357_1258_U61); 
assign P3_ADD_515_U50 = ~(P3_ADD_515_U115 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_515_U154 = ~(P3_ADD_515_U115 & P3_ADD_515_U49); 
assign P3_ADD_394_U50 = ~(P3_ADD_394_U118 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_394_U156 = ~(P3_ADD_394_U118 & P3_ADD_394_U49); 
assign P3_ADD_441_U50 = ~(P3_ADD_441_U115 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_441_U154 = ~(P3_ADD_441_U115 & P3_ADD_441_U49); 
assign P3_ADD_349_U51 = ~(P3_ADD_349_U119 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_349_U161 = ~(P3_ADD_349_U119 & P3_ADD_349_U50); 
assign P3_ADD_405_U50 = ~(P3_ADD_405_U118 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_405_U156 = ~(P3_ADD_405_U118 & P3_ADD_405_U49); 
assign P3_ADD_553_U51 = ~(P3_ADD_553_U119 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_553_U161 = ~(P3_ADD_553_U119 & P3_ADD_553_U50); 
assign P3_ADD_558_U51 = ~(P3_ADD_558_U119 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_558_U161 = ~(P3_ADD_558_U119 & P3_ADD_558_U50); 
assign P3_ADD_385_U51 = ~(P3_ADD_385_U119 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_385_U161 = ~(P3_ADD_385_U119 & P3_ADD_385_U50); 
assign P3_ADD_547_U51 = ~(P3_ADD_547_U119 & P3_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P3_ADD_547_U161 = ~(P3_ADD_547_U119 & P3_ADD_547_U50); 
assign P3_ADD_371_1212_U13 = P3_ADD_371_1212_U183 & P3_ADD_371_1212_U65; 
assign P3_ADD_371_1212_U68 = ~(P3_ADD_371_1212_U106 & P3_ADD_371_1212_U170); 
assign P3_ADD_371_1212_U180 = ~(P3_ADD_371_1212_U170 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_371_1212_U248 = ~(P3_ADD_371_1212_U170 & P3_ADD_371_1212_U67); 
assign P3_ADD_494_U50 = ~(P3_ADD_494_U115 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_494_U154 = ~(P3_ADD_494_U115 & P3_ADD_494_U49); 
assign P3_ADD_536_U50 = ~(P3_ADD_536_U115 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_536_U154 = ~(P3_ADD_536_U115 & P3_ADD_536_U49); 
assign P2_R2099_U90 = ~(P2_R2099_U217 & P2_R2099_U216); 
assign P2_R2099_U129 = ~P2_R2099_U33; 
assign P2_R2099_U214 = ~(P2_U2733 & P2_R2099_U33); 
assign P2_ADD_391_1196_U44 = ~P2_R2182_U93; 
assign P2_ADD_391_1196_U63 = ~P2_R2096_U87; 
assign P2_ADD_391_1196_U157 = P2_ADD_391_1196_U471 & P2_ADD_391_1196_U470; 
assign P2_ADD_391_1196_U187 = ~P2_ADD_391_1196_U112; 
assign P2_ADD_391_1196_U189 = ~(P2_ADD_391_1196_U188 & P2_ADD_391_1196_U112); 
assign P2_ADD_391_1196_U201 = ~(P2_ADD_391_1196_U185 & P2_ADD_391_1196_U200); 
assign P2_ADD_391_1196_U218 = P2_R2096_U94 | P2_R2182_U93; 
assign P2_ADD_391_1196_U220 = ~(P2_R2096_U94 & P2_R2182_U93); 
assign P2_ADD_391_1196_U295 = ~(P2_R2096_U94 & P2_R2182_U93); 
assign P2_ADD_391_1196_U314 = ~(P2_ADD_391_1196_U111 & P2_ADD_391_1196_U112); 
assign P2_ADD_391_1196_U462 = ~(P2_R2182_U93 & P2_ADD_391_1196_U45); 
assign P2_ADD_391_1196_U463 = ~(P2_R2096_U95 & P2_ADD_391_1196_U51); 
assign P2_ADD_391_1196_U465 = ~(P2_R2096_U95 & P2_ADD_391_1196_U51); 
assign P2_R2182_U17 = P2_U2696 & P2_R2182_U16; 
assign P2_R2182_U92 = ~(P2_R2182_U295 & P2_R2182_U294); 
assign P2_R2182_U147 = ~P2_R2182_U16; 
assign P2_R2182_U290 = ~(P2_R2182_U27 & P2_R2182_U16); 
assign P2_R2182_U293 = ~(P2_R2182_U146 & P2_U2666); 
assign P2_R2027_U51 = ~(P2_R2027_U119 & P2_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P2_R2027_U161 = ~(P2_R2027_U119 & P2_R2027_U50); 
assign P2_R2337_U51 = ~(P2_R2337_U116 & P2_PHYADDRPOINTER_REG_25__SCAN_IN); 
assign P2_R2337_U152 = ~(P2_R2337_U116 & P2_R2337_U50); 
assign P2_R2096_U10 = P2_U2626 & P2_R2096_U9; 
assign P2_R2096_U86 = ~(P2_R2096_U236 & P2_R2096_U235); 
assign P2_R2096_U158 = ~P2_R2096_U9; 
assign P2_R2096_U231 = ~(P2_R2096_U45 & P2_R2096_U9); 
assign P2_R2096_U234 = ~(P2_R2096_U157 & P2_U2627); 
assign P2_LT_563_U6 = P2_LT_563_U27 & P2_LT_563_U26; 
assign P2_R2256_U20 = ~(P2_R2256_U54 & P2_R2256_U53); 
assign P2_R2256_U42 = ~P2_R2256_U12; 
assign P2_R2256_U51 = ~(P2_U3624 & P2_R2256_U12); 
assign P2_R1957_U12 = P2_R1957_U114 & P2_R1957_U33; 
assign P2_R1957_U67 = ~P2_U3667; 
assign P2_R1957_U99 = ~P2_R1957_U33; 
assign P2_R1957_U144 = ~(P2_U3667 & P2_R1957_U33); 
assign P2_R2278_U18 = ~P2_U3636; 
assign P2_R2278_U20 = ~(P2_U3636 & P2_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P2_R2278_U41 = ~P2_U2804; 
assign P2_R2278_U126 = P2_R2278_U326 & P2_R2278_U257; 
assign P2_R2278_U165 = ~(P2_R2278_U310 & P2_R2278_U82 & P2_R2278_U311); 
assign P2_R2278_U193 = P2_R2278_U520 & P2_R2278_U519; 
assign P2_R2278_U207 = ~P2_R2278_U82; 
assign P2_R2278_U210 = P2_U3636 | P2_INSTADDRPOINTER_REG_2__SCAN_IN; 
assign P2_R2278_U261 = ~P2_R2278_U61; 
assign P2_R2278_U263 = P2_U2804 | P2_INSTADDRPOINTER_REG_17__SCAN_IN; 
assign P2_R2278_U264 = ~(P2_U2804 & P2_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P2_R2278_U410 = ~(P2_U3636 & P2_R2278_U19); 
assign P2_R2278_U412 = ~(P2_U3636 & P2_R2278_U19); 
assign P2_R2278_U490 = ~(P2_R2278_U488 & P2_R2278_U16); 
assign P2_R2278_U506 = ~(P2_U2804 & P2_R2278_U42); 
assign P2_R2278_U508 = ~(P2_U2804 & P2_R2278_U42); 
assign P2_R2278_U512 = ~(P2_R2278_U59 & P2_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P2_R2278_U514 = ~(P2_R2278_U59 & P2_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P2_R2278_U523 = ~(P2_R2278_U522 & P2_R2278_U521); 
assign P2_ADD_394_U50 = ~(P2_ADD_394_U118 & P2_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P2_ADD_394_U134 = ~(P2_ADD_394_U118 & P2_ADD_394_U49); 
assign P2_R2267_U10 = P2_R2267_U125 & P2_R2267_U35; 
assign P2_R2267_U36 = ~(P2_R2267_U50 & P2_R2267_U106); 
assign P2_R2267_U122 = ~(P2_R2267_U106 & P2_R2267_U74); 
assign P2_R2267_U154 = ~(P2_R2267_U106 & P2_R2267_U74); 
assign P2_ADD_371_1212_U25 = ~(P2_ADD_371_1212_U269 & P2_ADD_371_1212_U268 & P2_ADD_371_1212_U204); 
assign P2_ADD_371_1212_U33 = ~P2_R2256_U26; 
assign P2_ADD_371_1212_U115 = P2_ADD_371_1212_U221 & P2_ADD_371_1212_U220; 
assign P2_ADD_371_1212_U116 = ~(P2_ADD_371_1212_U67 & P2_ADD_371_1212_U139); 
assign P2_ADD_371_1212_U145 = P2_R2256_U26 | P2_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P2_ADD_371_1212_U147 = ~(P2_R2256_U26 & P2_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P2_ADD_371_1212_U224 = ~(P2_ADD_371_1212_U223 & P2_ADD_371_1212_U222); 
assign P2_ADD_371_1212_U259 = ~(P2_R2256_U26 & P2_ADD_371_1212_U34); 
assign P2_ADD_371_1212_U261 = ~(P2_R2256_U26 & P2_ADD_371_1212_U34); 
assign P1_R2278_U43 = ~(P1_R2278_U42 & P1_R2278_U248); 
assign P1_R2278_U63 = ~P1_U2785; 
assign P1_R2278_U93 = ~(P1_R2278_U11 & P1_R2278_U321 & P1_R2278_U377); 
assign P1_R2278_U94 = ~(P1_R2278_U132 & P1_R2278_U372); 
assign P1_R2278_U95 = ~(P1_R2278_U136 & P1_R2278_U368); 
assign P1_R2278_U96 = ~(P1_R2278_U11 & P1_R2278_U321 & P1_R2278_U378); 
assign P1_R2278_U104 = ~(P1_R2278_U454 & P1_R2278_U453); 
assign P1_R2278_U247 = ~P1_R2278_U42; 
assign P1_R2278_U286 = ~(P1_U2785 & P1_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P1_R2278_U287 = ~(P1_R2278_U391 & P1_R2278_U229 & P1_R2278_U285); 
assign P1_R2278_U337 = ~(P1_U2785 & P1_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P1_R2278_U355 = ~(P1_U2785 & P1_R2278_U284); 
assign P1_R2278_U369 = ~(P1_R2278_U368 & P1_R2278_U308); 
assign P1_R2278_U373 = ~(P1_R2278_U372 & P1_R2278_U317); 
assign P1_R2278_U374 = ~(P1_R2278_U372 & P1_R2278_U317); 
assign P1_R2278_U382 = ~(P1_R2278_U391 & P1_R2278_U229 & P1_R2278_U285); 
assign P1_R2278_U390 = ~(P1_R2278_U391 & P1_R2278_U229 & P1_R2278_U285); 
assign P1_R2278_U394 = ~(P1_R2278_U148 & P1_R2278_U372); 
assign P1_R2278_U395 = ~(P1_R2278_U383 & P1_R2278_U324); 
assign P1_R2278_U396 = ~(P1_R2278_U150 & P1_R2278_U368); 
assign P1_R2278_U399 = ~(P1_R2278_U154 & P1_R2278_U11 & P1_R2278_U378); 
assign P1_R2278_U402 = ~(P1_R2278_U391 & P1_R2278_U229 & P1_R2278_U285); 
assign P1_R2278_U588 = ~(P1_U2785 & P1_R2278_U62); 
assign P1_R2278_U592 = ~(P1_R2278_U591 & P1_R2278_U590); 
assign P1_R2278_U597 = ~(P1_R2278_U596 & P1_R2278_U595); 
assign P1_R2358_U6 = P1_R2358_U280 & P1_R2358_U278; 
assign P1_R2358_U35 = ~(P1_R2358_U236 & P1_R2358_U220); 
assign P1_R2358_U55 = ~P1_U2635; 
assign P1_R2358_U116 = P1_R2358_U59 & P1_R2358_U258; 
assign P1_R2358_U153 = ~(P1_R2358_U228 & P1_R2358_U230); 
assign P1_R2358_U256 = ~(P1_U2635 & P1_R2358_U474); 
assign P1_R2358_U267 = ~(P1_R2358_U360 & P1_R2358_U357 & P1_R2358_U266 & P1_R2358_U262); 
assign P1_R2358_U281 = ~(P1_U2630 & P1_R2358_U518); 
assign P1_R2358_U318 = ~(P1_R2358_U61 & P1_R2358_U255); 
assign P1_R2358_U351 = ~(P1_R2358_U59 & P1_R2358_U258); 
assign P1_R2358_U359 = ~P1_R2358_U70; 
assign P1_R2358_U361 = ~(P1_R2358_U70 & P1_R2358_U276); 
assign P1_R2358_U362 = ~(P1_R2358_U279 & P1_R2358_U280); 
assign P1_R2358_U452 = ~(P1_R2358_U79 & P1_R2358_U227); 
assign P1_R2358_U454 = ~(P1_R2358_U81 & P1_R2358_U235); 
assign P1_R2358_U504 = ~(P1_U2352 & P1_R2358_U167); 
assign P1_R2358_U513 = ~(P1_U2352 & P1_R2358_U167); 
assign P1_R2099_U20 = ~(P1_R2099_U174 & P1_R2099_U50); 
assign P1_R2099_U310 = ~(P1_R2099_U243 & P1_R2099_U174); 
assign P1_R2337_U50 = ~(P1_R2337_U115 & P1_PHYADDRPOINTER_REG_24__SCAN_IN); 
assign P1_R2337_U154 = ~(P1_R2337_U115 & P1_R2337_U49); 
assign P1_R2096_U50 = ~(P1_R2096_U115 & P1_REIP_REG_24__SCAN_IN); 
assign P1_R2096_U154 = ~(P1_R2096_U115 & P1_R2096_U49); 
assign P1_ADD_405_U50 = ~(P1_ADD_405_U118 & P1_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P1_ADD_405_U134 = ~(P1_ADD_405_U118 & P1_ADD_405_U49); 
assign P1_ADD_515_U50 = ~(P1_ADD_515_U115 & P1_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P1_ADD_515_U130 = ~(P1_ADD_515_U115 & P1_ADD_515_U49); 
assign P3_U2843 = ~(P3_U6111 & P3_U6109 & P3_U6110); 
assign P3_U3849 = P3_U6138 & P3_U3846 & P3_U3848 & P3_U6136 & P3_U3852; 
assign P3_U3854 = P3_U6164 & P3_U6163; 
assign P3_U3856 = P3_U6166 & P3_U6165 & P3_U6167 & P3_U3855; 
assign P3_U3860 = P3_U6176 & P3_U6175 & P3_U6177; 
assign P3_U3861 = P3_U6179 & P3_U6178; 
assign P3_U3865 = P3_U6193 & P3_U6192; 
assign P3_U3868 = P3_U6195 & P3_U6194 & P3_U6196; 
assign P3_U3869 = P3_U6198 & P3_U6197; 
assign P3_U3976 = P3_U6588 & P3_U6585 & P3_U6586 & P3_U6587; 
assign P3_U4108 = P3_U7294 & P3_U7293; 
assign P3_U6113 = ~(P3_SUB_357_1258_U17 & P3_U2393); 
assign P3_U6137 = ~(P3_SUB_357_1258_U85 & P3_U2393); 
assign P3_U6160 = ~(P3_ADD_360_1242_U80 & P3_U2395); 
assign P3_U6203 = ~(P3_ADD_371_1212_U13 & P3_U2360); 
assign P3_U6305 = ~(P3_SUB_357_1258_U19 & P3_U2393); 
assign P3_U6329 = ~(P3_SUB_357_1258_U79 & P3_U2393); 
assign P3_U6568 = ~(P3_U2394 & P3_SUB_357_1258_U17); 
assign P3_U6576 = ~(P3_U2394 & P3_SUB_357_1258_U85); 
assign P3_U6583 = ~(P3_U2396 & P3_ADD_360_1242_U80); 
assign P3_U6595 = ~(P3_U2387 & P3_ADD_371_1212_U13); 
assign P3_U6632 = ~(P3_U2394 & P3_SUB_357_1258_U19); 
assign P3_U6640 = ~(P3_U2394 & P3_SUB_357_1258_U79); 
assign P2_U2802 = P2_U3242 & P2_R2267_U10; 
assign P2_U3112 = ~(P2_U5112 & P2_U5111 & P2_U3793); 
assign P2_U3113 = ~(P2_U5107 & P2_U5106 & P2_U3792); 
assign P2_U3114 = ~(P2_U5102 & P2_U5101 & P2_U3791); 
assign P2_U3115 = ~(P2_U5097 & P2_U5096 & P2_U3790); 
assign P2_U3116 = ~(P2_U5092 & P2_U5091 & P2_U3789); 
assign P2_U3117 = ~(P2_U5087 & P2_U5086 & P2_U3788); 
assign P2_U3118 = ~(P2_U5082 & P2_U5081 & P2_U3787); 
assign P2_U3119 = ~(P2_U5077 & P2_U5076 & P2_U3786); 
assign P2_U3120 = ~(P2_U5055 & P2_U5054 & P2_U3784); 
assign P2_U3121 = ~(P2_U5050 & P2_U5049 & P2_U3783); 
assign P2_U3122 = ~(P2_U5045 & P2_U5044 & P2_U3782); 
assign P2_U3123 = ~(P2_U5040 & P2_U5039 & P2_U3781); 
assign P2_U3124 = ~(P2_U5035 & P2_U5034 & P2_U3780); 
assign P2_U3125 = ~(P2_U5030 & P2_U5029 & P2_U3779); 
assign P2_U3126 = ~(P2_U5025 & P2_U5024 & P2_U3778); 
assign P2_U3127 = ~(P2_U5020 & P2_U5019 & P2_U3777); 
assign P2_U3128 = ~(P2_U4997 & P2_U4996 & P2_U3775); 
assign P2_U3129 = ~(P2_U4992 & P2_U4991 & P2_U3774); 
assign P2_U3130 = ~(P2_U4987 & P2_U4986 & P2_U3773); 
assign P2_U3131 = ~(P2_U4982 & P2_U4981 & P2_U3772); 
assign P2_U3132 = ~(P2_U4977 & P2_U4976 & P2_U3771); 
assign P2_U3133 = ~(P2_U4972 & P2_U4971 & P2_U3770); 
assign P2_U3134 = ~(P2_U4967 & P2_U4966 & P2_U3769); 
assign P2_U3135 = ~(P2_U4962 & P2_U4961 & P2_U3768); 
assign P2_U3136 = ~(P2_U4940 & P2_U4939 & P2_U3766); 
assign P2_U3137 = ~(P2_U4935 & P2_U4934 & P2_U3765); 
assign P2_U3138 = ~(P2_U4930 & P2_U4929 & P2_U3764); 
assign P2_U3139 = ~(P2_U4925 & P2_U4924 & P2_U3763); 
assign P2_U3140 = ~(P2_U4920 & P2_U4919 & P2_U3762); 
assign P2_U3141 = ~(P2_U4915 & P2_U4914 & P2_U3761); 
assign P2_U3142 = ~(P2_U4910 & P2_U4909 & P2_U3760); 
assign P2_U3143 = ~(P2_U4905 & P2_U4904 & P2_U3759); 
assign P2_U3144 = ~(P2_U4882 & P2_U4881 & P2_U3757); 
assign P2_U3145 = ~(P2_U4877 & P2_U4876 & P2_U3756); 
assign P2_U3146 = ~(P2_U4872 & P2_U4871 & P2_U3755); 
assign P2_U3147 = ~(P2_U4867 & P2_U4866 & P2_U3754); 
assign P2_U3148 = ~(P2_U4862 & P2_U4861 & P2_U3753); 
assign P2_U3149 = ~(P2_U4857 & P2_U4856 & P2_U3752); 
assign P2_U3150 = ~(P2_U4852 & P2_U4851 & P2_U3751); 
assign P2_U3151 = ~(P2_U4847 & P2_U4846 & P2_U3750); 
assign P2_U3152 = ~(P2_U4825 & P2_U4824 & P2_U3748); 
assign P2_U3153 = ~(P2_U4820 & P2_U4819 & P2_U3747); 
assign P2_U3154 = ~(P2_U4815 & P2_U4814 & P2_U3746); 
assign P2_U3155 = ~(P2_U4810 & P2_U4809 & P2_U3745); 
assign P2_U3156 = ~(P2_U4805 & P2_U4804 & P2_U3744); 
assign P2_U3157 = ~(P2_U4800 & P2_U4799 & P2_U3743); 
assign P2_U3158 = ~(P2_U4795 & P2_U4794 & P2_U3742); 
assign P2_U3159 = ~(P2_U4790 & P2_U4789 & P2_U3741); 
assign P2_U3160 = ~(P2_U4766 & P2_U4765 & P2_U3739); 
assign P2_U3161 = ~(P2_U4761 & P2_U4760 & P2_U3738); 
assign P2_U3162 = ~(P2_U4756 & P2_U4755 & P2_U3737); 
assign P2_U3163 = ~(P2_U4751 & P2_U4750 & P2_U3736); 
assign P2_U3164 = ~(P2_U4746 & P2_U4745 & P2_U3735); 
assign P2_U3165 = ~(P2_U4741 & P2_U4740 & P2_U3734); 
assign P2_U3166 = ~(P2_U4736 & P2_U4735 & P2_U3733); 
assign P2_U3167 = ~(P2_U4731 & P2_U4730 & P2_U3732); 
assign P2_U3168 = ~(P2_U4708 & P2_U4707 & P2_U3730); 
assign P2_U3169 = ~(P2_U4703 & P2_U4702 & P2_U3729); 
assign P2_U3170 = ~(P2_U4698 & P2_U4697 & P2_U3728); 
assign P2_U3171 = ~(P2_U4693 & P2_U4692 & P2_U3727); 
assign P2_U3172 = ~(P2_U4688 & P2_U4687 & P2_U3726); 
assign P2_U3173 = ~(P2_U4683 & P2_U4682 & P2_U3725); 
assign P2_U3174 = ~(P2_U4678 & P2_U4677 & P2_U3724); 
assign P2_U3175 = ~(P2_U4673 & P2_U4672 & P2_U3723); 
assign P2_U3635 = ~(P2_U8324 & P2_U8323); 
assign P2_U3666 = ~(P2_U8388 & P2_U8387); 
assign P2_U4133 = P2_U6723 & P2_U4446; 
assign P2_U5132 = ~(P2_U2406 & P2_U5128); 
assign P2_U5133 = ~(P2_U5123 & P2_INSTQUEUE_REG_7__7__SCAN_IN); 
assign P2_U5137 = ~(P2_U2405 & P2_U5128); 
assign P2_U5138 = ~(P2_U5123 & P2_INSTQUEUE_REG_7__6__SCAN_IN); 
assign P2_U5142 = ~(P2_U2404 & P2_U5128); 
assign P2_U5143 = ~(P2_U5123 & P2_INSTQUEUE_REG_7__5__SCAN_IN); 
assign P2_U5147 = ~(P2_U2403 & P2_U5128); 
assign P2_U5148 = ~(P2_U5123 & P2_INSTQUEUE_REG_7__4__SCAN_IN); 
assign P2_U5152 = ~(P2_U2402 & P2_U5128); 
assign P2_U5153 = ~(P2_U5123 & P2_INSTQUEUE_REG_7__3__SCAN_IN); 
assign P2_U5157 = ~(P2_U2401 & P2_U5128); 
assign P2_U5158 = ~(P2_U5123 & P2_INSTQUEUE_REG_7__2__SCAN_IN); 
assign P2_U5162 = ~(P2_U2400 & P2_U5128); 
assign P2_U5163 = ~(P2_U5123 & P2_INSTQUEUE_REG_7__1__SCAN_IN); 
assign P2_U5167 = ~(P2_U2399 & P2_U5128); 
assign P2_U5168 = ~(P2_U5123 & P2_INSTQUEUE_REG_7__0__SCAN_IN); 
assign P2_U5189 = ~(P2_U2406 & P2_U5185); 
assign P2_U5190 = ~(P2_U5180 & P2_INSTQUEUE_REG_6__7__SCAN_IN); 
assign P2_U5194 = ~(P2_U2405 & P2_U5185); 
assign P2_U5195 = ~(P2_U5180 & P2_INSTQUEUE_REG_6__6__SCAN_IN); 
assign P2_U5199 = ~(P2_U2404 & P2_U5185); 
assign P2_U5200 = ~(P2_U5180 & P2_INSTQUEUE_REG_6__5__SCAN_IN); 
assign P2_U5204 = ~(P2_U2403 & P2_U5185); 
assign P2_U5205 = ~(P2_U5180 & P2_INSTQUEUE_REG_6__4__SCAN_IN); 
assign P2_U5209 = ~(P2_U2402 & P2_U5185); 
assign P2_U5210 = ~(P2_U5180 & P2_INSTQUEUE_REG_6__3__SCAN_IN); 
assign P2_U5214 = ~(P2_U2401 & P2_U5185); 
assign P2_U5215 = ~(P2_U5180 & P2_INSTQUEUE_REG_6__2__SCAN_IN); 
assign P2_U5219 = ~(P2_U2400 & P2_U5185); 
assign P2_U5220 = ~(P2_U5180 & P2_INSTQUEUE_REG_6__1__SCAN_IN); 
assign P2_U5224 = ~(P2_U2399 & P2_U5185); 
assign P2_U5225 = ~(P2_U5180 & P2_INSTQUEUE_REG_6__0__SCAN_IN); 
assign P2_U5247 = ~(P2_U2406 & P2_U5243); 
assign P2_U5248 = ~(P2_U5238 & P2_INSTQUEUE_REG_5__7__SCAN_IN); 
assign P2_U5252 = ~(P2_U2405 & P2_U5243); 
assign P2_U5253 = ~(P2_U5238 & P2_INSTQUEUE_REG_5__6__SCAN_IN); 
assign P2_U5257 = ~(P2_U2404 & P2_U5243); 
assign P2_U5258 = ~(P2_U5238 & P2_INSTQUEUE_REG_5__5__SCAN_IN); 
assign P2_U5262 = ~(P2_U2403 & P2_U5243); 
assign P2_U5263 = ~(P2_U5238 & P2_INSTQUEUE_REG_5__4__SCAN_IN); 
assign P2_U5267 = ~(P2_U2402 & P2_U5243); 
assign P2_U5268 = ~(P2_U5238 & P2_INSTQUEUE_REG_5__3__SCAN_IN); 
assign P2_U5272 = ~(P2_U2401 & P2_U5243); 
assign P2_U5273 = ~(P2_U5238 & P2_INSTQUEUE_REG_5__2__SCAN_IN); 
assign P2_U5277 = ~(P2_U2400 & P2_U5243); 
assign P2_U5278 = ~(P2_U5238 & P2_INSTQUEUE_REG_5__1__SCAN_IN); 
assign P2_U5282 = ~(P2_U2399 & P2_U5243); 
assign P2_U5283 = ~(P2_U5238 & P2_INSTQUEUE_REG_5__0__SCAN_IN); 
assign P2_U5304 = ~(P2_U2406 & P2_U5300); 
assign P2_U5305 = ~(P2_U5295 & P2_INSTQUEUE_REG_4__7__SCAN_IN); 
assign P2_U5309 = ~(P2_U2405 & P2_U5300); 
assign P2_U5310 = ~(P2_U5295 & P2_INSTQUEUE_REG_4__6__SCAN_IN); 
assign P2_U5314 = ~(P2_U2404 & P2_U5300); 
assign P2_U5315 = ~(P2_U5295 & P2_INSTQUEUE_REG_4__5__SCAN_IN); 
assign P2_U5319 = ~(P2_U2403 & P2_U5300); 
assign P2_U5320 = ~(P2_U5295 & P2_INSTQUEUE_REG_4__4__SCAN_IN); 
assign P2_U5324 = ~(P2_U2402 & P2_U5300); 
assign P2_U5325 = ~(P2_U5295 & P2_INSTQUEUE_REG_4__3__SCAN_IN); 
assign P2_U5329 = ~(P2_U2401 & P2_U5300); 
assign P2_U5330 = ~(P2_U5295 & P2_INSTQUEUE_REG_4__2__SCAN_IN); 
assign P2_U5334 = ~(P2_U2400 & P2_U5300); 
assign P2_U5335 = ~(P2_U5295 & P2_INSTQUEUE_REG_4__1__SCAN_IN); 
assign P2_U5339 = ~(P2_U2399 & P2_U5300); 
assign P2_U5340 = ~(P2_U5295 & P2_INSTQUEUE_REG_4__0__SCAN_IN); 
assign P2_U5362 = ~(P2_U2406 & P2_U5358); 
assign P2_U5363 = ~(P2_U5353 & P2_INSTQUEUE_REG_3__7__SCAN_IN); 
assign P2_U5367 = ~(P2_U2405 & P2_U5358); 
assign P2_U5368 = ~(P2_U5353 & P2_INSTQUEUE_REG_3__6__SCAN_IN); 
assign P2_U5372 = ~(P2_U2404 & P2_U5358); 
assign P2_U5373 = ~(P2_U5353 & P2_INSTQUEUE_REG_3__5__SCAN_IN); 
assign P2_U5377 = ~(P2_U2403 & P2_U5358); 
assign P2_U5378 = ~(P2_U5353 & P2_INSTQUEUE_REG_3__4__SCAN_IN); 
assign P2_U5382 = ~(P2_U2402 & P2_U5358); 
assign P2_U5383 = ~(P2_U5353 & P2_INSTQUEUE_REG_3__3__SCAN_IN); 
assign P2_U5387 = ~(P2_U2401 & P2_U5358); 
assign P2_U5388 = ~(P2_U5353 & P2_INSTQUEUE_REG_3__2__SCAN_IN); 
assign P2_U5392 = ~(P2_U2400 & P2_U5358); 
assign P2_U5393 = ~(P2_U5353 & P2_INSTQUEUE_REG_3__1__SCAN_IN); 
assign P2_U5397 = ~(P2_U2399 & P2_U5358); 
assign P2_U5398 = ~(P2_U5353 & P2_INSTQUEUE_REG_3__0__SCAN_IN); 
assign P2_U5419 = ~(P2_U2406 & P2_U5415); 
assign P2_U5420 = ~(P2_U5410 & P2_INSTQUEUE_REG_2__7__SCAN_IN); 
assign P2_U5424 = ~(P2_U2405 & P2_U5415); 
assign P2_U5425 = ~(P2_U5410 & P2_INSTQUEUE_REG_2__6__SCAN_IN); 
assign P2_U5429 = ~(P2_U2404 & P2_U5415); 
assign P2_U5430 = ~(P2_U5410 & P2_INSTQUEUE_REG_2__5__SCAN_IN); 
assign P2_U5434 = ~(P2_U2403 & P2_U5415); 
assign P2_U5435 = ~(P2_U5410 & P2_INSTQUEUE_REG_2__4__SCAN_IN); 
assign P2_U5439 = ~(P2_U2402 & P2_U5415); 
assign P2_U5440 = ~(P2_U5410 & P2_INSTQUEUE_REG_2__3__SCAN_IN); 
assign P2_U5444 = ~(P2_U2401 & P2_U5415); 
assign P2_U5445 = ~(P2_U5410 & P2_INSTQUEUE_REG_2__2__SCAN_IN); 
assign P2_U5449 = ~(P2_U2400 & P2_U5415); 
assign P2_U5450 = ~(P2_U5410 & P2_INSTQUEUE_REG_2__1__SCAN_IN); 
assign P2_U5454 = ~(P2_U2399 & P2_U5415); 
assign P2_U5455 = ~(P2_U5410 & P2_INSTQUEUE_REG_2__0__SCAN_IN); 
assign P2_U5477 = ~(P2_U2406 & P2_U5473); 
assign P2_U5478 = ~(P2_U5468 & P2_INSTQUEUE_REG_1__7__SCAN_IN); 
assign P2_U5482 = ~(P2_U2405 & P2_U5473); 
assign P2_U5483 = ~(P2_U5468 & P2_INSTQUEUE_REG_1__6__SCAN_IN); 
assign P2_U5487 = ~(P2_U2404 & P2_U5473); 
assign P2_U5488 = ~(P2_U5468 & P2_INSTQUEUE_REG_1__5__SCAN_IN); 
assign P2_U5492 = ~(P2_U2403 & P2_U5473); 
assign P2_U5493 = ~(P2_U5468 & P2_INSTQUEUE_REG_1__4__SCAN_IN); 
assign P2_U5497 = ~(P2_U2402 & P2_U5473); 
assign P2_U5498 = ~(P2_U5468 & P2_INSTQUEUE_REG_1__3__SCAN_IN); 
assign P2_U5502 = ~(P2_U2401 & P2_U5473); 
assign P2_U5503 = ~(P2_U5468 & P2_INSTQUEUE_REG_1__2__SCAN_IN); 
assign P2_U5507 = ~(P2_U2400 & P2_U5473); 
assign P2_U5508 = ~(P2_U5468 & P2_INSTQUEUE_REG_1__1__SCAN_IN); 
assign P2_U5512 = ~(P2_U2399 & P2_U5473); 
assign P2_U5513 = ~(P2_U5468 & P2_INSTQUEUE_REG_1__0__SCAN_IN); 
assign P2_U5534 = ~(P2_U2406 & P2_U5530); 
assign P2_U5535 = ~(P2_U5525 & P2_INSTQUEUE_REG_0__7__SCAN_IN); 
assign P2_U5539 = ~(P2_U2405 & P2_U5530); 
assign P2_U5540 = ~(P2_U5525 & P2_INSTQUEUE_REG_0__6__SCAN_IN); 
assign P2_U5544 = ~(P2_U2404 & P2_U5530); 
assign P2_U5545 = ~(P2_U5525 & P2_INSTQUEUE_REG_0__5__SCAN_IN); 
assign P2_U5549 = ~(P2_U2403 & P2_U5530); 
assign P2_U5550 = ~(P2_U5525 & P2_INSTQUEUE_REG_0__4__SCAN_IN); 
assign P2_U5554 = ~(P2_U2402 & P2_U5530); 
assign P2_U5555 = ~(P2_U5525 & P2_INSTQUEUE_REG_0__3__SCAN_IN); 
assign P2_U5559 = ~(P2_U2401 & P2_U5530); 
assign P2_U5560 = ~(P2_U5525 & P2_INSTQUEUE_REG_0__2__SCAN_IN); 
assign P2_U5564 = ~(P2_U2400 & P2_U5530); 
assign P2_U5565 = ~(P2_U5525 & P2_INSTQUEUE_REG_0__1__SCAN_IN); 
assign P2_U5569 = ~(P2_U2399 & P2_U5530); 
assign P2_U5570 = ~(P2_U5525 & P2_INSTQUEUE_REG_0__0__SCAN_IN); 
assign P2_U6419 = ~(P2_U2380 & P2_R2096_U86); 
assign P2_U6511 = ~(P2_U2379 & P2_R2099_U90); 
assign P2_U6513 = ~(P2_R2182_U92 & P2_U2393); 
assign P2_U6686 = ~(P2_U2392 & P2_R2099_U90); 
assign P2_U6731 = ~(P2_R2267_U10 & P2_U2587); 
assign P2_U6748 = ~(P2_U2588 & P2_R2096_U86); 
assign P2_U8321 = ~(P2_R2256_U20 & P2_U3572); 
assign P1_U2868 = ~(P1_U6278 & P1_U6279 & P1_U6277); 
assign P1_U2900 = ~(P1_U6168 & P1_U6166 & P1_U6167); 
assign P1_U3028 = ~(P1_U3775 & P1_U3776); 
assign P1_U3162 = ~(P1_U4520 & P1_U4519 & P1_U4518 & P1_U4244); 
assign P1_U3466 = ~(P1_U7686 & P1_U7685); 
assign P1_U3835 = P1_U5732 & P1_U5734; 
assign P1_U3837 = P1_U3836 & P1_U5735; 
assign P1_U3932 = P1_U6538 & P1_U6536; 
assign P1_U4017 = P1_U6805 & P1_U6806 & P1_U6807; 
assign P1_U4554 = ~(P1_U4551 & P1_U3587); 
assign P1_U4559 = ~(P1_U4558 & P1_U4557); 
assign P1_U4612 = ~(P1_U4609 & P1_U3596); 
assign P1_U4617 = ~(P1_U4616 & P1_U4615); 
assign P1_U4671 = ~(P1_U4668 & P1_U3605); 
assign P1_U4676 = ~(P1_U4675 & P1_U4674); 
assign P1_U4728 = ~(P1_U4725 & P1_U3614); 
assign P1_U4733 = ~(P1_U4732 & P1_U4731); 
assign P1_U4786 = ~(P1_U4783 & P1_U3623); 
assign P1_U4791 = ~(P1_U4790 & P1_U4789); 
assign P1_U4843 = ~(P1_U4840 & P1_U3632); 
assign P1_U4848 = ~(P1_U4847 & P1_U4846); 
assign P1_U4901 = ~(P1_U4898 & P1_U3641); 
assign P1_U4906 = ~(P1_U4905 & P1_U4904); 
assign P1_U4958 = ~(P1_U4955 & P1_U3650); 
assign P1_U4963 = ~(P1_U4962 & P1_U4961); 
assign P1_U5011 = ~(P1_U5006 & P1_U5010); 
assign P1_U5017 = ~(P1_U5016 & P1_U3361); 
assign P1_U5068 = ~(P1_U5063 & P1_U5067); 
assign P1_U5074 = ~(P1_U5073 & P1_U3365); 
assign P1_U5126 = ~(P1_U5120 & P1_U5125); 
assign P1_U5132 = ~(P1_U5131 & P1_U3368); 
assign P1_U5183 = ~(P1_U5178 & P1_U5182); 
assign P1_U5189 = ~(P1_U5188 & P1_U3372); 
assign P1_U5241 = ~(P1_U5235 & P1_U5240); 
assign P1_U5247 = ~(P1_U5246 & P1_U3375); 
assign P1_U5298 = ~(P1_U5293 & P1_U5297); 
assign P1_U5304 = ~(P1_U5303 & P1_U3379); 
assign P1_U5356 = ~(P1_U5350 & P1_U5355); 
assign P1_U5362 = ~(P1_U5361 & P1_U3382); 
assign P1_U5413 = ~(P1_U5408 & P1_U5412); 
assign P1_U5419 = ~(P1_U5418 & P1_U3386); 
assign P1_U5600 = ~(P1_R2278_U104 & P1_U2377); 
assign P1_U5820 = ~(P1_U2372 & P1_R2278_U104); 
assign P1_U7730 = ~(P1_U5545 & P1_U3404); 
assign P3_ADD_476_U77 = ~(P3_ADD_476_U154 & P3_ADD_476_U153); 
assign P3_ADD_476_U116 = ~P3_ADD_476_U50; 
assign P3_ADD_476_U151 = ~(P3_ADD_476_U50 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_531_U81 = ~(P3_ADD_531_U161 & P3_ADD_531_U160); 
assign P3_ADD_531_U120 = ~P3_ADD_531_U51; 
assign P3_ADD_531_U158 = ~(P3_ADD_531_U51 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_SUB_320_U111 = ~(P3_SUB_320_U99 & P3_SUB_320_U67); 
assign P3_SUB_320_U145 = ~(P3_SUB_320_U99 & P3_SUB_320_U67); 
assign P3_ADD_318_U77 = ~(P3_ADD_318_U154 & P3_ADD_318_U153); 
assign P3_ADD_318_U116 = ~P3_ADD_318_U50; 
assign P3_ADD_318_U151 = ~(P3_ADD_318_U50 & P3_PHYADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_315_U73 = ~(P3_ADD_315_U146 & P3_ADD_315_U145); 
assign P3_ADD_315_U113 = ~P3_ADD_315_U50; 
assign P3_ADD_315_U143 = ~(P3_ADD_315_U50 & P3_PHYADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_360_1242_U12 = P3_ADD_360_1242_U173 & P3_ADD_360_1242_U63; 
assign P3_ADD_360_1242_U66 = ~(P3_ADD_360_1242_U103 & P3_ADD_360_1242_U161); 
assign P3_ADD_360_1242_U170 = ~(P3_ADD_360_1242_U161 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_360_1242_U241 = ~(P3_ADD_360_1242_U161 & P3_ADD_360_1242_U65); 
assign P3_ADD_467_U77 = ~(P3_ADD_467_U154 & P3_ADD_467_U153); 
assign P3_ADD_467_U116 = ~P3_ADD_467_U50; 
assign P3_ADD_467_U151 = ~(P3_ADD_467_U50 & P3_REIP_REG_25__SCAN_IN); 
assign P3_ADD_430_U77 = ~(P3_ADD_430_U154 & P3_ADD_430_U153); 
assign P3_ADD_430_U116 = ~P3_ADD_430_U50; 
assign P3_ADD_430_U151 = ~(P3_ADD_430_U50 & P3_REIP_REG_25__SCAN_IN); 
assign P3_ADD_380_U81 = ~(P3_ADD_380_U161 & P3_ADD_380_U160); 
assign P3_ADD_380_U120 = ~P3_ADD_380_U51; 
assign P3_ADD_380_U158 = ~(P3_ADD_380_U51 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_344_U81 = ~(P3_ADD_344_U161 & P3_ADD_344_U160); 
assign P3_ADD_344_U120 = ~P3_ADD_344_U51; 
assign P3_ADD_344_U158 = ~(P3_ADD_344_U51 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_339_U77 = ~(P3_ADD_339_U154 & P3_ADD_339_U153); 
assign P3_ADD_339_U116 = ~P3_ADD_339_U50; 
assign P3_ADD_339_U151 = ~(P3_ADD_339_U50 & P3_PHYADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_541_U77 = ~(P3_ADD_541_U154 & P3_ADD_541_U153); 
assign P3_ADD_541_U116 = ~P3_ADD_541_U50; 
assign P3_ADD_541_U151 = ~(P3_ADD_541_U50 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_SUB_357_1258_U294 = ~(P3_SUB_357_1258_U223 & P3_SUB_357_1258_U60); 
assign P3_SUB_357_1258_U296 = ~(P3_SUB_357_1258_U352 & P3_SUB_357_1258_U351 & P3_SUB_357_1258_U295); 
assign P3_SUB_357_1258_U354 = ~(P3_SUB_357_1258_U297 & P3_SUB_357_1258_U39); 
assign P3_SUB_357_1258_U361 = ~(P3_SUB_357_1258_U359 & P3_SUB_357_1258_U223); 
assign P3_ADD_515_U77 = ~(P3_ADD_515_U154 & P3_ADD_515_U153); 
assign P3_ADD_515_U116 = ~P3_ADD_515_U50; 
assign P3_ADD_515_U151 = ~(P3_ADD_515_U50 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_394_U76 = ~(P3_ADD_394_U156 & P3_ADD_394_U155); 
assign P3_ADD_394_U119 = ~P3_ADD_394_U50; 
assign P3_ADD_394_U153 = ~(P3_ADD_394_U50 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_441_U77 = ~(P3_ADD_441_U154 & P3_ADD_441_U153); 
assign P3_ADD_441_U116 = ~P3_ADD_441_U50; 
assign P3_ADD_441_U151 = ~(P3_ADD_441_U50 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_349_U81 = ~(P3_ADD_349_U161 & P3_ADD_349_U160); 
assign P3_ADD_349_U120 = ~P3_ADD_349_U51; 
assign P3_ADD_349_U158 = ~(P3_ADD_349_U51 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_405_U76 = ~(P3_ADD_405_U156 & P3_ADD_405_U155); 
assign P3_ADD_405_U119 = ~P3_ADD_405_U50; 
assign P3_ADD_405_U153 = ~(P3_ADD_405_U50 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_553_U81 = ~(P3_ADD_553_U161 & P3_ADD_553_U160); 
assign P3_ADD_553_U120 = ~P3_ADD_553_U51; 
assign P3_ADD_553_U158 = ~(P3_ADD_553_U51 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_558_U81 = ~(P3_ADD_558_U161 & P3_ADD_558_U160); 
assign P3_ADD_558_U120 = ~P3_ADD_558_U51; 
assign P3_ADD_558_U158 = ~(P3_ADD_558_U51 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_385_U81 = ~(P3_ADD_385_U161 & P3_ADD_385_U160); 
assign P3_ADD_385_U120 = ~P3_ADD_385_U51; 
assign P3_ADD_385_U158 = ~(P3_ADD_385_U51 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_547_U81 = ~(P3_ADD_547_U161 & P3_ADD_547_U160); 
assign P3_ADD_547_U120 = ~P3_ADD_547_U51; 
assign P3_ADD_547_U158 = ~(P3_ADD_547_U51 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_371_1212_U81 = ~(P3_ADD_371_1212_U248 & P3_ADD_371_1212_U247); 
assign P3_ADD_371_1212_U171 = ~P3_ADD_371_1212_U68; 
assign P3_ADD_371_1212_U179 = ~(P3_ADD_371_1212_U69 & P3_ADD_371_1212_U68); 
assign P3_ADD_371_1212_U181 = ~(P3_ADD_371_1212_U66 & P3_ADD_371_1212_U180); 
assign P3_ADD_494_U77 = ~(P3_ADD_494_U154 & P3_ADD_494_U153); 
assign P3_ADD_494_U116 = ~P3_ADD_494_U50; 
assign P3_ADD_494_U151 = ~(P3_ADD_494_U50 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_536_U77 = ~(P3_ADD_536_U154 & P3_ADD_536_U153); 
assign P3_ADD_536_U116 = ~P3_ADD_536_U50; 
assign P3_ADD_536_U151 = ~(P3_ADD_536_U50 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P2_R2099_U35 = ~(P2_U2733 & P2_R2099_U129); 
assign P2_R2099_U215 = ~(P2_R2099_U129 & P2_R2099_U34); 
assign P2_ADD_391_1196_U10 = P2_ADD_391_1196_U201 & P2_ADD_391_1196_U199; 
assign P2_ADD_391_1196_U35 = ~(P2_ADD_391_1196_U190 & P2_ADD_391_1196_U189); 
assign P2_ADD_391_1196_U42 = ~P2_R2182_U92; 
assign P2_ADD_391_1196_U65 = ~P2_R2096_U86; 
assign P2_ADD_391_1196_U155 = P2_ADD_391_1196_U464 & P2_ADD_391_1196_U463; 
assign P2_ADD_391_1196_U159 = ~(P2_R2096_U93 & P2_R2182_U92); 
assign P2_ADD_391_1196_U224 = P2_R2096_U93 | P2_R2182_U92; 
assign P2_ADD_391_1196_U288 = P2_R2182_U92 | P2_R2096_U93; 
assign P2_ADD_391_1196_U293 = P2_R2096_U93 | P2_R2182_U92; 
assign P2_ADD_391_1196_U315 = ~(P2_ADD_391_1196_U187 & P2_ADD_391_1196_U313); 
assign P2_ADD_391_1196_U457 = ~(P2_R2182_U92 & P2_ADD_391_1196_U43); 
assign P2_ADD_391_1196_U461 = ~(P2_R2096_U94 & P2_ADD_391_1196_U44); 
assign P2_ADD_391_1196_U467 = ~(P2_ADD_391_1196_U466 & P2_ADD_391_1196_U465); 
assign P2_R2182_U18 = P2_U2695 & P2_R2182_U17; 
assign P2_R2182_U91 = ~(P2_R2182_U293 & P2_R2182_U292); 
assign P2_R2182_U148 = ~P2_R2182_U17; 
assign P2_R2182_U288 = ~(P2_R2182_U28 & P2_R2182_U17); 
assign P2_R2182_U291 = ~(P2_R2182_U147 & P2_U2696); 
assign P2_R2027_U81 = ~(P2_R2027_U161 & P2_R2027_U160); 
assign P2_R2027_U120 = ~P2_R2027_U51; 
assign P2_R2027_U158 = ~(P2_R2027_U51 & P2_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P2_R2337_U75 = ~(P2_R2337_U152 & P2_R2337_U151); 
assign P2_R2337_U117 = ~P2_R2337_U51; 
assign P2_R2337_U149 = ~(P2_R2337_U51 & P2_PHYADDRPOINTER_REG_26__SCAN_IN); 
assign P2_R2096_U11 = P2_U2625 & P2_R2096_U10; 
assign P2_R2096_U85 = ~(P2_R2096_U234 & P2_R2096_U233); 
assign P2_R2096_U159 = ~P2_R2096_U10; 
assign P2_R2096_U229 = ~(P2_R2096_U44 & P2_R2096_U10); 
assign P2_R2096_U232 = ~(P2_R2096_U158 & P2_U2626); 
assign P2_R2256_U14 = ~(P2_U3624 & P2_R2256_U42); 
assign P2_R2256_U52 = ~(P2_R2256_U42 & P2_R2256_U13); 
assign P2_R1957_U111 = ~(P2_R1957_U99 & P2_R1957_U67); 
assign P2_R1957_U145 = ~(P2_R1957_U99 & P2_R1957_U67); 
assign P2_R2278_U64 = ~P2_U2803; 
assign P2_R2278_U127 = P2_R2278_U259 & P2_R2278_U263; 
assign P2_R2278_U191 = P2_R2278_U513 & P2_R2278_U512; 
assign P2_R2278_U209 = ~P2_R2278_U165; 
assign P2_R2278_U211 = ~(P2_R2278_U210 & P2_R2278_U165); 
assign P2_R2278_U212 = ~P2_R2278_U20; 
assign P2_R2278_U266 = P2_U2803 | P2_INSTADDRPOINTER_REG_18__SCAN_IN; 
assign P2_R2278_U268 = ~(P2_U2803 & P2_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P2_R2278_U328 = ~(P2_R2278_U261 & P2_R2278_U263); 
assign P2_R2278_U345 = ~(P2_R2278_U207 & P2_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P2_R2278_U409 = ~(P2_R2278_U18 & P2_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P2_R2278_U411 = ~(P2_R2278_U18 & P2_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P2_R2278_U499 = ~(P2_U2803 & P2_R2278_U65); 
assign P2_R2278_U501 = ~(P2_U2803 & P2_R2278_U65); 
assign P2_R2278_U505 = ~(P2_R2278_U41 & P2_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P2_R2278_U507 = ~(P2_R2278_U41 & P2_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P2_R2278_U516 = ~(P2_R2278_U515 & P2_R2278_U514); 
assign P2_ADD_394_U66 = ~(P2_ADD_394_U134 & P2_ADD_394_U133); 
assign P2_ADD_394_U119 = ~P2_ADD_394_U50; 
assign P2_ADD_394_U183 = ~(P2_ADD_394_U50 & P2_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P2_R2267_U75 = P2_R2267_U154 & P2_R2267_U153; 
assign P2_R2267_U107 = ~P2_R2267_U36; 
assign P2_R2267_U123 = ~(P2_U2776 & P2_R2267_U122); 
assign P2_R2267_U151 = ~(P2_U2775 & P2_R2267_U36); 
assign P2_ADD_371_1212_U35 = ~P2_R2256_U20; 
assign P2_ADD_371_1212_U140 = ~P2_ADD_371_1212_U116; 
assign P2_ADD_371_1212_U142 = ~(P2_ADD_371_1212_U141 & P2_ADD_371_1212_U116); 
assign P2_ADD_371_1212_U149 = P2_R2256_U20 | P2_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P2_ADD_371_1212_U151 = ~(P2_R2256_U20 & P2_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P2_ADD_371_1212_U225 = ~(P2_ADD_371_1212_U115 & P2_ADD_371_1212_U116); 
assign P2_ADD_371_1212_U234 = ~(P2_R2256_U20 & P2_ADD_371_1212_U36); 
assign P2_ADD_371_1212_U236 = ~(P2_R2256_U20 & P2_ADD_371_1212_U36); 
assign P2_ADD_371_1212_U258 = ~(P2_ADD_371_1212_U33 & P2_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P2_ADD_371_1212_U260 = ~(P2_ADD_371_1212_U33 & P2_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P1_R2278_U40 = ~(P1_R2278_U43 & P1_R2278_U250); 
assign P1_R2278_U87 = ~(P1_R2278_U392 & P1_R2278_U92 & P1_R2278_U93); 
assign P1_R2278_U145 = P1_R2278_U95 & P1_R2278_U94; 
assign P1_R2278_U156 = P1_R2278_U14 & P1_R2278_U400 & P1_R2278_U399; 
assign P1_R2278_U162 = P1_R2278_U369 & P1_R2278_U76; 
assign P1_R2278_U227 = ~(P1_R2278_U356 & P1_R2278_U355); 
assign P1_R2278_U249 = ~P1_R2278_U43; 
assign P1_R2278_U270 = ~(P1_R2278_U180 & P1_R2278_U247); 
assign P1_R2278_U357 = ~(P1_R2278_U356 & P1_R2278_U63); 
assign P1_R2278_U380 = ~P1_R2278_U94; 
assign P1_R2278_U384 = ~P1_R2278_U95; 
assign P1_R2278_U386 = ~P1_R2278_U93; 
assign P1_R2278_U387 = ~P1_R2278_U96; 
assign P1_R2278_U408 = ~(P1_R2278_U374 & P1_R2278_U85); 
assign P1_R2278_U589 = ~(P1_R2278_U63 & P1_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P1_R2358_U36 = ~(P1_R2358_U35 & P1_R2358_U218); 
assign P1_R2358_U80 = ~(P1_R2358_U452 & P1_R2358_U451); 
assign P1_R2358_U82 = ~(P1_R2358_U454 & P1_R2358_U453); 
assign P1_R2358_U104 = P1_R2358_U281 & P1_R2358_U280; 
assign P1_R2358_U129 = P1_R2358_U361 & P1_R2358_U277; 
assign P1_R2358_U138 = P1_R2358_U362 & P1_R2358_U281; 
assign P1_R2358_U166 = ~P1_U2660; 
assign P1_R2358_U199 = ~(P1_R2358_U268 & P1_R2358_U264 & P1_R2358_U267); 
assign P1_R2358_U231 = ~P1_R2358_U153; 
assign P1_R2358_U237 = ~P1_R2358_U35; 
assign P1_R2358_U257 = ~(P1_R2358_U11 & P1_R2358_U55); 
assign P1_R2358_U282 = ~(P1_R2358_U505 & P1_R2358_U504 & P1_R2358_U44); 
assign P1_R2358_U321 = ~(P1_R2358_U54 & P1_R2358_U153); 
assign P1_R2358_U345 = ~(P1_R2358_U281 & P1_R2358_U280); 
assign P1_R2358_U356 = ~(P1_R2358_U11 & P1_R2358_U55); 
assign P1_R2358_U363 = ~(P1_R2358_U362 & P1_R2358_U281); 
assign P1_R2358_U449 = ~(P1_R2358_U332 & P1_R2358_U153); 
assign P1_R2358_U503 = ~(P1_U2660 & P1_R2358_U23); 
assign P1_R2358_U511 = ~(P1_U2660 & P1_R2358_U23); 
assign P1_R2358_U515 = ~(P1_R2358_U514 & P1_R2358_U513); 
assign P1_R2099_U72 = ~(P1_R2099_U311 & P1_R2099_U310); 
assign P1_R2099_U175 = ~P1_R2099_U20; 
assign P1_R2099_U309 = ~(P1_R2099_U49 & P1_R2099_U20); 
assign P1_R2337_U77 = ~(P1_R2337_U154 & P1_R2337_U153); 
assign P1_R2337_U116 = ~P1_R2337_U50; 
assign P1_R2337_U151 = ~(P1_R2337_U50 & P1_PHYADDRPOINTER_REG_25__SCAN_IN); 
assign P1_R2096_U77 = ~(P1_R2096_U154 & P1_R2096_U153); 
assign P1_R2096_U116 = ~P1_R2096_U50; 
assign P1_R2096_U151 = ~(P1_R2096_U50 & P1_REIP_REG_25__SCAN_IN); 
assign P1_ADD_405_U66 = ~(P1_ADD_405_U134 & P1_ADD_405_U133); 
assign P1_ADD_405_U119 = ~P1_ADD_405_U50; 
assign P1_ADD_405_U183 = ~(P1_ADD_405_U50 & P1_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P1_ADD_515_U65 = ~(P1_ADD_515_U130 & P1_ADD_515_U129); 
assign P1_ADD_515_U116 = ~P1_ADD_515_U50; 
assign P1_ADD_515_U179 = ~(P1_ADD_515_U50 & P1_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_U2808 = ~(P3_U6582 & P3_U6581 & P3_U6584 & P3_U6583 & P3_U3976); 
assign P3_U2809 = ~(P3_U6574 & P3_U6573 & P3_U6575 & P3_U3975 & P3_U6576); 
assign P3_U2810 = ~(P3_U6566 & P3_U6565 & P3_U6567 & P3_U3974 & P3_U6568); 
assign P3_U3857 = P3_U6161 & P3_U6162 & P3_U3854 & P3_U3856 & P3_U6160; 
assign P3_U3862 = P3_U3859 & P3_U3858 & P3_U3860 & P3_U3861; 
assign P3_U3977 = P3_U6596 & P3_U6593 & P3_U6594 & P3_U6595; 
assign P3_U6132 = ~(P3_U6113 & P3_U3841); 
assign P3_U6156 = ~(P3_U6137 & P3_U3849); 
assign P3_U6184 = ~(P3_ADD_360_1242_U12 & P3_U2395); 
assign P3_U6186 = ~(P3_ADD_558_U81 & P3_U3220); 
assign P3_U6187 = ~(P3_ADD_553_U81 & P3_U4298); 
assign P3_U6188 = ~(P3_ADD_547_U81 & P3_U4299); 
assign P3_U6191 = ~(P3_ADD_531_U81 & P3_U2354); 
assign P3_U6199 = ~(P3_ADD_385_U81 & P3_U2358); 
assign P3_U6200 = ~(P3_ADD_380_U81 & P3_U2359); 
assign P3_U6201 = ~(P3_ADD_349_U81 & P3_U4306); 
assign P3_U6202 = ~(P3_ADD_344_U81 & P3_U2362); 
assign P3_U6213 = ~(P3_ADD_541_U77 & P3_U4300); 
assign P3_U6214 = ~(P3_ADD_536_U77 & P3_U4301); 
assign P3_U6217 = ~(P3_ADD_515_U77 & P3_U4302); 
assign P3_U6218 = ~(P3_ADD_494_U77 & P3_U2356); 
assign P3_U6219 = ~(P3_ADD_476_U77 & P3_U4303); 
assign P3_U6220 = ~(P3_ADD_441_U77 & P3_U4304); 
assign P3_U6221 = ~(P3_ADD_405_U76 & P3_U4305); 
assign P3_U6222 = ~(P3_ADD_394_U76 & P3_U2357); 
assign P3_U6227 = ~(P3_ADD_371_1212_U81 & P3_U2360); 
assign P3_U6591 = ~(P3_U2396 & P3_ADD_360_1242_U12); 
assign P3_U6597 = ~(P3_ADD_318_U77 & P3_U2398); 
assign P3_U6602 = ~(P3_ADD_339_U77 & P3_U2388); 
assign P3_U6603 = ~(P3_U2387 & P3_ADD_371_1212_U81); 
assign P3_U6606 = ~(P3_ADD_315_U73 & P3_U2397); 
assign P3_U7302 = ~(P3_ADD_467_U77 & P3_U2601); 
assign P3_U7304 = ~(P3_ADD_430_U77 & P3_U2405); 
assign P2_U2801 = P2_U3242 & P2_R2267_U75; 
assign P2_U2874 = ~(P2_U6511 & P2_U6512 & P2_U6510); 
assign P2_U3048 = ~(P2_U5570 & P2_U5569 & P2_U3865); 
assign P2_U3049 = ~(P2_U5565 & P2_U5564 & P2_U3864); 
assign P2_U3050 = ~(P2_U5560 & P2_U5559 & P2_U3863); 
assign P2_U3051 = ~(P2_U5555 & P2_U5554 & P2_U3862); 
assign P2_U3052 = ~(P2_U5550 & P2_U5549 & P2_U3861); 
assign P2_U3053 = ~(P2_U5545 & P2_U5544 & P2_U3860); 
assign P2_U3054 = ~(P2_U5540 & P2_U5539 & P2_U3859); 
assign P2_U3055 = ~(P2_U5535 & P2_U5534 & P2_U3858); 
assign P2_U3056 = ~(P2_U5513 & P2_U5512 & P2_U3856); 
assign P2_U3057 = ~(P2_U5508 & P2_U5507 & P2_U3855); 
assign P2_U3058 = ~(P2_U5503 & P2_U5502 & P2_U3854); 
assign P2_U3059 = ~(P2_U5498 & P2_U5497 & P2_U3853); 
assign P2_U3060 = ~(P2_U5493 & P2_U5492 & P2_U3852); 
assign P2_U3061 = ~(P2_U5488 & P2_U5487 & P2_U3851); 
assign P2_U3062 = ~(P2_U5483 & P2_U5482 & P2_U3850); 
assign P2_U3063 = ~(P2_U5478 & P2_U5477 & P2_U3849); 
assign P2_U3064 = ~(P2_U5455 & P2_U5454 & P2_U3847); 
assign P2_U3065 = ~(P2_U5450 & P2_U5449 & P2_U3846); 
assign P2_U3066 = ~(P2_U5445 & P2_U5444 & P2_U3845); 
assign P2_U3067 = ~(P2_U5440 & P2_U5439 & P2_U3844); 
assign P2_U3068 = ~(P2_U5435 & P2_U5434 & P2_U3843); 
assign P2_U3069 = ~(P2_U5430 & P2_U5429 & P2_U3842); 
assign P2_U3070 = ~(P2_U5425 & P2_U5424 & P2_U3841); 
assign P2_U3071 = ~(P2_U5420 & P2_U5419 & P2_U3840); 
assign P2_U3072 = ~(P2_U5398 & P2_U5397 & P2_U3838); 
assign P2_U3073 = ~(P2_U5393 & P2_U5392 & P2_U3837); 
assign P2_U3074 = ~(P2_U5388 & P2_U5387 & P2_U3836); 
assign P2_U3075 = ~(P2_U5383 & P2_U5382 & P2_U3835); 
assign P2_U3076 = ~(P2_U5378 & P2_U5377 & P2_U3834); 
assign P2_U3077 = ~(P2_U5373 & P2_U5372 & P2_U3833); 
assign P2_U3078 = ~(P2_U5368 & P2_U5367 & P2_U3832); 
assign P2_U3079 = ~(P2_U5363 & P2_U5362 & P2_U3831); 
assign P2_U3080 = ~(P2_U5340 & P2_U5339 & P2_U3829); 
assign P2_U3081 = ~(P2_U5335 & P2_U5334 & P2_U3828); 
assign P2_U3082 = ~(P2_U5330 & P2_U5329 & P2_U3827); 
assign P2_U3083 = ~(P2_U5325 & P2_U5324 & P2_U3826); 
assign P2_U3084 = ~(P2_U5320 & P2_U5319 & P2_U3825); 
assign P2_U3085 = ~(P2_U5315 & P2_U5314 & P2_U3824); 
assign P2_U3086 = ~(P2_U5310 & P2_U5309 & P2_U3823); 
assign P2_U3087 = ~(P2_U5305 & P2_U5304 & P2_U3822); 
assign P2_U3088 = ~(P2_U5283 & P2_U5282 & P2_U3820); 
assign P2_U3089 = ~(P2_U5278 & P2_U5277 & P2_U3819); 
assign P2_U3090 = ~(P2_U5273 & P2_U5272 & P2_U3818); 
assign P2_U3091 = ~(P2_U5268 & P2_U5267 & P2_U3817); 
assign P2_U3092 = ~(P2_U5263 & P2_U5262 & P2_U3816); 
assign P2_U3093 = ~(P2_U5258 & P2_U5257 & P2_U3815); 
assign P2_U3094 = ~(P2_U5253 & P2_U5252 & P2_U3814); 
assign P2_U3095 = ~(P2_U5248 & P2_U5247 & P2_U3813); 
assign P2_U3096 = ~(P2_U5225 & P2_U5224 & P2_U3811); 
assign P2_U3097 = ~(P2_U5220 & P2_U5219 & P2_U3810); 
assign P2_U3098 = ~(P2_U5215 & P2_U5214 & P2_U3809); 
assign P2_U3099 = ~(P2_U5210 & P2_U5209 & P2_U3808); 
assign P2_U3100 = ~(P2_U5205 & P2_U5204 & P2_U3807); 
assign P2_U3101 = ~(P2_U5200 & P2_U5199 & P2_U3806); 
assign P2_U3102 = ~(P2_U5195 & P2_U5194 & P2_U3805); 
assign P2_U3103 = ~(P2_U5190 & P2_U5189 & P2_U3804); 
assign P2_U3104 = ~(P2_U5168 & P2_U5167 & P2_U3802); 
assign P2_U3105 = ~(P2_U5163 & P2_U5162 & P2_U3801); 
assign P2_U3106 = ~(P2_U5158 & P2_U5157 & P2_U3800); 
assign P2_U3107 = ~(P2_U5153 & P2_U5152 & P2_U3799); 
assign P2_U3108 = ~(P2_U5148 & P2_U5147 & P2_U3798); 
assign P2_U3109 = ~(P2_U5143 & P2_U5142 & P2_U3797); 
assign P2_U3110 = ~(P2_U5138 & P2_U5137 & P2_U3796); 
assign P2_U3111 = ~(P2_U5133 & P2_U5132 & P2_U3795); 
assign P2_U3634 = ~(P2_U8322 & P2_U8321); 
assign P2_U4115 = P2_U6683 & P2_U4446 & P2_U6686; 
assign P2_U4137 = P2_U6731 & P2_U4446; 
assign P2_U6356 = ~(P2_ADD_391_1196_U10 & P2_U2397); 
assign P2_U6424 = ~(P2_U2380 & P2_R2096_U85); 
assign P2_U6516 = ~(P2_R2182_U91 & P2_U2393); 
assign P2_U6739 = ~(P2_R2267_U75 & P2_U2587); 
assign P2_U6756 = ~(P2_U2588 & P2_R2096_U85); 
assign P2_U8385 = ~(P2_R2337_U75 & P2_U3284); 
assign P1_U2659 = ~(P1_U6804 & P1_U4017); 
assign P1_U2995 = ~(P1_U5821 & P1_U5819 & P1_U5820 & P1_U5823 & P1_U5822); 
assign P1_U3027 = ~(P1_U3778 & P1_U3780 & P1_U5600); 
assign P1_U3475 = ~(P1_U7730 & P1_U7729); 
assign P1_U4563 = ~(P1_U2397 & P1_U4559); 
assign P1_U4564 = ~(P1_U4554 & P1_INSTQUEUE_REG_15__7__SCAN_IN); 
assign P1_U4568 = ~(P1_U2396 & P1_U4559); 
assign P1_U4569 = ~(P1_U4554 & P1_INSTQUEUE_REG_15__6__SCAN_IN); 
assign P1_U4573 = ~(P1_U2395 & P1_U4559); 
assign P1_U4574 = ~(P1_U4554 & P1_INSTQUEUE_REG_15__5__SCAN_IN); 
assign P1_U4578 = ~(P1_U2394 & P1_U4559); 
assign P1_U4579 = ~(P1_U4554 & P1_INSTQUEUE_REG_15__4__SCAN_IN); 
assign P1_U4583 = ~(P1_U2393 & P1_U4559); 
assign P1_U4584 = ~(P1_U4554 & P1_INSTQUEUE_REG_15__3__SCAN_IN); 
assign P1_U4588 = ~(P1_U2392 & P1_U4559); 
assign P1_U4589 = ~(P1_U4554 & P1_INSTQUEUE_REG_15__2__SCAN_IN); 
assign P1_U4593 = ~(P1_U2391 & P1_U4559); 
assign P1_U4594 = ~(P1_U4554 & P1_INSTQUEUE_REG_15__1__SCAN_IN); 
assign P1_U4598 = ~(P1_U2390 & P1_U4559); 
assign P1_U4599 = ~(P1_U4554 & P1_INSTQUEUE_REG_15__0__SCAN_IN); 
assign P1_U4621 = ~(P1_U2397 & P1_U4617); 
assign P1_U4622 = ~(P1_U4612 & P1_INSTQUEUE_REG_14__7__SCAN_IN); 
assign P1_U4626 = ~(P1_U2396 & P1_U4617); 
assign P1_U4627 = ~(P1_U4612 & P1_INSTQUEUE_REG_14__6__SCAN_IN); 
assign P1_U4631 = ~(P1_U2395 & P1_U4617); 
assign P1_U4632 = ~(P1_U4612 & P1_INSTQUEUE_REG_14__5__SCAN_IN); 
assign P1_U4636 = ~(P1_U2394 & P1_U4617); 
assign P1_U4637 = ~(P1_U4612 & P1_INSTQUEUE_REG_14__4__SCAN_IN); 
assign P1_U4641 = ~(P1_U2393 & P1_U4617); 
assign P1_U4642 = ~(P1_U4612 & P1_INSTQUEUE_REG_14__3__SCAN_IN); 
assign P1_U4646 = ~(P1_U2392 & P1_U4617); 
assign P1_U4647 = ~(P1_U4612 & P1_INSTQUEUE_REG_14__2__SCAN_IN); 
assign P1_U4651 = ~(P1_U2391 & P1_U4617); 
assign P1_U4652 = ~(P1_U4612 & P1_INSTQUEUE_REG_14__1__SCAN_IN); 
assign P1_U4656 = ~(P1_U2390 & P1_U4617); 
assign P1_U4657 = ~(P1_U4612 & P1_INSTQUEUE_REG_14__0__SCAN_IN); 
assign P1_U4680 = ~(P1_U2397 & P1_U4676); 
assign P1_U4681 = ~(P1_U4671 & P1_INSTQUEUE_REG_13__7__SCAN_IN); 
assign P1_U4685 = ~(P1_U2396 & P1_U4676); 
assign P1_U4686 = ~(P1_U4671 & P1_INSTQUEUE_REG_13__6__SCAN_IN); 
assign P1_U4690 = ~(P1_U2395 & P1_U4676); 
assign P1_U4691 = ~(P1_U4671 & P1_INSTQUEUE_REG_13__5__SCAN_IN); 
assign P1_U4695 = ~(P1_U2394 & P1_U4676); 
assign P1_U4696 = ~(P1_U4671 & P1_INSTQUEUE_REG_13__4__SCAN_IN); 
assign P1_U4700 = ~(P1_U2393 & P1_U4676); 
assign P1_U4701 = ~(P1_U4671 & P1_INSTQUEUE_REG_13__3__SCAN_IN); 
assign P1_U4705 = ~(P1_U2392 & P1_U4676); 
assign P1_U4706 = ~(P1_U4671 & P1_INSTQUEUE_REG_13__2__SCAN_IN); 
assign P1_U4710 = ~(P1_U2391 & P1_U4676); 
assign P1_U4711 = ~(P1_U4671 & P1_INSTQUEUE_REG_13__1__SCAN_IN); 
assign P1_U4715 = ~(P1_U2390 & P1_U4676); 
assign P1_U4716 = ~(P1_U4671 & P1_INSTQUEUE_REG_13__0__SCAN_IN); 
assign P1_U4737 = ~(P1_U2397 & P1_U4733); 
assign P1_U4738 = ~(P1_U4728 & P1_INSTQUEUE_REG_12__7__SCAN_IN); 
assign P1_U4742 = ~(P1_U2396 & P1_U4733); 
assign P1_U4743 = ~(P1_U4728 & P1_INSTQUEUE_REG_12__6__SCAN_IN); 
assign P1_U4747 = ~(P1_U2395 & P1_U4733); 
assign P1_U4748 = ~(P1_U4728 & P1_INSTQUEUE_REG_12__5__SCAN_IN); 
assign P1_U4752 = ~(P1_U2394 & P1_U4733); 
assign P1_U4753 = ~(P1_U4728 & P1_INSTQUEUE_REG_12__4__SCAN_IN); 
assign P1_U4757 = ~(P1_U2393 & P1_U4733); 
assign P1_U4758 = ~(P1_U4728 & P1_INSTQUEUE_REG_12__3__SCAN_IN); 
assign P1_U4762 = ~(P1_U2392 & P1_U4733); 
assign P1_U4763 = ~(P1_U4728 & P1_INSTQUEUE_REG_12__2__SCAN_IN); 
assign P1_U4767 = ~(P1_U2391 & P1_U4733); 
assign P1_U4768 = ~(P1_U4728 & P1_INSTQUEUE_REG_12__1__SCAN_IN); 
assign P1_U4772 = ~(P1_U2390 & P1_U4733); 
assign P1_U4773 = ~(P1_U4728 & P1_INSTQUEUE_REG_12__0__SCAN_IN); 
assign P1_U4795 = ~(P1_U2397 & P1_U4791); 
assign P1_U4796 = ~(P1_U4786 & P1_INSTQUEUE_REG_11__7__SCAN_IN); 
assign P1_U4800 = ~(P1_U2396 & P1_U4791); 
assign P1_U4801 = ~(P1_U4786 & P1_INSTQUEUE_REG_11__6__SCAN_IN); 
assign P1_U4805 = ~(P1_U2395 & P1_U4791); 
assign P1_U4806 = ~(P1_U4786 & P1_INSTQUEUE_REG_11__5__SCAN_IN); 
assign P1_U4810 = ~(P1_U2394 & P1_U4791); 
assign P1_U4811 = ~(P1_U4786 & P1_INSTQUEUE_REG_11__4__SCAN_IN); 
assign P1_U4815 = ~(P1_U2393 & P1_U4791); 
assign P1_U4816 = ~(P1_U4786 & P1_INSTQUEUE_REG_11__3__SCAN_IN); 
assign P1_U4820 = ~(P1_U2392 & P1_U4791); 
assign P1_U4821 = ~(P1_U4786 & P1_INSTQUEUE_REG_11__2__SCAN_IN); 
assign P1_U4825 = ~(P1_U2391 & P1_U4791); 
assign P1_U4826 = ~(P1_U4786 & P1_INSTQUEUE_REG_11__1__SCAN_IN); 
assign P1_U4830 = ~(P1_U2390 & P1_U4791); 
assign P1_U4831 = ~(P1_U4786 & P1_INSTQUEUE_REG_11__0__SCAN_IN); 
assign P1_U4852 = ~(P1_U2397 & P1_U4848); 
assign P1_U4853 = ~(P1_U4843 & P1_INSTQUEUE_REG_10__7__SCAN_IN); 
assign P1_U4857 = ~(P1_U2396 & P1_U4848); 
assign P1_U4858 = ~(P1_U4843 & P1_INSTQUEUE_REG_10__6__SCAN_IN); 
assign P1_U4862 = ~(P1_U2395 & P1_U4848); 
assign P1_U4863 = ~(P1_U4843 & P1_INSTQUEUE_REG_10__5__SCAN_IN); 
assign P1_U4867 = ~(P1_U2394 & P1_U4848); 
assign P1_U4868 = ~(P1_U4843 & P1_INSTQUEUE_REG_10__4__SCAN_IN); 
assign P1_U4872 = ~(P1_U2393 & P1_U4848); 
assign P1_U4873 = ~(P1_U4843 & P1_INSTQUEUE_REG_10__3__SCAN_IN); 
assign P1_U4877 = ~(P1_U2392 & P1_U4848); 
assign P1_U4878 = ~(P1_U4843 & P1_INSTQUEUE_REG_10__2__SCAN_IN); 
assign P1_U4882 = ~(P1_U2391 & P1_U4848); 
assign P1_U4883 = ~(P1_U4843 & P1_INSTQUEUE_REG_10__1__SCAN_IN); 
assign P1_U4887 = ~(P1_U2390 & P1_U4848); 
assign P1_U4888 = ~(P1_U4843 & P1_INSTQUEUE_REG_10__0__SCAN_IN); 
assign P1_U4910 = ~(P1_U2397 & P1_U4906); 
assign P1_U4911 = ~(P1_U4901 & P1_INSTQUEUE_REG_9__7__SCAN_IN); 
assign P1_U4915 = ~(P1_U2396 & P1_U4906); 
assign P1_U4916 = ~(P1_U4901 & P1_INSTQUEUE_REG_9__6__SCAN_IN); 
assign P1_U4920 = ~(P1_U2395 & P1_U4906); 
assign P1_U4921 = ~(P1_U4901 & P1_INSTQUEUE_REG_9__5__SCAN_IN); 
assign P1_U4925 = ~(P1_U2394 & P1_U4906); 
assign P1_U4926 = ~(P1_U4901 & P1_INSTQUEUE_REG_9__4__SCAN_IN); 
assign P1_U4930 = ~(P1_U2393 & P1_U4906); 
assign P1_U4931 = ~(P1_U4901 & P1_INSTQUEUE_REG_9__3__SCAN_IN); 
assign P1_U4935 = ~(P1_U2392 & P1_U4906); 
assign P1_U4936 = ~(P1_U4901 & P1_INSTQUEUE_REG_9__2__SCAN_IN); 
assign P1_U4940 = ~(P1_U2391 & P1_U4906); 
assign P1_U4941 = ~(P1_U4901 & P1_INSTQUEUE_REG_9__1__SCAN_IN); 
assign P1_U4945 = ~(P1_U2390 & P1_U4906); 
assign P1_U4946 = ~(P1_U4901 & P1_INSTQUEUE_REG_9__0__SCAN_IN); 
assign P1_U4967 = ~(P1_U2397 & P1_U4963); 
assign P1_U4968 = ~(P1_U4958 & P1_INSTQUEUE_REG_8__7__SCAN_IN); 
assign P1_U4972 = ~(P1_U2396 & P1_U4963); 
assign P1_U4973 = ~(P1_U4958 & P1_INSTQUEUE_REG_8__6__SCAN_IN); 
assign P1_U4977 = ~(P1_U2395 & P1_U4963); 
assign P1_U4978 = ~(P1_U4958 & P1_INSTQUEUE_REG_8__5__SCAN_IN); 
assign P1_U4982 = ~(P1_U2394 & P1_U4963); 
assign P1_U4983 = ~(P1_U4958 & P1_INSTQUEUE_REG_8__4__SCAN_IN); 
assign P1_U4987 = ~(P1_U2393 & P1_U4963); 
assign P1_U4988 = ~(P1_U4958 & P1_INSTQUEUE_REG_8__3__SCAN_IN); 
assign P1_U4992 = ~(P1_U2392 & P1_U4963); 
assign P1_U4993 = ~(P1_U4958 & P1_INSTQUEUE_REG_8__2__SCAN_IN); 
assign P1_U4997 = ~(P1_U2391 & P1_U4963); 
assign P1_U4998 = ~(P1_U4958 & P1_INSTQUEUE_REG_8__1__SCAN_IN); 
assign P1_U5002 = ~(P1_U2390 & P1_U4963); 
assign P1_U5003 = ~(P1_U4958 & P1_INSTQUEUE_REG_8__0__SCAN_IN); 
assign P1_U5014 = ~(P1_U5011 & P1_U3659); 
assign P1_U5019 = ~(P1_U5018 & P1_U5017); 
assign P1_U5071 = ~(P1_U5068 & P1_U3668); 
assign P1_U5076 = ~(P1_U5075 & P1_U5074); 
assign P1_U5129 = ~(P1_U5126 & P1_U3677); 
assign P1_U5134 = ~(P1_U5133 & P1_U5132); 
assign P1_U5186 = ~(P1_U5183 & P1_U3686); 
assign P1_U5191 = ~(P1_U5190 & P1_U5189); 
assign P1_U5244 = ~(P1_U5241 & P1_U3695); 
assign P1_U5249 = ~(P1_U5248 & P1_U5247); 
assign P1_U5301 = ~(P1_U5298 & P1_U3704); 
assign P1_U5306 = ~(P1_U5305 & P1_U5304); 
assign P1_U5359 = ~(P1_U5356 & P1_U3713); 
assign P1_U5364 = ~(P1_U5363 & P1_U5362); 
assign P1_U5416 = ~(P1_U5413 & P1_U3722); 
assign P1_U5421 = ~(P1_U5420 & P1_U5419); 
assign P1_U5731 = ~(P1_R2099_U72 & P1_U2380); 
assign P1_U5741 = ~(P1_ADD_405_U66 & P1_U2375); 
assign P1_U5742 = ~(P1_ADD_515_U65 & P1_U2374); 
assign P1_U5827 = ~(P1_R2358_U82 & P1_U2364); 
assign P1_U5842 = ~(P1_R2358_U80 & P1_U2364); 
assign P1_U5919 = ~(P1_R2337_U77 & P1_U2376); 
assign P1_U6170 = ~(P1_U2386 & P1_R2358_U82); 
assign P1_U6179 = ~(P1_U2386 & P1_R2358_U80); 
assign P1_U6280 = ~(P1_U2383 & P1_R2358_U82); 
assign P1_U6289 = ~(P1_U2383 & P1_R2358_U80); 
assign P1_U6335 = ~(P1_U2371 & P1_R2099_U72); 
assign P1_U6535 = ~(P1_U2604 & P1_R2099_U72); 
assign P1_U6543 = ~(P1_R2096_U77 & P1_U7485); 
assign P1_U6803 = ~(P1_R2337_U77 & P1_U2352); 
assign P3_ADD_476_U52 = ~(P3_ADD_476_U116 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_476_U152 = ~(P3_ADD_476_U116 & P3_ADD_476_U51); 
assign P3_ADD_531_U53 = ~(P3_ADD_531_U120 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_531_U159 = ~(P3_ADD_531_U120 & P3_ADD_531_U52); 
assign P3_SUB_320_U42 = ~P3_ADD_318_U77; 
assign P3_SUB_320_U68 = P3_SUB_320_U145 & P3_SUB_320_U144; 
assign P3_SUB_320_U112 = ~(P3_ADD_318_U77 & P3_SUB_320_U111); 
assign P3_ADD_318_U52 = ~(P3_ADD_318_U116 & P3_PHYADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_318_U152 = ~(P3_ADD_318_U116 & P3_ADD_318_U51); 
assign P3_ADD_315_U52 = ~(P3_ADD_315_U113 & P3_PHYADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_315_U144 = ~(P3_ADD_315_U113 & P3_ADD_315_U51); 
assign P3_ADD_360_1242_U79 = ~(P3_ADD_360_1242_U241 & P3_ADD_360_1242_U240); 
assign P3_ADD_360_1242_U162 = ~P3_ADD_360_1242_U66; 
assign P3_ADD_360_1242_U169 = ~(P3_ADD_360_1242_U67 & P3_ADD_360_1242_U66); 
assign P3_ADD_360_1242_U171 = ~(P3_ADD_360_1242_U64 & P3_ADD_360_1242_U170); 
assign P3_ADD_467_U52 = ~(P3_ADD_467_U116 & P3_REIP_REG_25__SCAN_IN); 
assign P3_ADD_467_U152 = ~(P3_ADD_467_U116 & P3_ADD_467_U51); 
assign P3_ADD_430_U52 = ~(P3_ADD_430_U116 & P3_REIP_REG_25__SCAN_IN); 
assign P3_ADD_430_U152 = ~(P3_ADD_430_U116 & P3_ADD_430_U51); 
assign P3_ADD_380_U53 = ~(P3_ADD_380_U120 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_380_U159 = ~(P3_ADD_380_U120 & P3_ADD_380_U52); 
assign P3_ADD_344_U53 = ~(P3_ADD_344_U120 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_344_U159 = ~(P3_ADD_344_U120 & P3_ADD_344_U52); 
assign P3_ADD_339_U52 = ~(P3_ADD_339_U116 & P3_PHYADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_339_U152 = ~(P3_ADD_339_U116 & P3_ADD_339_U51); 
assign P3_ADD_541_U52 = ~(P3_ADD_541_U116 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_541_U152 = ~(P3_ADD_541_U116 & P3_ADD_541_U51); 
assign P3_SUB_357_1258_U77 = ~(P3_SUB_357_1258_U361 & P3_SUB_357_1258_U360); 
assign P3_SUB_357_1258_U225 = ~(P3_SUB_357_1258_U354 & P3_SUB_357_1258_U353 & P3_SUB_357_1258_U294); 
assign P3_ADD_515_U52 = ~(P3_ADD_515_U116 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_515_U152 = ~(P3_ADD_515_U116 & P3_ADD_515_U51); 
assign P3_ADD_394_U52 = ~(P3_ADD_394_U119 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_394_U154 = ~(P3_ADD_394_U119 & P3_ADD_394_U51); 
assign P3_ADD_441_U52 = ~(P3_ADD_441_U116 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_441_U152 = ~(P3_ADD_441_U116 & P3_ADD_441_U51); 
assign P3_ADD_349_U53 = ~(P3_ADD_349_U120 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_349_U159 = ~(P3_ADD_349_U120 & P3_ADD_349_U52); 
assign P3_ADD_405_U52 = ~(P3_ADD_405_U119 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_405_U154 = ~(P3_ADD_405_U119 & P3_ADD_405_U51); 
assign P3_ADD_553_U53 = ~(P3_ADD_553_U120 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_553_U159 = ~(P3_ADD_553_U120 & P3_ADD_553_U52); 
assign P3_ADD_558_U53 = ~(P3_ADD_558_U120 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_558_U159 = ~(P3_ADD_558_U120 & P3_ADD_558_U52); 
assign P3_ADD_385_U53 = ~(P3_ADD_385_U120 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_385_U159 = ~(P3_ADD_385_U120 & P3_ADD_385_U52); 
assign P3_ADD_547_U53 = ~(P3_ADD_547_U120 & P3_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P3_ADD_547_U159 = ~(P3_ADD_547_U120 & P3_ADD_547_U52); 
assign P3_ADD_371_1212_U14 = P3_ADD_371_1212_U181 & P3_ADD_371_1212_U68; 
assign P3_ADD_371_1212_U70 = ~(P3_ADD_371_1212_U171 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_494_U52 = ~(P3_ADD_494_U116 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_494_U152 = ~(P3_ADD_494_U116 & P3_ADD_494_U51); 
assign P3_ADD_536_U52 = ~(P3_ADD_536_U116 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_536_U152 = ~(P3_ADD_536_U116 & P3_ADD_536_U51); 
assign P2_R2099_U89 = ~(P2_R2099_U215 & P2_R2099_U214); 
assign P2_R2099_U130 = ~P2_R2099_U35; 
assign P2_R2099_U212 = ~(P2_U2732 & P2_R2099_U35); 
assign P2_ADD_391_1196_U36 = ~(P2_ADD_391_1196_U35 & P2_ADD_391_1196_U193); 
assign P2_ADD_391_1196_U40 = ~P2_R2182_U91; 
assign P2_ADD_391_1196_U67 = ~P2_R2096_U85; 
assign P2_ADD_391_1196_U88 = ~(P2_ADD_391_1196_U315 & P2_ADD_391_1196_U314); 
assign P2_ADD_391_1196_U154 = P2_ADD_391_1196_U462 & P2_ADD_391_1196_U461; 
assign P2_ADD_391_1196_U191 = ~P2_ADD_391_1196_U35; 
assign P2_ADD_391_1196_U223 = P2_R2096_U92 | P2_R2182_U91; 
assign P2_ADD_391_1196_U226 = ~(P2_R2096_U92 & P2_R2182_U91); 
assign P2_ADD_391_1196_U291 = ~(P2_R2096_U92 & P2_R2182_U91); 
assign P2_ADD_391_1196_U304 = ~(P2_ADD_391_1196_U293 & P2_ADD_391_1196_U159); 
assign P2_ADD_391_1196_U455 = ~(P2_R2182_U91 & P2_ADD_391_1196_U41); 
assign P2_ADD_391_1196_U456 = ~(P2_R2096_U93 & P2_ADD_391_1196_U42); 
assign P2_R2182_U12 = P2_U2694 & P2_R2182_U18; 
assign P2_R2182_U90 = ~(P2_R2182_U291 & P2_R2182_U290); 
assign P2_R2182_U149 = ~P2_R2182_U18; 
assign P2_R2182_U286 = ~(P2_R2182_U29 & P2_R2182_U18); 
assign P2_R2182_U289 = ~(P2_R2182_U148 & P2_U2695); 
assign P2_R2027_U53 = ~(P2_R2027_U120 & P2_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P2_R2027_U159 = ~(P2_R2027_U120 & P2_R2027_U52); 
assign P2_R2337_U53 = ~(P2_R2337_U117 & P2_PHYADDRPOINTER_REG_26__SCAN_IN); 
assign P2_R2337_U150 = ~(P2_R2337_U117 & P2_R2337_U52); 
assign P2_R2096_U12 = P2_U2624 & P2_R2096_U11; 
assign P2_R2096_U84 = ~(P2_R2096_U232 & P2_R2096_U231); 
assign P2_R2096_U160 = ~P2_R2096_U11; 
assign P2_R2096_U227 = ~(P2_R2096_U43 & P2_R2096_U11); 
assign P2_R2096_U230 = ~(P2_R2096_U159 & P2_U2625); 
assign P2_R2256_U19 = ~(P2_R2256_U52 & P2_R2256_U51); 
assign P2_R2256_U43 = ~P2_R2256_U14; 
assign P2_R2256_U49 = ~(P2_U3623 & P2_R2256_U14); 
assign P2_R1957_U41 = ~P2_U3666; 
assign P2_R1957_U68 = P2_R1957_U145 & P2_R1957_U144; 
assign P2_R1957_U112 = ~(P2_U3666 & P2_R1957_U111); 
assign P2_R2278_U6 = ~(P2_R2278_U490 & P2_R2278_U489 & P2_R2278_U345); 
assign P2_R2278_U11 = ~P2_U3635; 
assign P2_R2278_U62 = ~P2_U2802; 
assign P2_R2278_U128 = P2_R2278_U328 & P2_R2278_U264; 
assign P2_R2278_U158 = ~(P2_R2278_U20 & P2_R2278_U211); 
assign P2_R2278_U164 = P2_R2278_U410 & P2_R2278_U409; 
assign P2_R2278_U189 = P2_R2278_U506 & P2_R2278_U505; 
assign P2_R2278_U214 = P2_U3635 | P2_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P2_R2278_U215 = ~(P2_U3635 & P2_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P2_R2278_U270 = P2_U2802 | P2_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P2_R2278_U271 = ~(P2_U2802 & P2_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P2_R2278_U314 = P2_U3635 | P2_INSTADDRPOINTER_REG_3__SCAN_IN; 
assign P2_R2278_U331 = P2_U2802 | P2_INSTADDRPOINTER_REG_19__SCAN_IN; 
assign P2_R2278_U389 = ~(P2_U3635 & P2_R2278_U12); 
assign P2_R2278_U391 = ~(P2_U3635 & P2_R2278_U12); 
assign P2_R2278_U413 = ~(P2_R2278_U412 & P2_R2278_U411); 
assign P2_R2278_U492 = ~(P2_U2802 & P2_R2278_U63); 
assign P2_R2278_U494 = ~(P2_U2802 & P2_R2278_U63); 
assign P2_R2278_U498 = ~(P2_R2278_U64 & P2_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P2_R2278_U500 = ~(P2_R2278_U64 & P2_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P2_R2278_U509 = ~(P2_R2278_U508 & P2_R2278_U507); 
assign P2_ADD_394_U52 = ~(P2_ADD_394_U119 & P2_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P2_ADD_394_U184 = ~(P2_ADD_394_U119 & P2_ADD_394_U51); 
assign P2_R2267_U11 = P2_R2267_U123 & P2_R2267_U36; 
assign P2_R2267_U37 = ~(P2_R2267_U51 & P2_R2267_U107); 
assign P2_R2267_U120 = ~(P2_R2267_U107 & P2_R2267_U72); 
assign P2_R2267_U152 = ~(P2_R2267_U107 & P2_R2267_U72); 
assign P2_ADD_371_1212_U129 = P2_ADD_371_1212_U259 & P2_ADD_371_1212_U258; 
assign P2_ADD_371_1212_U130 = ~(P2_ADD_371_1212_U143 & P2_ADD_371_1212_U142); 
assign P2_ADD_371_1212_U226 = ~(P2_ADD_371_1212_U140 & P2_ADD_371_1212_U224); 
assign P2_ADD_371_1212_U233 = ~(P2_ADD_371_1212_U35 & P2_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P2_ADD_371_1212_U235 = ~(P2_ADD_371_1212_U35 & P2_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P2_ADD_371_1212_U262 = ~(P2_ADD_371_1212_U261 & P2_ADD_371_1212_U260); 
assign P1_R2278_U139 = P1_R2278_U357 & P1_R2278_U140; 
assign P1_R2278_U173 = P1_R2278_U589 & P1_R2278_U588 & P1_R2278_U285; 
assign P1_R2278_U174 = P1_R2278_U337 & P1_R2278_U227; 
assign P1_R2278_U251 = ~P1_R2278_U40; 
assign P1_R2278_U265 = ~(P1_R2278_U264 & P1_R2278_U40); 
assign P1_R2278_U272 = ~(P1_R2278_U249 & P1_R2278_U271); 
assign P1_R2278_U398 = ~(P1_R2278_U386 & P1_R2278_U324); 
assign P1_R2278_U401 = ~P1_R2278_U87; 
assign P1_R2278_U403 = ~(P1_R2278_U380 & P1_R2278_U324); 
assign P1_R2278_U404 = ~(P1_R2278_U384 & P1_R2278_U324); 
assign P1_R2278_U406 = ~(P1_R2278_U387 & P1_R2278_U324); 
assign P1_R2278_U407 = ~(P1_R2278_U87 & P1_R2278_U324); 
assign P1_R2278_U409 = ~(P1_R2278_U408 & P1_R2278_U319); 
assign P1_R2278_U410 = ~(P1_R2278_U402 & P1_R2278_U227); 
assign P1_R2278_U412 = ~(P1_R2278_U390 & P1_R2278_U227); 
assign P1_R2278_U415 = ~(P1_R2278_U287 & P1_R2278_U227); 
assign P1_R2278_U417 = ~(P1_R2278_U382 & P1_R2278_U227); 
assign P1_R2278_U444 = ~(P1_R2278_U347 & P1_R2278_U40); 
assign P1_R2358_U7 = P1_R2358_U6 & P1_R2358_U282; 
assign P1_R2358_U73 = ~(P1_R2358_U233 & P1_R2358_U321); 
assign P1_R2358_U126 = P1_R2358_U258 & P1_R2358_U259 & P1_R2358_U255 & P1_R2358_U356; 
assign P1_R2358_U139 = P1_R2358_U257 & P1_R2358_U256; 
assign P1_R2358_U238 = ~P1_R2358_U36; 
assign P1_R2358_U239 = ~(P1_R2358_U36 & P1_R2358_U215); 
assign P1_R2358_U242 = ~(P1_R2358_U36 & P1_R2358_U215 & P1_R2358_U241); 
assign P1_R2358_U244 = ~(P1_R2358_U237 & P1_R2358_U243); 
assign P1_R2358_U269 = ~P1_R2358_U199; 
assign P1_R2358_U283 = ~(P1_U2629 & P1_R2358_U515); 
assign P1_R2358_U309 = ~(P1_R2358_U199 & P1_R2358_U259); 
assign P1_R2358_U316 = ~(P1_R2358_U257 & P1_R2358_U256); 
assign P1_R2358_U353 = ~(P1_R2358_U270 & P1_R2358_U258 & P1_R2358_U255 & P1_R2358_U257); 
assign P1_R2358_U354 = ~(P1_R2358_U260 & P1_R2358_U255 & P1_R2358_U257); 
assign P1_R2358_U355 = ~(P1_R2358_U261 & P1_R2358_U257); 
assign P1_R2358_U364 = ~(P1_R2358_U363 & P1_R2358_U282); 
assign P1_R2358_U450 = ~(P1_R2358_U77 & P1_R2358_U231); 
assign P1_R2358_U502 = ~(P1_U2352 & P1_R2358_U166); 
assign P1_R2358_U510 = ~(P1_U2352 & P1_R2358_U166); 
assign P1_R2358_U608 = ~(P1_R2358_U352 & P1_R2358_U199); 
assign P1_R2099_U21 = ~(P1_R2099_U175 & P1_R2099_U49); 
assign P1_R2099_U308 = ~(P1_R2099_U240 & P1_R2099_U175); 
assign P1_R2337_U52 = ~(P1_R2337_U116 & P1_PHYADDRPOINTER_REG_25__SCAN_IN); 
assign P1_R2337_U152 = ~(P1_R2337_U116 & P1_R2337_U51); 
assign P1_R2096_U52 = ~(P1_R2096_U116 & P1_REIP_REG_25__SCAN_IN); 
assign P1_R2096_U152 = ~(P1_R2096_U116 & P1_R2096_U51); 
assign P1_ADD_405_U52 = ~(P1_ADD_405_U119 & P1_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P1_ADD_405_U184 = ~(P1_ADD_405_U119 & P1_ADD_405_U51); 
assign P1_ADD_515_U52 = ~(P1_ADD_515_U116 & P1_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P1_ADD_515_U180 = ~(P1_ADD_515_U116 & P1_ADD_515_U51); 
assign P3_U2807 = ~(P3_U6590 & P3_U6589 & P3_U6592 & P3_U6591 & P3_U3977); 
assign P3_U3864 = P3_U6188 & P3_U6187; 
assign P3_U3866 = P3_U6190 & P3_U6189 & P3_U6191 & P3_U3865; 
assign P3_U3870 = P3_U6200 & P3_U6199 & P3_U6201; 
assign P3_U3871 = P3_U6203 & P3_U6202; 
assign P3_U3875 = P3_U6217 & P3_U6216; 
assign P3_U3878 = P3_U6219 & P3_U6218 & P3_U6220; 
assign P3_U3879 = P3_U6222 & P3_U6221; 
assign P3_U3978 = P3_U6604 & P3_U6601 & P3_U6602 & P3_U6603; 
assign P3_U4111 = P3_U7302 & P3_U7301; 
assign P3_U6134 = ~(P3_U4318 & P3_U6132); 
assign P3_U6158 = ~(P3_U4318 & P3_U6156); 
assign P3_U6180 = ~(P3_U3862 & P3_U3857); 
assign P3_U6208 = ~(P3_ADD_360_1242_U79 & P3_U2395); 
assign P3_U6251 = ~(P3_ADD_371_1212_U14 & P3_U2360); 
assign P3_U6353 = ~(P3_SUB_357_1258_U77 & P3_U2393); 
assign P3_U6599 = ~(P3_U2396 & P3_ADD_360_1242_U79); 
assign P3_U6611 = ~(P3_U2387 & P3_ADD_371_1212_U14); 
assign P3_U6648 = ~(P3_U2394 & P3_SUB_357_1258_U77); 
assign P2_U2800 = P2_U3242 & P2_R2267_U11; 
assign P2_U2912 = ~(P2_U4066 & P2_U6355 & P2_U6356); 
assign P2_U3665 = ~(P2_U8386 & P2_U8385); 
assign P2_U6360 = ~(P2_ADD_391_1196_U88 & P2_U2397); 
assign P2_U6429 = ~(P2_U2380 & P2_R2096_U84); 
assign P2_U6514 = ~(P2_U2379 & P2_R2099_U89); 
assign P2_U6519 = ~(P2_R2182_U90 & P2_U2393); 
assign P2_U6694 = ~(P2_U2392 & P2_R2099_U89); 
assign P2_U6747 = ~(P2_R2267_U11 & P2_U2587); 
assign P2_U6764 = ~(P2_U2588 & P2_R2096_U84); 
assign P2_U8319 = ~(P2_R2256_U19 & P2_U3572); 
assign P1_U2864 = ~(P1_U6290 & P1_U6291 & P1_U6289); 
assign P1_U2867 = ~(P1_U6281 & P1_U6282 & P1_U6280); 
assign P1_U2896 = ~(P1_U6180 & P1_U6178 & P1_U6179); 
assign P1_U2899 = ~(P1_U6171 & P1_U6169 & P1_U6170); 
assign P1_U3097 = ~(P1_U5003 & P1_U5002 & P1_U3658); 
assign P1_U3098 = ~(P1_U4998 & P1_U4997 & P1_U3657); 
assign P1_U3099 = ~(P1_U4993 & P1_U4992 & P1_U3656); 
assign P1_U3100 = ~(P1_U4988 & P1_U4987 & P1_U3655); 
assign P1_U3101 = ~(P1_U4983 & P1_U4982 & P1_U3654); 
assign P1_U3102 = ~(P1_U4978 & P1_U4977 & P1_U3653); 
assign P1_U3103 = ~(P1_U4973 & P1_U4972 & P1_U3652); 
assign P1_U3104 = ~(P1_U4968 & P1_U4967 & P1_U3651); 
assign P1_U3105 = ~(P1_U4946 & P1_U4945 & P1_U3649); 
assign P1_U3106 = ~(P1_U4941 & P1_U4940 & P1_U3648); 
assign P1_U3107 = ~(P1_U4936 & P1_U4935 & P1_U3647); 
assign P1_U3108 = ~(P1_U4931 & P1_U4930 & P1_U3646); 
assign P1_U3109 = ~(P1_U4926 & P1_U4925 & P1_U3645); 
assign P1_U3110 = ~(P1_U4921 & P1_U4920 & P1_U3644); 
assign P1_U3111 = ~(P1_U4916 & P1_U4915 & P1_U3643); 
assign P1_U3112 = ~(P1_U4911 & P1_U4910 & P1_U3642); 
assign P1_U3113 = ~(P1_U4888 & P1_U4887 & P1_U3640); 
assign P1_U3114 = ~(P1_U4883 & P1_U4882 & P1_U3639); 
assign P1_U3115 = ~(P1_U4878 & P1_U4877 & P1_U3638); 
assign P1_U3116 = ~(P1_U4873 & P1_U4872 & P1_U3637); 
assign P1_U3117 = ~(P1_U4868 & P1_U4867 & P1_U3636); 
assign P1_U3118 = ~(P1_U4863 & P1_U4862 & P1_U3635); 
assign P1_U3119 = ~(P1_U4858 & P1_U4857 & P1_U3634); 
assign P1_U3120 = ~(P1_U4853 & P1_U4852 & P1_U3633); 
assign P1_U3121 = ~(P1_U4831 & P1_U4830 & P1_U3631); 
assign P1_U3122 = ~(P1_U4826 & P1_U4825 & P1_U3630); 
assign P1_U3123 = ~(P1_U4821 & P1_U4820 & P1_U3629); 
assign P1_U3124 = ~(P1_U4816 & P1_U4815 & P1_U3628); 
assign P1_U3125 = ~(P1_U4811 & P1_U4810 & P1_U3627); 
assign P1_U3126 = ~(P1_U4806 & P1_U4805 & P1_U3626); 
assign P1_U3127 = ~(P1_U4801 & P1_U4800 & P1_U3625); 
assign P1_U3128 = ~(P1_U4796 & P1_U4795 & P1_U3624); 
assign P1_U3129 = ~(P1_U4773 & P1_U4772 & P1_U3622); 
assign P1_U3130 = ~(P1_U4768 & P1_U4767 & P1_U3621); 
assign P1_U3131 = ~(P1_U4763 & P1_U4762 & P1_U3620); 
assign P1_U3132 = ~(P1_U4758 & P1_U4757 & P1_U3619); 
assign P1_U3133 = ~(P1_U4753 & P1_U4752 & P1_U3618); 
assign P1_U3134 = ~(P1_U4748 & P1_U4747 & P1_U3617); 
assign P1_U3135 = ~(P1_U4743 & P1_U4742 & P1_U3616); 
assign P1_U3136 = ~(P1_U4738 & P1_U4737 & P1_U3615); 
assign P1_U3137 = ~(P1_U4716 & P1_U4715 & P1_U3613); 
assign P1_U3138 = ~(P1_U4711 & P1_U4710 & P1_U3612); 
assign P1_U3139 = ~(P1_U4706 & P1_U4705 & P1_U3611); 
assign P1_U3140 = ~(P1_U4701 & P1_U4700 & P1_U3610); 
assign P1_U3141 = ~(P1_U4696 & P1_U4695 & P1_U3609); 
assign P1_U3142 = ~(P1_U4691 & P1_U4690 & P1_U3608); 
assign P1_U3143 = ~(P1_U4686 & P1_U4685 & P1_U3607); 
assign P1_U3144 = ~(P1_U4681 & P1_U4680 & P1_U3606); 
assign P1_U3145 = ~(P1_U4657 & P1_U4656 & P1_U3604); 
assign P1_U3146 = ~(P1_U4652 & P1_U4651 & P1_U3603); 
assign P1_U3147 = ~(P1_U4647 & P1_U4646 & P1_U3602); 
assign P1_U3148 = ~(P1_U4642 & P1_U4641 & P1_U3601); 
assign P1_U3149 = ~(P1_U4637 & P1_U4636 & P1_U3600); 
assign P1_U3150 = ~(P1_U4632 & P1_U4631 & P1_U3599); 
assign P1_U3151 = ~(P1_U4627 & P1_U4626 & P1_U3598); 
assign P1_U3152 = ~(P1_U4622 & P1_U4621 & P1_U3597); 
assign P1_U3153 = ~(P1_U4599 & P1_U4598 & P1_U3595); 
assign P1_U3154 = ~(P1_U4594 & P1_U4593 & P1_U3594); 
assign P1_U3155 = ~(P1_U4589 & P1_U4588 & P1_U3593); 
assign P1_U3156 = ~(P1_U4584 & P1_U4583 & P1_U3592); 
assign P1_U3157 = ~(P1_U4579 & P1_U4578 & P1_U3591); 
assign P1_U3158 = ~(P1_U4574 & P1_U4573 & P1_U3590); 
assign P1_U3159 = ~(P1_U4569 & P1_U4568 & P1_U3589); 
assign P1_U3160 = ~(P1_U4564 & P1_U4563 & P1_U3588); 
assign P1_U3838 = P1_U5739 & P1_U5741; 
assign P1_U3840 = P1_U3839 & P1_U5742; 
assign P1_U3934 = P1_U6545 & P1_U6543; 
assign P1_U4016 = P1_U6801 & P1_U6802 & P1_U6803; 
assign P1_U5023 = ~(P1_U2397 & P1_U5019); 
assign P1_U5024 = ~(P1_U5014 & P1_INSTQUEUE_REG_7__7__SCAN_IN); 
assign P1_U5028 = ~(P1_U2396 & P1_U5019); 
assign P1_U5029 = ~(P1_U5014 & P1_INSTQUEUE_REG_7__6__SCAN_IN); 
assign P1_U5033 = ~(P1_U2395 & P1_U5019); 
assign P1_U5034 = ~(P1_U5014 & P1_INSTQUEUE_REG_7__5__SCAN_IN); 
assign P1_U5038 = ~(P1_U2394 & P1_U5019); 
assign P1_U5039 = ~(P1_U5014 & P1_INSTQUEUE_REG_7__4__SCAN_IN); 
assign P1_U5043 = ~(P1_U2393 & P1_U5019); 
assign P1_U5044 = ~(P1_U5014 & P1_INSTQUEUE_REG_7__3__SCAN_IN); 
assign P1_U5048 = ~(P1_U2392 & P1_U5019); 
assign P1_U5049 = ~(P1_U5014 & P1_INSTQUEUE_REG_7__2__SCAN_IN); 
assign P1_U5053 = ~(P1_U2391 & P1_U5019); 
assign P1_U5054 = ~(P1_U5014 & P1_INSTQUEUE_REG_7__1__SCAN_IN); 
assign P1_U5058 = ~(P1_U2390 & P1_U5019); 
assign P1_U5059 = ~(P1_U5014 & P1_INSTQUEUE_REG_7__0__SCAN_IN); 
assign P1_U5080 = ~(P1_U2397 & P1_U5076); 
assign P1_U5081 = ~(P1_U5071 & P1_INSTQUEUE_REG_6__7__SCAN_IN); 
assign P1_U5085 = ~(P1_U2396 & P1_U5076); 
assign P1_U5086 = ~(P1_U5071 & P1_INSTQUEUE_REG_6__6__SCAN_IN); 
assign P1_U5090 = ~(P1_U2395 & P1_U5076); 
assign P1_U5091 = ~(P1_U5071 & P1_INSTQUEUE_REG_6__5__SCAN_IN); 
assign P1_U5095 = ~(P1_U2394 & P1_U5076); 
assign P1_U5096 = ~(P1_U5071 & P1_INSTQUEUE_REG_6__4__SCAN_IN); 
assign P1_U5100 = ~(P1_U2393 & P1_U5076); 
assign P1_U5101 = ~(P1_U5071 & P1_INSTQUEUE_REG_6__3__SCAN_IN); 
assign P1_U5105 = ~(P1_U2392 & P1_U5076); 
assign P1_U5106 = ~(P1_U5071 & P1_INSTQUEUE_REG_6__2__SCAN_IN); 
assign P1_U5110 = ~(P1_U2391 & P1_U5076); 
assign P1_U5111 = ~(P1_U5071 & P1_INSTQUEUE_REG_6__1__SCAN_IN); 
assign P1_U5115 = ~(P1_U2390 & P1_U5076); 
assign P1_U5116 = ~(P1_U5071 & P1_INSTQUEUE_REG_6__0__SCAN_IN); 
assign P1_U5138 = ~(P1_U2397 & P1_U5134); 
assign P1_U5139 = ~(P1_U5129 & P1_INSTQUEUE_REG_5__7__SCAN_IN); 
assign P1_U5143 = ~(P1_U2396 & P1_U5134); 
assign P1_U5144 = ~(P1_U5129 & P1_INSTQUEUE_REG_5__6__SCAN_IN); 
assign P1_U5148 = ~(P1_U2395 & P1_U5134); 
assign P1_U5149 = ~(P1_U5129 & P1_INSTQUEUE_REG_5__5__SCAN_IN); 
assign P1_U5153 = ~(P1_U2394 & P1_U5134); 
assign P1_U5154 = ~(P1_U5129 & P1_INSTQUEUE_REG_5__4__SCAN_IN); 
assign P1_U5158 = ~(P1_U2393 & P1_U5134); 
assign P1_U5159 = ~(P1_U5129 & P1_INSTQUEUE_REG_5__3__SCAN_IN); 
assign P1_U5163 = ~(P1_U2392 & P1_U5134); 
assign P1_U5164 = ~(P1_U5129 & P1_INSTQUEUE_REG_5__2__SCAN_IN); 
assign P1_U5168 = ~(P1_U2391 & P1_U5134); 
assign P1_U5169 = ~(P1_U5129 & P1_INSTQUEUE_REG_5__1__SCAN_IN); 
assign P1_U5173 = ~(P1_U2390 & P1_U5134); 
assign P1_U5174 = ~(P1_U5129 & P1_INSTQUEUE_REG_5__0__SCAN_IN); 
assign P1_U5195 = ~(P1_U2397 & P1_U5191); 
assign P1_U5196 = ~(P1_U5186 & P1_INSTQUEUE_REG_4__7__SCAN_IN); 
assign P1_U5200 = ~(P1_U2396 & P1_U5191); 
assign P1_U5201 = ~(P1_U5186 & P1_INSTQUEUE_REG_4__6__SCAN_IN); 
assign P1_U5205 = ~(P1_U2395 & P1_U5191); 
assign P1_U5206 = ~(P1_U5186 & P1_INSTQUEUE_REG_4__5__SCAN_IN); 
assign P1_U5210 = ~(P1_U2394 & P1_U5191); 
assign P1_U5211 = ~(P1_U5186 & P1_INSTQUEUE_REG_4__4__SCAN_IN); 
assign P1_U5215 = ~(P1_U2393 & P1_U5191); 
assign P1_U5216 = ~(P1_U5186 & P1_INSTQUEUE_REG_4__3__SCAN_IN); 
assign P1_U5220 = ~(P1_U2392 & P1_U5191); 
assign P1_U5221 = ~(P1_U5186 & P1_INSTQUEUE_REG_4__2__SCAN_IN); 
assign P1_U5225 = ~(P1_U2391 & P1_U5191); 
assign P1_U5226 = ~(P1_U5186 & P1_INSTQUEUE_REG_4__1__SCAN_IN); 
assign P1_U5230 = ~(P1_U2390 & P1_U5191); 
assign P1_U5231 = ~(P1_U5186 & P1_INSTQUEUE_REG_4__0__SCAN_IN); 
assign P1_U5253 = ~(P1_U2397 & P1_U5249); 
assign P1_U5254 = ~(P1_U5244 & P1_INSTQUEUE_REG_3__7__SCAN_IN); 
assign P1_U5258 = ~(P1_U2396 & P1_U5249); 
assign P1_U5259 = ~(P1_U5244 & P1_INSTQUEUE_REG_3__6__SCAN_IN); 
assign P1_U5263 = ~(P1_U2395 & P1_U5249); 
assign P1_U5264 = ~(P1_U5244 & P1_INSTQUEUE_REG_3__5__SCAN_IN); 
assign P1_U5268 = ~(P1_U2394 & P1_U5249); 
assign P1_U5269 = ~(P1_U5244 & P1_INSTQUEUE_REG_3__4__SCAN_IN); 
assign P1_U5273 = ~(P1_U2393 & P1_U5249); 
assign P1_U5274 = ~(P1_U5244 & P1_INSTQUEUE_REG_3__3__SCAN_IN); 
assign P1_U5278 = ~(P1_U2392 & P1_U5249); 
assign P1_U5279 = ~(P1_U5244 & P1_INSTQUEUE_REG_3__2__SCAN_IN); 
assign P1_U5283 = ~(P1_U2391 & P1_U5249); 
assign P1_U5284 = ~(P1_U5244 & P1_INSTQUEUE_REG_3__1__SCAN_IN); 
assign P1_U5288 = ~(P1_U2390 & P1_U5249); 
assign P1_U5289 = ~(P1_U5244 & P1_INSTQUEUE_REG_3__0__SCAN_IN); 
assign P1_U5310 = ~(P1_U2397 & P1_U5306); 
assign P1_U5311 = ~(P1_U5301 & P1_INSTQUEUE_REG_2__7__SCAN_IN); 
assign P1_U5315 = ~(P1_U2396 & P1_U5306); 
assign P1_U5316 = ~(P1_U5301 & P1_INSTQUEUE_REG_2__6__SCAN_IN); 
assign P1_U5320 = ~(P1_U2395 & P1_U5306); 
assign P1_U5321 = ~(P1_U5301 & P1_INSTQUEUE_REG_2__5__SCAN_IN); 
assign P1_U5325 = ~(P1_U2394 & P1_U5306); 
assign P1_U5326 = ~(P1_U5301 & P1_INSTQUEUE_REG_2__4__SCAN_IN); 
assign P1_U5330 = ~(P1_U2393 & P1_U5306); 
assign P1_U5331 = ~(P1_U5301 & P1_INSTQUEUE_REG_2__3__SCAN_IN); 
assign P1_U5335 = ~(P1_U2392 & P1_U5306); 
assign P1_U5336 = ~(P1_U5301 & P1_INSTQUEUE_REG_2__2__SCAN_IN); 
assign P1_U5340 = ~(P1_U2391 & P1_U5306); 
assign P1_U5341 = ~(P1_U5301 & P1_INSTQUEUE_REG_2__1__SCAN_IN); 
assign P1_U5345 = ~(P1_U2390 & P1_U5306); 
assign P1_U5346 = ~(P1_U5301 & P1_INSTQUEUE_REG_2__0__SCAN_IN); 
assign P1_U5368 = ~(P1_U2397 & P1_U5364); 
assign P1_U5369 = ~(P1_U5359 & P1_INSTQUEUE_REG_1__7__SCAN_IN); 
assign P1_U5373 = ~(P1_U2396 & P1_U5364); 
assign P1_U5374 = ~(P1_U5359 & P1_INSTQUEUE_REG_1__6__SCAN_IN); 
assign P1_U5378 = ~(P1_U2395 & P1_U5364); 
assign P1_U5379 = ~(P1_U5359 & P1_INSTQUEUE_REG_1__5__SCAN_IN); 
assign P1_U5383 = ~(P1_U2394 & P1_U5364); 
assign P1_U5384 = ~(P1_U5359 & P1_INSTQUEUE_REG_1__4__SCAN_IN); 
assign P1_U5388 = ~(P1_U2393 & P1_U5364); 
assign P1_U5389 = ~(P1_U5359 & P1_INSTQUEUE_REG_1__3__SCAN_IN); 
assign P1_U5393 = ~(P1_U2392 & P1_U5364); 
assign P1_U5394 = ~(P1_U5359 & P1_INSTQUEUE_REG_1__2__SCAN_IN); 
assign P1_U5398 = ~(P1_U2391 & P1_U5364); 
assign P1_U5399 = ~(P1_U5359 & P1_INSTQUEUE_REG_1__1__SCAN_IN); 
assign P1_U5403 = ~(P1_U2390 & P1_U5364); 
assign P1_U5404 = ~(P1_U5359 & P1_INSTQUEUE_REG_1__0__SCAN_IN); 
assign P1_U5425 = ~(P1_U2397 & P1_U5421); 
assign P1_U5426 = ~(P1_U5416 & P1_INSTQUEUE_REG_0__7__SCAN_IN); 
assign P1_U5430 = ~(P1_U2396 & P1_U5421); 
assign P1_U5431 = ~(P1_U5416 & P1_INSTQUEUE_REG_0__6__SCAN_IN); 
assign P1_U5435 = ~(P1_U2395 & P1_U5421); 
assign P1_U5436 = ~(P1_U5416 & P1_INSTQUEUE_REG_0__5__SCAN_IN); 
assign P1_U5440 = ~(P1_U2394 & P1_U5421); 
assign P1_U5444 = ~(P1_U2393 & P1_U5421); 
assign P1_U5445 = ~(P1_U5416 & P1_INSTQUEUE_REG_0__3__SCAN_IN); 
assign P1_U5449 = ~(P1_U2392 & P1_U5421); 
assign P1_U5450 = ~(P1_U5416 & P1_INSTQUEUE_REG_0__2__SCAN_IN); 
assign P1_U5454 = ~(P1_U2391 & P1_U5421); 
assign P1_U5455 = ~(P1_U5416 & P1_INSTQUEUE_REG_0__1__SCAN_IN); 
assign P1_U5459 = ~(P1_U2390 & P1_U5421); 
assign P1_U5460 = ~(P1_U5416 & P1_INSTQUEUE_REG_0__0__SCAN_IN); 
assign P1_U7612 = ~(P1_U5416 & P1_INSTQUEUE_REG_0__4__SCAN_IN); 
assign P3_ADD_476_U76 = ~(P3_ADD_476_U152 & P3_ADD_476_U151); 
assign P3_ADD_476_U117 = ~P3_ADD_476_U52; 
assign P3_ADD_476_U149 = ~(P3_ADD_476_U52 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_531_U80 = ~(P3_ADD_531_U159 & P3_ADD_531_U158); 
assign P3_ADD_531_U121 = ~P3_ADD_531_U53; 
assign P3_ADD_531_U156 = ~(P3_ADD_531_U53 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_SUB_320_U35 = ~(P3_SUB_320_U42 & P3_SUB_320_U67 & P3_SUB_320_U99); 
assign P3_ADD_318_U76 = ~(P3_ADD_318_U152 & P3_ADD_318_U151); 
assign P3_ADD_318_U117 = ~P3_ADD_318_U52; 
assign P3_ADD_318_U149 = ~(P3_ADD_318_U52 & P3_PHYADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_315_U72 = ~(P3_ADD_315_U144 & P3_ADD_315_U143); 
assign P3_ADD_315_U114 = ~P3_ADD_315_U52; 
assign P3_ADD_315_U141 = ~(P3_ADD_315_U52 & P3_PHYADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_360_1242_U13 = P3_ADD_360_1242_U171 & P3_ADD_360_1242_U66; 
assign P3_ADD_360_1242_U68 = ~(P3_ADD_360_1242_U162 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_467_U76 = ~(P3_ADD_467_U152 & P3_ADD_467_U151); 
assign P3_ADD_467_U117 = ~P3_ADD_467_U52; 
assign P3_ADD_467_U149 = ~(P3_ADD_467_U52 & P3_REIP_REG_26__SCAN_IN); 
assign P3_ADD_430_U76 = ~(P3_ADD_430_U152 & P3_ADD_430_U151); 
assign P3_ADD_430_U117 = ~P3_ADD_430_U52; 
assign P3_ADD_430_U149 = ~(P3_ADD_430_U52 & P3_REIP_REG_26__SCAN_IN); 
assign P3_ADD_380_U80 = ~(P3_ADD_380_U159 & P3_ADD_380_U158); 
assign P3_ADD_380_U121 = ~P3_ADD_380_U53; 
assign P3_ADD_380_U156 = ~(P3_ADD_380_U53 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_344_U80 = ~(P3_ADD_344_U159 & P3_ADD_344_U158); 
assign P3_ADD_344_U121 = ~P3_ADD_344_U53; 
assign P3_ADD_344_U156 = ~(P3_ADD_344_U53 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_339_U76 = ~(P3_ADD_339_U152 & P3_ADD_339_U151); 
assign P3_ADD_339_U117 = ~P3_ADD_339_U52; 
assign P3_ADD_339_U149 = ~(P3_ADD_339_U52 & P3_PHYADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_541_U76 = ~(P3_ADD_541_U152 & P3_ADD_541_U151); 
assign P3_ADD_541_U117 = ~P3_ADD_541_U52; 
assign P3_ADD_541_U149 = ~(P3_ADD_541_U52 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_SUB_357_1258_U20 = P3_SUB_357_1258_U225 & P3_SUB_357_1258_U296; 
assign P3_ADD_515_U76 = ~(P3_ADD_515_U152 & P3_ADD_515_U151); 
assign P3_ADD_515_U117 = ~P3_ADD_515_U52; 
assign P3_ADD_515_U149 = ~(P3_ADD_515_U52 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_394_U75 = ~(P3_ADD_394_U154 & P3_ADD_394_U153); 
assign P3_ADD_394_U120 = ~P3_ADD_394_U52; 
assign P3_ADD_394_U151 = ~(P3_ADD_394_U52 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_441_U76 = ~(P3_ADD_441_U152 & P3_ADD_441_U151); 
assign P3_ADD_441_U117 = ~P3_ADD_441_U52; 
assign P3_ADD_441_U149 = ~(P3_ADD_441_U52 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_349_U80 = ~(P3_ADD_349_U159 & P3_ADD_349_U158); 
assign P3_ADD_349_U121 = ~P3_ADD_349_U53; 
assign P3_ADD_349_U156 = ~(P3_ADD_349_U53 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_405_U75 = ~(P3_ADD_405_U154 & P3_ADD_405_U153); 
assign P3_ADD_405_U120 = ~P3_ADD_405_U52; 
assign P3_ADD_405_U151 = ~(P3_ADD_405_U52 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_553_U80 = ~(P3_ADD_553_U159 & P3_ADD_553_U158); 
assign P3_ADD_553_U121 = ~P3_ADD_553_U53; 
assign P3_ADD_553_U156 = ~(P3_ADD_553_U53 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_558_U80 = ~(P3_ADD_558_U159 & P3_ADD_558_U158); 
assign P3_ADD_558_U121 = ~P3_ADD_558_U53; 
assign P3_ADD_558_U156 = ~(P3_ADD_558_U53 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_385_U80 = ~(P3_ADD_385_U159 & P3_ADD_385_U158); 
assign P3_ADD_385_U121 = ~P3_ADD_385_U53; 
assign P3_ADD_385_U156 = ~(P3_ADD_385_U53 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_547_U80 = ~(P3_ADD_547_U159 & P3_ADD_547_U158); 
assign P3_ADD_547_U121 = ~P3_ADD_547_U53; 
assign P3_ADD_547_U156 = ~(P3_ADD_547_U53 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_371_1212_U15 = P3_ADD_371_1212_U179 & P3_ADD_371_1212_U70; 
assign P3_ADD_371_1212_U172 = ~P3_ADD_371_1212_U70; 
assign P3_ADD_371_1212_U245 = ~(P3_ADD_371_1212_U70 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_494_U76 = ~(P3_ADD_494_U152 & P3_ADD_494_U151); 
assign P3_ADD_494_U117 = ~P3_ADD_494_U52; 
assign P3_ADD_494_U149 = ~(P3_ADD_494_U52 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_536_U76 = ~(P3_ADD_536_U152 & P3_ADD_536_U151); 
assign P3_ADD_536_U117 = ~P3_ADD_536_U52; 
assign P3_ADD_536_U149 = ~(P3_ADD_536_U52 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P2_R2099_U37 = ~(P2_U2732 & P2_R2099_U130); 
assign P2_R2099_U213 = ~(P2_R2099_U130 & P2_R2099_U36); 
assign P2_ADD_391_1196_U50 = ~(P2_ADD_391_1196_U36 & P2_ADD_391_1196_U206); 
assign P2_ADD_391_1196_U54 = ~P2_R2182_U90; 
assign P2_ADD_391_1196_U69 = ~P2_R2096_U84; 
assign P2_ADD_391_1196_U192 = ~(P2_ADD_391_1196_U110 & P2_ADD_391_1196_U191); 
assign P2_ADD_391_1196_U194 = ~P2_ADD_391_1196_U36; 
assign P2_ADD_391_1196_U228 = P2_R2182_U90 | P2_R2096_U91; 
assign P2_ADD_391_1196_U230 = ~(P2_R2096_U91 & P2_R2182_U90); 
assign P2_ADD_391_1196_U448 = ~(P2_R2182_U90 & P2_ADD_391_1196_U55); 
assign P2_ADD_391_1196_U450 = ~(P2_R2182_U90 & P2_ADD_391_1196_U55); 
assign P2_ADD_391_1196_U454 = ~(P2_R2096_U92 & P2_ADD_391_1196_U40); 
assign P2_ADD_391_1196_U458 = ~(P2_ADD_391_1196_U457 & P2_ADD_391_1196_U456); 
assign P2_R2182_U13 = P2_U2693 & P2_R2182_U12; 
assign P2_R2182_U89 = ~(P2_R2182_U289 & P2_R2182_U288); 
assign P2_R2182_U150 = ~P2_R2182_U12; 
assign P2_R2182_U284 = ~(P2_R2182_U30 & P2_R2182_U12); 
assign P2_R2182_U287 = ~(P2_R2182_U149 & P2_U2694); 
assign P2_R2027_U80 = ~(P2_R2027_U159 & P2_R2027_U158); 
assign P2_R2027_U121 = ~P2_R2027_U53; 
assign P2_R2027_U156 = ~(P2_R2027_U53 & P2_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P2_R2337_U74 = ~(P2_R2337_U150 & P2_R2337_U149); 
assign P2_R2337_U118 = ~P2_R2337_U53; 
assign P2_R2337_U147 = ~(P2_R2337_U53 & P2_PHYADDRPOINTER_REG_27__SCAN_IN); 
assign P2_R2096_U15 = P2_U2623 & P2_R2096_U12; 
assign P2_R2096_U83 = ~(P2_R2096_U230 & P2_R2096_U229); 
assign P2_R2096_U161 = ~P2_R2096_U12; 
assign P2_R2096_U225 = ~(P2_R2096_U42 & P2_R2096_U12); 
assign P2_R2096_U228 = ~(P2_R2096_U160 & P2_U2624); 
assign P2_R2256_U5 = P2_R2256_U23 & P2_R2256_U43; 
assign P2_R2256_U24 = ~(P2_U3623 & P2_R2256_U43); 
assign P2_R2256_U50 = ~(P2_R2256_U43 & P2_R2256_U16); 
assign P2_R1957_U34 = ~(P2_R1957_U99 & P2_R1957_U67 & P2_R1957_U41); 
assign P2_R2278_U21 = ~P2_U3634; 
assign P2_R2278_U23 = ~(P2_U3634 & P2_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P2_R2278_U39 = ~P2_U2801; 
assign P2_R2278_U113 = P2_R2278_U210 & P2_R2278_U314; 
assign P2_R2278_U144 = P2_R2278_U266 & P2_R2278_U270; 
assign P2_R2278_U187 = P2_R2278_U499 & P2_R2278_U498; 
assign P2_R2278_U213 = ~P2_R2278_U158; 
assign P2_R2278_U217 = P2_U3634 | P2_INSTADDRPOINTER_REG_4__SCAN_IN; 
assign P2_R2278_U273 = P2_U2801 | P2_INSTADDRPOINTER_REG_20__SCAN_IN; 
assign P2_R2278_U274 = ~(P2_U2801 & P2_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P2_R2278_U313 = ~(P2_R2278_U212 & P2_R2278_U214); 
assign P2_R2278_U332 = ~(P2_R2278_U268 & P2_R2278_U271); 
assign P2_R2278_U382 = ~(P2_U3634 & P2_R2278_U22); 
assign P2_R2278_U384 = ~(P2_U3634 & P2_R2278_U22); 
assign P2_R2278_U388 = ~(P2_R2278_U11 & P2_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P2_R2278_U390 = ~(P2_R2278_U11 & P2_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P2_R2278_U414 = ~(P2_R2278_U164 & P2_R2278_U165); 
assign P2_R2278_U415 = ~(P2_R2278_U209 & P2_R2278_U413); 
assign P2_R2278_U480 = ~(P2_U2801 & P2_R2278_U40); 
assign P2_R2278_U482 = ~(P2_U2801 & P2_R2278_U40); 
assign P2_R2278_U491 = ~(P2_R2278_U62 & P2_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P2_R2278_U493 = ~(P2_R2278_U62 & P2_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P2_R2278_U502 = ~(P2_R2278_U501 & P2_R2278_U500); 
assign P2_ADD_394_U90 = ~(P2_ADD_394_U184 & P2_ADD_394_U183); 
assign P2_ADD_394_U120 = ~P2_ADD_394_U52; 
assign P2_ADD_394_U149 = ~(P2_ADD_394_U52 & P2_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P2_R2267_U73 = P2_R2267_U152 & P2_R2267_U151; 
assign P2_R2267_U108 = ~P2_R2267_U37; 
assign P2_R2267_U121 = ~(P2_U2774 & P2_R2267_U120); 
assign P2_R2267_U149 = ~(P2_U2773 & P2_R2267_U37); 
assign P2_ADD_371_1212_U37 = ~P2_R2256_U19; 
assign P2_ADD_371_1212_U79 = ~(P2_ADD_371_1212_U226 & P2_ADD_371_1212_U225); 
assign P2_ADD_371_1212_U121 = P2_ADD_371_1212_U234 & P2_ADD_371_1212_U233; 
assign P2_ADD_371_1212_U144 = ~P2_ADD_371_1212_U130; 
assign P2_ADD_371_1212_U146 = ~(P2_ADD_371_1212_U145 & P2_ADD_371_1212_U130); 
assign P2_ADD_371_1212_U153 = P2_R2256_U19 | P2_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P2_ADD_371_1212_U155 = ~(P2_R2256_U19 & P2_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P2_ADD_371_1212_U237 = ~(P2_ADD_371_1212_U236 & P2_ADD_371_1212_U235); 
assign P2_ADD_371_1212_U243 = ~(P2_R2256_U19 & P2_ADD_371_1212_U38); 
assign P2_ADD_371_1212_U245 = ~(P2_R2256_U19 & P2_ADD_371_1212_U38); 
assign P2_ADD_371_1212_U263 = ~(P2_ADD_371_1212_U129 & P2_ADD_371_1212_U130); 
assign P1_R2278_U17 = P1_R2278_U272 & P1_R2278_U270; 
assign P1_R2278_U141 = P1_R2278_U286 & P1_R2278_U410; 
assign P1_R2278_U146 = P1_R2278_U401 & P1_R2278_U96; 
assign P1_R2278_U151 = P1_R2278_U286 & P1_R2278_U412; 
assign P1_R2278_U155 = P1_R2278_U394 & P1_R2278_U393 & P1_R2278_U395 & P1_R2278_U398 & P1_R2278_U156; 
assign P1_R2278_U159 = P1_R2278_U403 & P1_R2278_U187 & P1_R2278_U404; 
assign P1_R2278_U160 = P1_R2278_U286 & P1_R2278_U417; 
assign P1_R2278_U168 = P1_R2278_U286 & P1_R2278_U415; 
assign P1_R2278_U252 = ~(P1_R2278_U251 & P1_R2278_U231); 
assign P1_R2278_U266 = ~(P1_R2278_U265 & P1_R2278_U231 & P1_R2278_U179); 
assign P1_R2278_U445 = ~(P1_R2278_U443 & P1_R2278_U251); 
assign P1_R2358_U69 = ~(P1_R2358_U364 & P1_R2358_U283); 
assign P1_R2358_U74 = ~(P1_R2358_U73 & P1_R2358_U262); 
assign P1_R2358_U78 = ~(P1_R2358_U450 & P1_R2358_U449); 
assign P1_R2358_U102 = P1_R2358_U283 & P1_R2358_U282; 
assign P1_R2358_U127 = P1_R2358_U256 & P1_R2358_U353 & P1_R2358_U355 & P1_R2358_U354; 
assign P1_R2358_U140 = P1_R2358_U316 & P1_R2358_U61; 
assign P1_R2358_U173 = ~P1_U2659; 
assign P1_R2358_U198 = ~(P1_R2358_U57 & P1_R2358_U309); 
assign P1_R2358_U201 = ~(P1_R2358_U126 & P1_R2358_U199); 
assign P1_R2358_U240 = ~(P1_R2358_U122 & P1_R2358_U239); 
assign P1_R2358_U245 = ~(P1_R2358_U238 & P1_R2358_U215); 
assign P1_R2358_U284 = ~(P1_R2358_U503 & P1_R2358_U502 & P1_R2358_U43); 
assign P1_R2358_U322 = ~P1_R2358_U73; 
assign P1_R2358_U344 = ~(P1_R2358_U283 & P1_R2358_U282); 
assign P1_R2358_U512 = ~(P1_R2358_U511 & P1_R2358_U510); 
assign P1_R2358_U529 = ~(P1_U2659 & P1_R2358_U23); 
assign P1_R2358_U545 = ~(P1_U2659 & P1_R2358_U23); 
assign P1_R2358_U609 = ~(P1_R2358_U118 & P1_R2358_U269); 
assign P1_R2099_U71 = ~(P1_R2099_U309 & P1_R2099_U308); 
assign P1_R2099_U176 = ~P1_R2099_U21; 
assign P1_R2099_U307 = ~(P1_R2099_U48 & P1_R2099_U21); 
assign P1_R2337_U76 = ~(P1_R2337_U152 & P1_R2337_U151); 
assign P1_R2337_U117 = ~P1_R2337_U52; 
assign P1_R2337_U149 = ~(P1_R2337_U52 & P1_PHYADDRPOINTER_REG_26__SCAN_IN); 
assign P1_R2096_U76 = ~(P1_R2096_U152 & P1_R2096_U151); 
assign P1_R2096_U117 = ~P1_R2096_U52; 
assign P1_R2096_U149 = ~(P1_R2096_U52 & P1_REIP_REG_26__SCAN_IN); 
assign P1_ADD_405_U90 = ~(P1_ADD_405_U184 & P1_ADD_405_U183); 
assign P1_ADD_405_U120 = ~P1_ADD_405_U52; 
assign P1_ADD_405_U149 = ~(P1_ADD_405_U52 & P1_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P1_ADD_515_U90 = ~(P1_ADD_515_U180 & P1_ADD_515_U179); 
assign P1_ADD_515_U117 = ~P1_ADD_515_U52; 
assign P1_ADD_515_U147 = ~(P1_ADD_515_U52 & P1_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_U2806 = ~(P3_U6598 & P3_U6600 & P3_U6597 & P3_U6599 & P3_U3978); 
assign P3_U2841 = ~(P3_U3853 & P3_U6158); 
assign P3_U2842 = ~(P3_U3845 & P3_U6134); 
assign P3_U3867 = P3_U6185 & P3_U6186 & P3_U3864 & P3_U3866 & P3_U6184; 
assign P3_U3872 = P3_U3869 & P3_U3868 & P3_U3870 & P3_U3871; 
assign P3_U6182 = ~(P3_U4318 & P3_U6180); 
assign P3_U6210 = ~(P3_ADD_558_U80 & P3_U3220); 
assign P3_U6211 = ~(P3_ADD_553_U80 & P3_U4298); 
assign P3_U6212 = ~(P3_ADD_547_U80 & P3_U4299); 
assign P3_U6215 = ~(P3_ADD_531_U80 & P3_U2354); 
assign P3_U6223 = ~(P3_ADD_385_U80 & P3_U2358); 
assign P3_U6224 = ~(P3_ADD_380_U80 & P3_U2359); 
assign P3_U6225 = ~(P3_ADD_349_U80 & P3_U4306); 
assign P3_U6226 = ~(P3_ADD_344_U80 & P3_U2362); 
assign P3_U6232 = ~(P3_ADD_360_1242_U13 & P3_U2395); 
assign P3_U6237 = ~(P3_ADD_541_U76 & P3_U4300); 
assign P3_U6238 = ~(P3_ADD_536_U76 & P3_U4301); 
assign P3_U6241 = ~(P3_ADD_515_U76 & P3_U4302); 
assign P3_U6242 = ~(P3_ADD_494_U76 & P3_U2356); 
assign P3_U6243 = ~(P3_ADD_476_U76 & P3_U4303); 
assign P3_U6244 = ~(P3_ADD_441_U76 & P3_U4304); 
assign P3_U6245 = ~(P3_ADD_405_U75 & P3_U4305); 
assign P3_U6246 = ~(P3_ADD_394_U75 & P3_U2357); 
assign P3_U6275 = ~(P3_ADD_371_1212_U15 & P3_U2360); 
assign P3_U6377 = ~(P3_SUB_357_1258_U20 & P3_U2393); 
assign P3_U6605 = ~(P3_ADD_318_U76 & P3_U2398); 
assign P3_U6607 = ~(P3_U2396 & P3_ADD_360_1242_U13); 
assign P3_U6610 = ~(P3_ADD_339_U76 & P3_U2388); 
assign P3_U6614 = ~(P3_ADD_315_U72 & P3_U2397); 
assign P3_U6619 = ~(P3_U2387 & P3_ADD_371_1212_U15); 
assign P3_U6656 = ~(P3_U2394 & P3_SUB_357_1258_U20); 
assign P3_U7310 = ~(P3_ADD_467_U76 & P3_U2601); 
assign P3_U7312 = ~(P3_ADD_430_U76 & P3_U2405); 
assign P2_U2799 = P2_U3242 & P2_R2267_U73; 
assign P2_U2873 = ~(P2_U6514 & P2_U6515 & P2_U6513); 
assign P2_U2911 = ~(P2_U4067 & P2_U6359 & P2_U6360); 
assign P2_U3633 = ~(P2_U8320 & P2_U8319); 
assign P2_U4118 = P2_U6691 & P2_U4446 & P2_U6694; 
assign P2_U6434 = ~(P2_U2380 & P2_R2096_U83); 
assign P2_U6522 = ~(P2_R2182_U89 & P2_U2393); 
assign P2_U6755 = ~(P2_R2267_U73 & P2_U2587); 
assign P2_U6772 = ~(P2_U2588 & P2_R2096_U83); 
assign P2_U8313 = ~(P2_R2256_U5 & P2_U3572); 
assign P2_U8383 = ~(P2_R2337_U74 & P2_U3284); 
assign P1_U2658 = ~(P1_U6800 & P1_U4016); 
assign P1_U3033 = ~(P1_U5460 & P1_U5459 & P1_U3730); 
assign P1_U3034 = ~(P1_U5455 & P1_U5454 & P1_U3729); 
assign P1_U3035 = ~(P1_U5450 & P1_U5449 & P1_U3728); 
assign P1_U3036 = ~(P1_U5445 & P1_U5444 & P1_U3727); 
assign P1_U3037 = ~(P1_U7612 & P1_U5440 & P1_U3726); 
assign P1_U3038 = ~(P1_U5436 & P1_U5435 & P1_U3725); 
assign P1_U3039 = ~(P1_U5431 & P1_U5430 & P1_U3724); 
assign P1_U3040 = ~(P1_U5426 & P1_U5425 & P1_U3723); 
assign P1_U3041 = ~(P1_U5404 & P1_U5403 & P1_U3721); 
assign P1_U3042 = ~(P1_U5399 & P1_U5398 & P1_U3720); 
assign P1_U3043 = ~(P1_U5394 & P1_U5393 & P1_U3719); 
assign P1_U3044 = ~(P1_U5389 & P1_U5388 & P1_U3718); 
assign P1_U3045 = ~(P1_U5384 & P1_U5383 & P1_U3717); 
assign P1_U3046 = ~(P1_U5379 & P1_U5378 & P1_U3716); 
assign P1_U3047 = ~(P1_U5374 & P1_U5373 & P1_U3715); 
assign P1_U3048 = ~(P1_U5369 & P1_U5368 & P1_U3714); 
assign P1_U3049 = ~(P1_U5346 & P1_U5345 & P1_U3712); 
assign P1_U3050 = ~(P1_U5341 & P1_U5340 & P1_U3711); 
assign P1_U3051 = ~(P1_U5336 & P1_U5335 & P1_U3710); 
assign P1_U3052 = ~(P1_U5331 & P1_U5330 & P1_U3709); 
assign P1_U3053 = ~(P1_U5326 & P1_U5325 & P1_U3708); 
assign P1_U3054 = ~(P1_U5321 & P1_U5320 & P1_U3707); 
assign P1_U3055 = ~(P1_U5316 & P1_U5315 & P1_U3706); 
assign P1_U3056 = ~(P1_U5311 & P1_U5310 & P1_U3705); 
assign P1_U3057 = ~(P1_U5289 & P1_U5288 & P1_U3703); 
assign P1_U3058 = ~(P1_U5284 & P1_U5283 & P1_U3702); 
assign P1_U3059 = ~(P1_U5279 & P1_U5278 & P1_U3701); 
assign P1_U3060 = ~(P1_U5274 & P1_U5273 & P1_U3700); 
assign P1_U3061 = ~(P1_U5269 & P1_U5268 & P1_U3699); 
assign P1_U3062 = ~(P1_U5264 & P1_U5263 & P1_U3698); 
assign P1_U3063 = ~(P1_U5259 & P1_U5258 & P1_U3697); 
assign P1_U3064 = ~(P1_U5254 & P1_U5253 & P1_U3696); 
assign P1_U3065 = ~(P1_U5231 & P1_U5230 & P1_U3694); 
assign P1_U3066 = ~(P1_U5226 & P1_U5225 & P1_U3693); 
assign P1_U3067 = ~(P1_U5221 & P1_U5220 & P1_U3692); 
assign P1_U3068 = ~(P1_U5216 & P1_U5215 & P1_U3691); 
assign P1_U3069 = ~(P1_U5211 & P1_U5210 & P1_U3690); 
assign P1_U3070 = ~(P1_U5206 & P1_U5205 & P1_U3689); 
assign P1_U3071 = ~(P1_U5201 & P1_U5200 & P1_U3688); 
assign P1_U3072 = ~(P1_U5196 & P1_U5195 & P1_U3687); 
assign P1_U3073 = ~(P1_U5174 & P1_U5173 & P1_U3685); 
assign P1_U3074 = ~(P1_U5169 & P1_U5168 & P1_U3684); 
assign P1_U3075 = ~(P1_U5164 & P1_U5163 & P1_U3683); 
assign P1_U3076 = ~(P1_U5159 & P1_U5158 & P1_U3682); 
assign P1_U3077 = ~(P1_U5154 & P1_U5153 & P1_U3681); 
assign P1_U3078 = ~(P1_U5149 & P1_U5148 & P1_U3680); 
assign P1_U3079 = ~(P1_U5144 & P1_U5143 & P1_U3679); 
assign P1_U3080 = ~(P1_U5139 & P1_U5138 & P1_U3678); 
assign P1_U3081 = ~(P1_U5116 & P1_U5115 & P1_U3676); 
assign P1_U3082 = ~(P1_U5111 & P1_U5110 & P1_U3675); 
assign P1_U3083 = ~(P1_U5106 & P1_U5105 & P1_U3674); 
assign P1_U3084 = ~(P1_U5101 & P1_U5100 & P1_U3673); 
assign P1_U3085 = ~(P1_U5096 & P1_U5095 & P1_U3672); 
assign P1_U3086 = ~(P1_U5091 & P1_U5090 & P1_U3671); 
assign P1_U3087 = ~(P1_U5086 & P1_U5085 & P1_U3670); 
assign P1_U3088 = ~(P1_U5081 & P1_U5080 & P1_U3669); 
assign P1_U3089 = ~(P1_U5059 & P1_U5058 & P1_U3667); 
assign P1_U3090 = ~(P1_U5054 & P1_U5053 & P1_U3666); 
assign P1_U3091 = ~(P1_U5049 & P1_U5048 & P1_U3665); 
assign P1_U3092 = ~(P1_U5044 & P1_U5043 & P1_U3664); 
assign P1_U3093 = ~(P1_U5039 & P1_U5038 & P1_U3663); 
assign P1_U3094 = ~(P1_U5034 & P1_U5033 & P1_U3662); 
assign P1_U3095 = ~(P1_U5029 & P1_U5028 & P1_U3661); 
assign P1_U3096 = ~(P1_U5024 & P1_U5023 & P1_U3660); 
assign P1_U5607 = ~(P1_R2278_U17 & P1_U2377); 
assign P1_U5738 = ~(P1_R2099_U71 & P1_U2380); 
assign P1_U5748 = ~(P1_ADD_405_U90 & P1_U2375); 
assign P1_U5749 = ~(P1_ADD_515_U90 & P1_U2374); 
assign P1_U5825 = ~(P1_U2372 & P1_R2278_U17); 
assign P1_U5847 = ~(P1_R2358_U78 & P1_U2364); 
assign P1_U5924 = ~(P1_R2337_U76 & P1_U2376); 
assign P1_U6182 = ~(P1_U2386 & P1_R2358_U78); 
assign P1_U6292 = ~(P1_U2383 & P1_R2358_U78); 
assign P1_U6338 = ~(P1_U2371 & P1_R2099_U71); 
assign P1_U6542 = ~(P1_U2604 & P1_R2099_U71); 
assign P1_U6550 = ~(P1_R2096_U76 & P1_U7485); 
assign P1_U6799 = ~(P1_R2337_U76 & P1_U2352); 
assign P3_ADD_476_U54 = ~(P3_ADD_476_U117 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_476_U150 = ~(P3_ADD_476_U117 & P3_ADD_476_U53); 
assign P3_ADD_531_U55 = ~(P3_ADD_531_U121 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_531_U157 = ~(P3_ADD_531_U121 & P3_ADD_531_U54); 
assign P3_SUB_320_U13 = P3_SUB_320_U112 & P3_SUB_320_U35; 
assign P3_SUB_320_U65 = ~P3_ADD_318_U76; 
assign P3_SUB_320_U100 = ~P3_SUB_320_U35; 
assign P3_SUB_320_U142 = ~(P3_ADD_318_U76 & P3_SUB_320_U35); 
assign P3_ADD_318_U54 = ~(P3_ADD_318_U117 & P3_PHYADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_318_U150 = ~(P3_ADD_318_U117 & P3_ADD_318_U53); 
assign P3_ADD_315_U54 = ~(P3_ADD_315_U114 & P3_PHYADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_315_U142 = ~(P3_ADD_315_U114 & P3_ADD_315_U53); 
assign P3_ADD_360_1242_U14 = P3_ADD_360_1242_U169 & P3_ADD_360_1242_U68; 
assign P3_ADD_360_1242_U163 = ~P3_ADD_360_1242_U68; 
assign P3_ADD_360_1242_U238 = ~(P3_ADD_360_1242_U68 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_467_U54 = ~(P3_ADD_467_U117 & P3_REIP_REG_26__SCAN_IN); 
assign P3_ADD_467_U150 = ~(P3_ADD_467_U117 & P3_ADD_467_U53); 
assign P3_ADD_430_U54 = ~(P3_ADD_430_U117 & P3_REIP_REG_26__SCAN_IN); 
assign P3_ADD_430_U150 = ~(P3_ADD_430_U117 & P3_ADD_430_U53); 
assign P3_ADD_380_U55 = ~(P3_ADD_380_U121 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_380_U157 = ~(P3_ADD_380_U121 & P3_ADD_380_U54); 
assign P3_ADD_344_U55 = ~(P3_ADD_344_U121 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_344_U157 = ~(P3_ADD_344_U121 & P3_ADD_344_U54); 
assign P3_ADD_339_U54 = ~(P3_ADD_339_U117 & P3_PHYADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_339_U150 = ~(P3_ADD_339_U117 & P3_ADD_339_U53); 
assign P3_ADD_541_U54 = ~(P3_ADD_541_U117 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_541_U150 = ~(P3_ADD_541_U117 & P3_ADD_541_U53); 
assign P3_ADD_515_U54 = ~(P3_ADD_515_U117 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_515_U150 = ~(P3_ADD_515_U117 & P3_ADD_515_U53); 
assign P3_ADD_394_U54 = ~(P3_ADD_394_U120 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_394_U152 = ~(P3_ADD_394_U120 & P3_ADD_394_U53); 
assign P3_ADD_441_U54 = ~(P3_ADD_441_U117 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_441_U150 = ~(P3_ADD_441_U117 & P3_ADD_441_U53); 
assign P3_ADD_349_U55 = ~(P3_ADD_349_U121 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_349_U157 = ~(P3_ADD_349_U121 & P3_ADD_349_U54); 
assign P3_ADD_405_U54 = ~(P3_ADD_405_U120 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_405_U152 = ~(P3_ADD_405_U120 & P3_ADD_405_U53); 
assign P3_ADD_553_U55 = ~(P3_ADD_553_U121 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_553_U157 = ~(P3_ADD_553_U121 & P3_ADD_553_U54); 
assign P3_ADD_558_U55 = ~(P3_ADD_558_U121 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_558_U157 = ~(P3_ADD_558_U121 & P3_ADD_558_U54); 
assign P3_ADD_385_U55 = ~(P3_ADD_385_U121 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_385_U157 = ~(P3_ADD_385_U121 & P3_ADD_385_U54); 
assign P3_ADD_547_U55 = ~(P3_ADD_547_U121 & P3_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P3_ADD_547_U157 = ~(P3_ADD_547_U121 & P3_ADD_547_U54); 
assign P3_ADD_371_1212_U73 = ~(P3_ADD_371_1212_U107 & P3_ADD_371_1212_U172); 
assign P3_ADD_371_1212_U177 = ~(P3_ADD_371_1212_U172 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_371_1212_U246 = ~(P3_ADD_371_1212_U172 & P3_ADD_371_1212_U72); 
assign P3_ADD_494_U54 = ~(P3_ADD_494_U117 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_494_U150 = ~(P3_ADD_494_U117 & P3_ADD_494_U53); 
assign P3_ADD_536_U54 = ~(P3_ADD_536_U117 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_536_U150 = ~(P3_ADD_536_U117 & P3_ADD_536_U53); 
assign P2_R2099_U88 = ~(P2_R2099_U213 & P2_R2099_U212); 
assign P2_R2099_U131 = ~P2_R2099_U37; 
assign P2_R2099_U210 = ~(P2_U2731 & P2_R2099_U37); 
assign P2_ADD_391_1196_U56 = ~P2_R2182_U89; 
assign P2_ADD_391_1196_U71 = ~P2_R2096_U83; 
assign P2_ADD_391_1196_U153 = P2_ADD_391_1196_U455 & P2_ADD_391_1196_U454; 
assign P2_ADD_391_1196_U196 = ~(P2_ADD_391_1196_U194 & P2_ADD_391_1196_U195); 
assign P2_ADD_391_1196_U207 = ~P2_ADD_391_1196_U50; 
assign P2_ADD_391_1196_U232 = P2_R2182_U89 | P2_R2096_U90; 
assign P2_ADD_391_1196_U234 = ~(P2_R2096_U90 & P2_R2182_U89); 
assign P2_ADD_391_1196_U298 = ~(P2_ADD_391_1196_U297 & P2_ADD_391_1196_U50); 
assign P2_ADD_391_1196_U441 = ~(P2_R2182_U89 & P2_ADD_391_1196_U57); 
assign P2_ADD_391_1196_U443 = ~(P2_R2182_U89 & P2_ADD_391_1196_U57); 
assign P2_ADD_391_1196_U447 = ~(P2_R2096_U91 & P2_ADD_391_1196_U54); 
assign P2_ADD_391_1196_U449 = ~(P2_R2096_U91 & P2_ADD_391_1196_U54); 
assign P2_ADD_391_1196_U475 = ~(P2_ADD_391_1196_U305 & P2_ADD_391_1196_U50); 
assign P2_R2182_U11 = P2_U2692 & P2_R2182_U13; 
assign P2_R2182_U88 = ~(P2_R2182_U287 & P2_R2182_U286); 
assign P2_R2182_U151 = ~P2_R2182_U13; 
assign P2_R2182_U277 = ~(P2_R2182_U31 & P2_R2182_U13); 
assign P2_R2182_U285 = ~(P2_R2182_U150 & P2_U2693); 
assign P2_R2027_U55 = ~(P2_R2027_U121 & P2_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P2_R2027_U157 = ~(P2_R2027_U121 & P2_R2027_U54); 
assign P2_R2337_U55 = ~(P2_R2337_U118 & P2_PHYADDRPOINTER_REG_27__SCAN_IN); 
assign P2_R2337_U148 = ~(P2_R2337_U118 & P2_R2337_U54); 
assign P2_R2096_U13 = P2_U2622 & P2_R2096_U15; 
assign P2_R2096_U82 = ~(P2_R2096_U228 & P2_R2096_U227); 
assign P2_R2096_U162 = ~P2_R2096_U15; 
assign P2_R2096_U223 = ~(P2_R2096_U38 & P2_R2096_U15); 
assign P2_R2096_U226 = ~(P2_R2096_U161 & P2_U2623); 
assign P2_R2256_U18 = ~(P2_R2256_U50 & P2_R2256_U49); 
assign P2_R2256_U44 = ~P2_R2256_U24; 
assign P2_R2256_U47 = ~(P2_U3622 & P2_R2256_U24); 
assign P2_R1957_U13 = P2_R1957_U112 & P2_R1957_U34; 
assign P2_R1957_U65 = ~P2_U3665; 
assign P2_R1957_U100 = ~P2_R1957_U34; 
assign P2_R1957_U142 = ~(P2_U3665 & P2_R1957_U34); 
assign P2_R2278_U66 = ~P2_U2800; 
assign P2_R2278_U68 = ~(P2_U2800 & P2_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P2_R2278_U92 = ~(P2_R2278_U415 & P2_R2278_U414); 
assign P2_R2278_U114 = P2_R2278_U313 & P2_R2278_U215; 
assign P2_R2278_U129 = P2_R2278_U273 & P2_R2278_U270; 
assign P2_R2278_U130 = P2_R2278_U331 & P2_R2278_U273; 
assign P2_R2278_U157 = P2_R2278_U389 & P2_R2278_U388; 
assign P2_R2278_U185 = P2_R2278_U492 & P2_R2278_U491; 
assign P2_R2278_U219 = ~P2_R2278_U23; 
assign P2_R2278_U276 = P2_U2800 | P2_INSTADDRPOINTER_REG_21__SCAN_IN; 
assign P2_R2278_U312 = ~(P2_R2278_U113 & P2_R2278_U165); 
assign P2_R2278_U330 = ~(P2_R2278_U331 & P2_R2278_U332); 
assign P2_R2278_U381 = ~(P2_R2278_U21 & P2_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P2_R2278_U383 = ~(P2_R2278_U21 & P2_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P2_R2278_U392 = ~(P2_R2278_U391 & P2_R2278_U390); 
assign P2_R2278_U473 = ~(P2_U2800 & P2_R2278_U67); 
assign P2_R2278_U475 = ~(P2_U2800 & P2_R2278_U67); 
assign P2_R2278_U479 = ~(P2_R2278_U39 & P2_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P2_R2278_U481 = ~(P2_R2278_U39 & P2_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P2_R2278_U495 = ~(P2_R2278_U494 & P2_R2278_U493); 
assign P2_ADD_394_U54 = ~(P2_ADD_394_U120 & P2_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P2_ADD_394_U150 = ~(P2_ADD_394_U120 & P2_ADD_394_U53); 
assign P2_R2267_U12 = P2_R2267_U121 & P2_R2267_U37; 
assign P2_R2267_U38 = ~(P2_R2267_U52 & P2_R2267_U108); 
assign P2_R2267_U118 = ~(P2_R2267_U108 & P2_R2267_U70); 
assign P2_R2267_U150 = ~(P2_R2267_U108 & P2_R2267_U70); 
assign P2_ADD_371_1212_U41 = ~P2_R2256_U5; 
assign P2_ADD_371_1212_U122 = ~(P2_ADD_371_1212_U147 & P2_ADD_371_1212_U146); 
assign P2_ADD_371_1212_U165 = P2_R2256_U5 | P2_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P2_ADD_371_1212_U166 = ~(P2_R2256_U5 & P2_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P2_ADD_371_1212_U242 = ~(P2_ADD_371_1212_U37 & P2_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P2_ADD_371_1212_U244 = ~(P2_ADD_371_1212_U37 & P2_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P2_ADD_371_1212_U250 = ~(P2_R2256_U5 & P2_ADD_371_1212_U42); 
assign P2_ADD_371_1212_U252 = ~(P2_R2256_U5 & P2_ADD_371_1212_U42); 
assign P2_ADD_371_1212_U264 = ~(P2_ADD_371_1212_U144 & P2_ADD_371_1212_U262); 
assign P1_R2278_U41 = ~(P1_R2278_U254 & P1_R2278_U252 & P1_R2278_U253); 
assign P1_R2278_U103 = ~(P1_R2278_U445 & P1_R2278_U444); 
assign P1_R2278_U353 = ~(P1_R2278_U253 & P1_R2278_U252 & P1_R2278_U128); 
assign P1_R2358_U20 = P1_R2358_U245 & P1_R2358_U244; 
assign P1_R2358_U21 = P1_R2358_U242 & P1_R2358_U240; 
assign P1_R2358_U119 = ~(P1_R2358_U609 & P1_R2358_U608); 
assign P1_R2358_U130 = P1_R2358_U7 & P1_R2358_U284; 
assign P1_R2358_U197 = ~(P1_R2358_U201 & P1_R2358_U127); 
assign P1_R2358_U285 = ~(P1_U2628 & P1_R2358_U512); 
assign P1_R2358_U310 = ~P1_R2358_U198; 
assign P1_R2358_U311 = ~(P1_R2358_U198 & P1_R2358_U258); 
assign P1_R2358_U323 = ~P1_R2358_U74; 
assign P1_R2358_U324 = ~(P1_R2358_U74 & P1_R2358_U263); 
assign P1_R2358_U327 = ~(P1_R2358_U142 & P1_R2358_U74); 
assign P1_R2358_U329 = ~(P1_R2358_U322 & P1_R2358_U328); 
assign P1_R2358_U365 = ~P1_R2358_U69; 
assign P1_R2358_U366 = ~(P1_R2358_U69 & P1_R2358_U284); 
assign P1_R2358_U528 = ~(P1_U2352 & P1_R2358_U173); 
assign P1_R2358_U544 = ~(P1_U2352 & P1_R2358_U173); 
assign P1_R2358_U606 = ~(P1_R2358_U351 & P1_R2358_U198); 
assign P1_R2099_U22 = ~(P1_R2099_U176 & P1_R2099_U48); 
assign P1_R2099_U306 = ~(P1_R2099_U237 & P1_R2099_U176); 
assign P1_R2337_U54 = ~(P1_R2337_U117 & P1_PHYADDRPOINTER_REG_26__SCAN_IN); 
assign P1_R2337_U150 = ~(P1_R2337_U117 & P1_R2337_U53); 
assign P1_R2096_U54 = ~(P1_R2096_U117 & P1_REIP_REG_26__SCAN_IN); 
assign P1_R2096_U150 = ~(P1_R2096_U117 & P1_R2096_U53); 
assign P1_ADD_405_U54 = ~(P1_ADD_405_U120 & P1_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P1_ADD_405_U150 = ~(P1_ADD_405_U120 & P1_ADD_405_U53); 
assign P1_ADD_515_U54 = ~(P1_ADD_515_U117 & P1_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P1_ADD_515_U148 = ~(P1_ADD_515_U117 & P1_ADD_515_U53); 
assign P3_U2840 = ~(P3_U3863 & P3_U6182); 
assign P3_U3874 = P3_U6212 & P3_U6211; 
assign P3_U3876 = P3_U6214 & P3_U6213 & P3_U6215 & P3_U3875; 
assign P3_U3880 = P3_U6224 & P3_U6223 & P3_U6225; 
assign P3_U3881 = P3_U6227 & P3_U6226; 
assign P3_U3885 = P3_U6241 & P3_U6240; 
assign P3_U3888 = P3_U6243 & P3_U6242 & P3_U6244; 
assign P3_U3889 = P3_U6246 & P3_U6245; 
assign P3_U3979 = P3_U6612 & P3_U6609 & P3_U6610 & P3_U6611; 
assign P3_U4114 = P3_U7310 & P3_U7309; 
assign P3_U6204 = ~(P3_U3872 & P3_U3867); 
assign P3_U6256 = ~(P3_ADD_360_1242_U14 & P3_U2395); 
assign P3_U6615 = ~(P3_U2396 & P3_ADD_360_1242_U14); 
assign P2_U2798 = P2_U3242 & P2_R2267_U12; 
assign P2_U3630 = ~(P2_U8314 & P2_U8313); 
assign P2_U3664 = ~(P2_U8384 & P2_U8383); 
assign P2_U6439 = ~(P2_U2380 & P2_R2096_U82); 
assign P2_U6517 = ~(P2_U2379 & P2_R2099_U88); 
assign P2_U6525 = ~(P2_R2182_U88 & P2_U2393); 
assign P2_U6702 = ~(P2_U2392 & P2_R2099_U88); 
assign P2_U6763 = ~(P2_R2267_U12 & P2_U2587); 
assign P2_U6780 = ~(P2_U2588 & P2_R2096_U82); 
assign P2_U8317 = ~(P2_R2256_U18 & P2_U3572); 
assign P1_U2863 = ~(P1_U6293 & P1_U6294 & P1_U6292); 
assign P1_U2895 = ~(P1_U6183 & P1_U6181 & P1_U6182); 
assign P1_U2994 = ~(P1_U5826 & P1_U5824 & P1_U5825 & P1_U5828 & P1_U5827); 
assign P1_U3026 = ~(P1_U3781 & P1_U3783 & P1_U5607); 
assign P1_U3841 = P1_U5746 & P1_U5748; 
assign P1_U3843 = P1_U3842 & P1_U5749; 
assign P1_U3936 = P1_U6552 & P1_U6550; 
assign P1_U4015 = P1_U6797 & P1_U6798 & P1_U6799; 
assign P1_U5614 = ~(P1_R2278_U103 & P1_U2377); 
assign P1_U5830 = ~(P1_U2372 & P1_R2278_U103); 
assign P1_U5832 = ~(P1_R2358_U20 & P1_U2364); 
assign P1_U5837 = ~(P1_R2358_U21 & P1_U2364); 
assign P1_U5862 = ~(P1_R2358_U119 & P1_U2364); 
assign P1_U6173 = ~(P1_U2386 & P1_R2358_U20); 
assign P1_U6176 = ~(P1_U2386 & P1_R2358_U21); 
assign P1_U6191 = ~(P1_U2386 & P1_R2358_U119); 
assign P1_U6283 = ~(P1_U2383 & P1_R2358_U20); 
assign P1_U6286 = ~(P1_U2383 & P1_R2358_U21); 
assign P1_U6301 = ~(P1_U2383 & P1_R2358_U119); 
assign P3_ADD_476_U75 = ~(P3_ADD_476_U150 & P3_ADD_476_U149); 
assign P3_ADD_476_U118 = ~P3_ADD_476_U54; 
assign P3_ADD_476_U147 = ~(P3_ADD_476_U54 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_531_U79 = ~(P3_ADD_531_U157 & P3_ADD_531_U156); 
assign P3_ADD_531_U122 = ~P3_ADD_531_U55; 
assign P3_ADD_531_U154 = ~(P3_ADD_531_U55 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_SUB_320_U109 = ~(P3_SUB_320_U100 & P3_SUB_320_U65); 
assign P3_SUB_320_U143 = ~(P3_SUB_320_U100 & P3_SUB_320_U65); 
assign P3_ADD_318_U75 = ~(P3_ADD_318_U150 & P3_ADD_318_U149); 
assign P3_ADD_318_U118 = ~P3_ADD_318_U54; 
assign P3_ADD_318_U147 = ~(P3_ADD_318_U54 & P3_PHYADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_315_U71 = ~(P3_ADD_315_U142 & P3_ADD_315_U141); 
assign P3_ADD_315_U115 = ~P3_ADD_315_U54; 
assign P3_ADD_315_U139 = ~(P3_ADD_315_U54 & P3_PHYADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_360_1242_U71 = ~(P3_ADD_360_1242_U104 & P3_ADD_360_1242_U163); 
assign P3_ADD_360_1242_U167 = ~(P3_ADD_360_1242_U163 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_360_1242_U239 = ~(P3_ADD_360_1242_U163 & P3_ADD_360_1242_U70); 
assign P3_ADD_467_U75 = ~(P3_ADD_467_U150 & P3_ADD_467_U149); 
assign P3_ADD_467_U118 = ~P3_ADD_467_U54; 
assign P3_ADD_467_U147 = ~(P3_ADD_467_U54 & P3_REIP_REG_27__SCAN_IN); 
assign P3_ADD_430_U75 = ~(P3_ADD_430_U150 & P3_ADD_430_U149); 
assign P3_ADD_430_U118 = ~P3_ADD_430_U54; 
assign P3_ADD_430_U147 = ~(P3_ADD_430_U54 & P3_REIP_REG_27__SCAN_IN); 
assign P3_ADD_380_U79 = ~(P3_ADD_380_U157 & P3_ADD_380_U156); 
assign P3_ADD_380_U122 = ~P3_ADD_380_U55; 
assign P3_ADD_380_U154 = ~(P3_ADD_380_U55 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_344_U79 = ~(P3_ADD_344_U157 & P3_ADD_344_U156); 
assign P3_ADD_344_U122 = ~P3_ADD_344_U55; 
assign P3_ADD_344_U154 = ~(P3_ADD_344_U55 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_339_U75 = ~(P3_ADD_339_U150 & P3_ADD_339_U149); 
assign P3_ADD_339_U118 = ~P3_ADD_339_U54; 
assign P3_ADD_339_U147 = ~(P3_ADD_339_U54 & P3_PHYADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_541_U75 = ~(P3_ADD_541_U150 & P3_ADD_541_U149); 
assign P3_ADD_541_U118 = ~P3_ADD_541_U54; 
assign P3_ADD_541_U147 = ~(P3_ADD_541_U54 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_515_U75 = ~(P3_ADD_515_U150 & P3_ADD_515_U149); 
assign P3_ADD_515_U118 = ~P3_ADD_515_U54; 
assign P3_ADD_515_U147 = ~(P3_ADD_515_U54 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_394_U74 = ~(P3_ADD_394_U152 & P3_ADD_394_U151); 
assign P3_ADD_394_U121 = ~P3_ADD_394_U54; 
assign P3_ADD_394_U149 = ~(P3_ADD_394_U54 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_441_U75 = ~(P3_ADD_441_U150 & P3_ADD_441_U149); 
assign P3_ADD_441_U118 = ~P3_ADD_441_U54; 
assign P3_ADD_441_U147 = ~(P3_ADD_441_U54 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_349_U79 = ~(P3_ADD_349_U157 & P3_ADD_349_U156); 
assign P3_ADD_349_U122 = ~P3_ADD_349_U55; 
assign P3_ADD_349_U154 = ~(P3_ADD_349_U55 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_405_U74 = ~(P3_ADD_405_U152 & P3_ADD_405_U151); 
assign P3_ADD_405_U121 = ~P3_ADD_405_U54; 
assign P3_ADD_405_U149 = ~(P3_ADD_405_U54 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_553_U79 = ~(P3_ADD_553_U157 & P3_ADD_553_U156); 
assign P3_ADD_553_U122 = ~P3_ADD_553_U55; 
assign P3_ADD_553_U154 = ~(P3_ADD_553_U55 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_558_U79 = ~(P3_ADD_558_U157 & P3_ADD_558_U156); 
assign P3_ADD_558_U122 = ~P3_ADD_558_U55; 
assign P3_ADD_558_U154 = ~(P3_ADD_558_U55 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_385_U79 = ~(P3_ADD_385_U157 & P3_ADD_385_U156); 
assign P3_ADD_385_U122 = ~P3_ADD_385_U55; 
assign P3_ADD_385_U154 = ~(P3_ADD_385_U55 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_547_U79 = ~(P3_ADD_547_U157 & P3_ADD_547_U156); 
assign P3_ADD_547_U122 = ~P3_ADD_547_U55; 
assign P3_ADD_547_U154 = ~(P3_ADD_547_U55 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_371_1212_U80 = ~(P3_ADD_371_1212_U246 & P3_ADD_371_1212_U245); 
assign P3_ADD_371_1212_U173 = ~P3_ADD_371_1212_U73; 
assign P3_ADD_371_1212_U176 = ~(P3_ADD_371_1212_U74 & P3_ADD_371_1212_U73); 
assign P3_ADD_371_1212_U178 = ~(P3_ADD_371_1212_U71 & P3_ADD_371_1212_U177); 
assign P3_ADD_494_U75 = ~(P3_ADD_494_U150 & P3_ADD_494_U149); 
assign P3_ADD_494_U118 = ~P3_ADD_494_U54; 
assign P3_ADD_494_U147 = ~(P3_ADD_494_U54 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_536_U75 = ~(P3_ADD_536_U150 & P3_ADD_536_U149); 
assign P3_ADD_536_U118 = ~P3_ADD_536_U54; 
assign P3_ADD_536_U147 = ~(P3_ADD_536_U54 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P2_R2099_U39 = ~(P2_U2731 & P2_R2099_U131); 
assign P2_R2099_U211 = ~(P2_R2099_U131 & P2_R2099_U38); 
assign P2_ADD_391_1196_U11 = P2_ADD_391_1196_U196 & P2_ADD_391_1196_U192; 
assign P2_ADD_391_1196_U58 = ~P2_R2182_U88; 
assign P2_ADD_391_1196_U73 = ~P2_R2096_U82; 
assign P2_ADD_391_1196_U151 = P2_ADD_391_1196_U448 & P2_ADD_391_1196_U447; 
assign P2_ADD_391_1196_U208 = ~(P2_ADD_391_1196_U207 & P2_ADD_391_1196_U158); 
assign P2_ADD_391_1196_U236 = P2_R2182_U88 | P2_R2096_U89; 
assign P2_ADD_391_1196_U238 = ~(P2_R2096_U89 & P2_R2182_U88); 
assign P2_ADD_391_1196_U299 = ~(P2_ADD_391_1196_U298 & P2_ADD_391_1196_U158 & P2_ADD_391_1196_U157); 
assign P2_ADD_391_1196_U434 = ~(P2_R2182_U88 & P2_ADD_391_1196_U59); 
assign P2_ADD_391_1196_U436 = ~(P2_R2182_U88 & P2_ADD_391_1196_U59); 
assign P2_ADD_391_1196_U440 = ~(P2_R2096_U90 & P2_ADD_391_1196_U56); 
assign P2_ADD_391_1196_U442 = ~(P2_R2096_U90 & P2_ADD_391_1196_U56); 
assign P2_ADD_391_1196_U451 = ~(P2_ADD_391_1196_U450 & P2_ADD_391_1196_U449); 
assign P2_ADD_391_1196_U476 = ~(P2_ADD_391_1196_U474 & P2_ADD_391_1196_U207); 
assign P2_R2182_U8 = P2_U2691 & P2_R2182_U11; 
assign P2_R2182_U87 = ~(P2_R2182_U285 & P2_R2182_U284); 
assign P2_R2182_U152 = ~P2_R2182_U11; 
assign P2_R2182_U275 = ~(P2_R2182_U32 & P2_R2182_U11); 
assign P2_R2182_U278 = ~(P2_R2182_U151 & P2_U2692); 
assign P2_R2027_U79 = ~(P2_R2027_U157 & P2_R2027_U156); 
assign P2_R2027_U122 = ~P2_R2027_U55; 
assign P2_R2027_U154 = ~(P2_R2027_U55 & P2_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P2_R2337_U73 = ~(P2_R2337_U148 & P2_R2337_U147); 
assign P2_R2337_U119 = ~P2_R2337_U55; 
assign P2_R2337_U145 = ~(P2_R2337_U55 & P2_PHYADDRPOINTER_REG_28__SCAN_IN); 
assign P2_R2096_U14 = P2_U2621 & P2_R2096_U13; 
assign P2_R2096_U81 = ~(P2_R2096_U226 & P2_R2096_U225); 
assign P2_R2096_U163 = ~P2_R2096_U13; 
assign P2_R2096_U221 = ~(P2_R2096_U41 & P2_R2096_U13); 
assign P2_R2096_U224 = ~(P2_R2096_U162 & P2_U2622); 
assign P2_R2256_U48 = ~(P2_R2256_U44 & P2_R2256_U15); 
assign P2_R1957_U109 = ~(P2_R1957_U100 & P2_R1957_U65); 
assign P2_R1957_U143 = ~(P2_R1957_U100 & P2_R1957_U65); 
assign P2_R2278_U9 = ~P2_U3633; 
assign P2_R2278_U37 = ~P2_U2799; 
assign P2_R2278_U155 = P2_R2278_U382 & P2_R2278_U381; 
assign P2_R2278_U156 = ~(P2_R2278_U114 & P2_R2278_U312); 
assign P2_R2278_U183 = P2_R2278_U480 & P2_R2278_U479; 
assign P2_R2278_U221 = P2_U3633 | P2_INSTADDRPOINTER_REG_5__SCAN_IN; 
assign P2_R2278_U222 = ~(P2_U3633 & P2_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P2_R2278_U278 = ~P2_R2278_U68; 
assign P2_R2278_U280 = P2_U2799 | P2_INSTADDRPOINTER_REG_22__SCAN_IN; 
assign P2_R2278_U281 = ~(P2_U2799 & P2_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P2_R2278_U334 = ~(P2_R2278_U130 & P2_R2278_U332); 
assign P2_R2278_U375 = ~(P2_U3633 & P2_R2278_U10); 
assign P2_R2278_U377 = ~(P2_U3633 & P2_R2278_U10); 
assign P2_R2278_U385 = ~(P2_R2278_U384 & P2_R2278_U383); 
assign P2_R2278_U393 = ~(P2_R2278_U157 & P2_R2278_U158); 
assign P2_R2278_U394 = ~(P2_R2278_U213 & P2_R2278_U392); 
assign P2_R2278_U466 = ~(P2_U2799 & P2_R2278_U38); 
assign P2_R2278_U468 = ~(P2_U2799 & P2_R2278_U38); 
assign P2_R2278_U472 = ~(P2_R2278_U66 & P2_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P2_R2278_U474 = ~(P2_R2278_U66 & P2_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P2_R2278_U483 = ~(P2_R2278_U482 & P2_R2278_U481); 
assign P2_ADD_394_U74 = ~(P2_ADD_394_U150 & P2_ADD_394_U149); 
assign P2_ADD_394_U121 = ~P2_ADD_394_U54; 
assign P2_ADD_394_U155 = ~(P2_ADD_394_U54 & P2_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P2_R2267_U71 = P2_R2267_U150 & P2_R2267_U149; 
assign P2_R2267_U109 = ~P2_R2267_U38; 
assign P2_R2267_U119 = ~(P2_U2772 & P2_R2267_U118); 
assign P2_R2267_U147 = ~(P2_U2771 & P2_R2267_U38); 
assign P2_ADD_371_1212_U40 = ~P2_R2256_U18; 
assign P2_ADD_371_1212_U84 = ~(P2_ADD_371_1212_U264 & P2_ADD_371_1212_U263); 
assign P2_ADD_371_1212_U124 = P2_ADD_371_1212_U243 & P2_ADD_371_1212_U242; 
assign P2_ADD_371_1212_U148 = ~P2_ADD_371_1212_U122; 
assign P2_ADD_371_1212_U150 = ~(P2_ADD_371_1212_U149 & P2_ADD_371_1212_U122); 
assign P2_ADD_371_1212_U157 = P2_R2256_U18 | P2_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P2_ADD_371_1212_U159 = ~(P2_R2256_U18 & P2_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P2_ADD_371_1212_U208 = ~(P2_R2256_U18 & P2_ADD_371_1212_U39); 
assign P2_ADD_371_1212_U210 = ~(P2_R2256_U18 & P2_ADD_371_1212_U39); 
assign P2_ADD_371_1212_U238 = ~(P2_ADD_371_1212_U121 & P2_ADD_371_1212_U122); 
assign P2_ADD_371_1212_U246 = ~(P2_ADD_371_1212_U245 & P2_ADD_371_1212_U244); 
assign P2_ADD_371_1212_U249 = ~(P2_ADD_371_1212_U41 & P2_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P2_ADD_371_1212_U251 = ~(P2_ADD_371_1212_U41 & P2_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P1_R2278_U176 = ~(P1_R2278_U129 & P1_R2278_U353); 
assign P1_R2278_U178 = ~(P1_R2278_U41 & P1_R2278_U256); 
assign P1_R2278_U255 = ~P1_R2278_U41; 
assign P1_R2278_U354 = ~(P1_R2278_U353 & P1_R2278_U352 & P1_R2278_U137); 
assign P1_R2358_U71 = ~(P1_R2358_U59 & P1_R2358_U311); 
assign P1_R2358_U100 = P1_R2358_U285 & P1_R2358_U284; 
assign P1_R2358_U131 = P1_R2358_U366 & P1_R2358_U285; 
assign P1_R2358_U174 = ~P1_U2658; 
assign P1_R2358_U271 = ~P1_R2358_U197; 
assign P1_R2358_U286 = ~(P1_R2358_U529 & P1_R2358_U528 & P1_R2358_U41); 
assign P1_R2358_U325 = ~(P1_R2358_U141 & P1_R2358_U324); 
assign P1_R2358_U330 = ~(P1_R2358_U323 & P1_R2358_U263); 
assign P1_R2358_U343 = ~(P1_R2358_U285 & P1_R2358_U284); 
assign P1_R2358_U393 = ~(P1_R2358_U128 & P1_R2358_U197); 
assign P1_R2358_U395 = ~(P1_R2358_U5 & P1_R2358_U197); 
assign P1_R2358_U397 = ~(P1_R2358_U272 & P1_R2358_U197); 
assign P1_R2358_U531 = ~(P1_U2658 & P1_R2358_U23); 
assign P1_R2358_U542 = ~(P1_U2658 & P1_R2358_U23); 
assign P1_R2358_U546 = ~(P1_R2358_U545 & P1_R2358_U544); 
assign P1_R2358_U604 = ~(P1_R2358_U350 & P1_R2358_U197); 
assign P1_R2358_U607 = ~(P1_R2358_U116 & P1_R2358_U310); 
assign P1_R2099_U70 = ~(P1_R2099_U307 & P1_R2099_U306); 
assign P1_R2099_U177 = ~P1_R2099_U22; 
assign P1_R2099_U305 = ~(P1_R2099_U47 & P1_R2099_U22); 
assign P1_R2337_U75 = ~(P1_R2337_U150 & P1_R2337_U149); 
assign P1_R2337_U118 = ~P1_R2337_U54; 
assign P1_R2337_U147 = ~(P1_R2337_U54 & P1_PHYADDRPOINTER_REG_27__SCAN_IN); 
assign P1_R2096_U75 = ~(P1_R2096_U150 & P1_R2096_U149); 
assign P1_R2096_U118 = ~P1_R2096_U54; 
assign P1_R2096_U147 = ~(P1_R2096_U54 & P1_REIP_REG_27__SCAN_IN); 
assign P1_ADD_405_U74 = ~(P1_ADD_405_U150 & P1_ADD_405_U149); 
assign P1_ADD_405_U121 = ~P1_ADD_405_U54; 
assign P1_ADD_405_U155 = ~(P1_ADD_405_U54 & P1_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P1_ADD_515_U74 = ~(P1_ADD_515_U148 & P1_ADD_515_U147); 
assign P1_ADD_515_U118 = ~P1_ADD_515_U54; 
assign P1_ADD_515_U153 = ~(P1_ADD_515_U54 & P1_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_U2805 = ~(P3_U6606 & P3_U6608 & P3_U6605 & P3_U6607 & P3_U3979); 
assign P3_U3877 = P3_U6209 & P3_U6210 & P3_U3874 & P3_U6208 & P3_U3876; 
assign P3_U3882 = P3_U3879 & P3_U3878 & P3_U3881 & P3_U3880; 
assign P3_U3894 = P3_U6257 & P3_U6256; 
assign P3_U6206 = ~(P3_U4318 & P3_U6204); 
assign P3_U6234 = ~(P3_ADD_558_U79 & P3_U3220); 
assign P3_U6235 = ~(P3_ADD_553_U79 & P3_U4298); 
assign P3_U6236 = ~(P3_ADD_547_U79 & P3_U4299); 
assign P3_U6239 = ~(P3_ADD_531_U79 & P3_U2354); 
assign P3_U6247 = ~(P3_ADD_385_U79 & P3_U2358); 
assign P3_U6248 = ~(P3_ADD_380_U79 & P3_U2359); 
assign P3_U6249 = ~(P3_ADD_349_U79 & P3_U4306); 
assign P3_U6250 = ~(P3_ADD_344_U79 & P3_U2362); 
assign P3_U6261 = ~(P3_ADD_541_U75 & P3_U4300); 
assign P3_U6262 = ~(P3_ADD_536_U75 & P3_U4301); 
assign P3_U6265 = ~(P3_ADD_515_U75 & P3_U4302); 
assign P3_U6266 = ~(P3_ADD_494_U75 & P3_U2356); 
assign P3_U6267 = ~(P3_ADD_476_U75 & P3_U4303); 
assign P3_U6268 = ~(P3_ADD_441_U75 & P3_U4304); 
assign P3_U6269 = ~(P3_ADD_405_U74 & P3_U4305); 
assign P3_U6270 = ~(P3_ADD_394_U74 & P3_U2357); 
assign P3_U6299 = ~(P3_ADD_371_1212_U80 & P3_U2360); 
assign P3_U6613 = ~(P3_ADD_318_U75 & P3_U2398); 
assign P3_U6618 = ~(P3_ADD_339_U75 & P3_U2388); 
assign P3_U6622 = ~(P3_ADD_315_U71 & P3_U2397); 
assign P3_U6627 = ~(P3_U2387 & P3_ADD_371_1212_U80); 
assign P3_U7318 = ~(P3_ADD_467_U75 & P3_U2601); 
assign P3_U7320 = ~(P3_ADD_430_U75 & P3_U2405); 
assign P2_U2797 = P2_U3242 & P2_R2267_U71; 
assign P2_U2872 = ~(P2_U6517 & P2_U6518 & P2_U6516); 
assign P2_U3632 = ~(P2_U8318 & P2_U8317); 
assign P2_U6364 = ~(P2_ADD_391_1196_U11 & P2_U2397); 
assign P2_U6444 = ~(P2_U2380 & P2_R2096_U81); 
assign P2_U6528 = ~(P2_R2182_U87 & P2_U2393); 
assign P2_U6771 = ~(P2_R2267_U71 & P2_U2587); 
assign P2_U6788 = ~(P2_U2588 & P2_R2096_U81); 
assign P2_U8381 = ~(P2_R2337_U73 & P2_U3284); 
assign P1_U2657 = ~(P1_U6796 & P1_U4015); 
assign P1_U2860 = ~(P1_U6302 & P1_U6303 & P1_U6301); 
assign P1_U2865 = ~(P1_U6287 & P1_U6288 & P1_U6286); 
assign P1_U2866 = ~(P1_U6284 & P1_U6285 & P1_U6283); 
assign P1_U2892 = ~(P1_U6192 & P1_U6190 & P1_U6191); 
assign P1_U2897 = ~(P1_U6177 & P1_U6175 & P1_U6176); 
assign P1_U2898 = ~(P1_U6174 & P1_U6172 & P1_U6173); 
assign P1_U2993 = ~(P1_U5831 & P1_U5829 & P1_U5830 & P1_U5833 & P1_U5832); 
assign P1_U3025 = ~(P1_U3784 & P1_U3786 & P1_U5614); 
assign P1_U5745 = ~(P1_R2099_U70 & P1_U2380); 
assign P1_U5755 = ~(P1_ADD_405_U74 & P1_U2375); 
assign P1_U5756 = ~(P1_ADD_515_U74 & P1_U2374); 
assign P1_U5929 = ~(P1_R2337_U75 & P1_U2376); 
assign P1_U6341 = ~(P1_U2371 & P1_R2099_U70); 
assign P1_U6549 = ~(P1_U2604 & P1_R2099_U70); 
assign P1_U6557 = ~(P1_R2096_U75 & P1_U7485); 
assign P1_U6795 = ~(P1_R2337_U75 & P1_U2352); 
assign P3_ADD_476_U56 = ~(P3_ADD_476_U118 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_476_U148 = ~(P3_ADD_476_U118 & P3_ADD_476_U55); 
assign P3_ADD_531_U57 = ~(P3_ADD_531_U122 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_531_U155 = ~(P3_ADD_531_U122 & P3_ADD_531_U56); 
assign P3_SUB_320_U41 = ~P3_ADD_318_U75; 
assign P3_SUB_320_U66 = P3_SUB_320_U143 & P3_SUB_320_U142; 
assign P3_SUB_320_U110 = ~(P3_ADD_318_U75 & P3_SUB_320_U109); 
assign P3_ADD_318_U56 = ~(P3_ADD_318_U118 & P3_PHYADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_318_U148 = ~(P3_ADD_318_U118 & P3_ADD_318_U55); 
assign P3_ADD_315_U56 = ~(P3_ADD_315_U115 & P3_PHYADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_315_U140 = ~(P3_ADD_315_U115 & P3_ADD_315_U55); 
assign P3_ADD_360_1242_U78 = ~(P3_ADD_360_1242_U239 & P3_ADD_360_1242_U238); 
assign P3_ADD_360_1242_U164 = ~P3_ADD_360_1242_U71; 
assign P3_ADD_360_1242_U166 = ~(P3_ADD_360_1242_U72 & P3_ADD_360_1242_U71); 
assign P3_ADD_360_1242_U168 = ~(P3_ADD_360_1242_U69 & P3_ADD_360_1242_U167); 
assign P3_ADD_467_U56 = ~(P3_ADD_467_U118 & P3_REIP_REG_27__SCAN_IN); 
assign P3_ADD_467_U148 = ~(P3_ADD_467_U118 & P3_ADD_467_U55); 
assign P3_ADD_430_U56 = ~(P3_ADD_430_U118 & P3_REIP_REG_27__SCAN_IN); 
assign P3_ADD_430_U148 = ~(P3_ADD_430_U118 & P3_ADD_430_U55); 
assign P3_ADD_380_U57 = ~(P3_ADD_380_U122 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_380_U155 = ~(P3_ADD_380_U122 & P3_ADD_380_U56); 
assign P3_ADD_344_U57 = ~(P3_ADD_344_U122 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_344_U155 = ~(P3_ADD_344_U122 & P3_ADD_344_U56); 
assign P3_ADD_339_U56 = ~(P3_ADD_339_U118 & P3_PHYADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_339_U148 = ~(P3_ADD_339_U118 & P3_ADD_339_U55); 
assign P3_ADD_541_U56 = ~(P3_ADD_541_U118 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_541_U148 = ~(P3_ADD_541_U118 & P3_ADD_541_U55); 
assign P3_ADD_515_U56 = ~(P3_ADD_515_U118 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_515_U148 = ~(P3_ADD_515_U118 & P3_ADD_515_U55); 
assign P3_ADD_394_U56 = ~(P3_ADD_394_U121 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_394_U150 = ~(P3_ADD_394_U121 & P3_ADD_394_U55); 
assign P3_ADD_441_U56 = ~(P3_ADD_441_U118 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_441_U148 = ~(P3_ADD_441_U118 & P3_ADD_441_U55); 
assign P3_ADD_349_U57 = ~(P3_ADD_349_U122 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_349_U155 = ~(P3_ADD_349_U122 & P3_ADD_349_U56); 
assign P3_ADD_405_U56 = ~(P3_ADD_405_U121 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_405_U150 = ~(P3_ADD_405_U121 & P3_ADD_405_U55); 
assign P3_ADD_553_U57 = ~(P3_ADD_553_U122 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_553_U155 = ~(P3_ADD_553_U122 & P3_ADD_553_U56); 
assign P3_ADD_558_U57 = ~(P3_ADD_558_U122 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_558_U155 = ~(P3_ADD_558_U122 & P3_ADD_558_U56); 
assign P3_ADD_385_U57 = ~(P3_ADD_385_U122 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_385_U155 = ~(P3_ADD_385_U122 & P3_ADD_385_U56); 
assign P3_ADD_547_U57 = ~(P3_ADD_547_U122 & P3_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P3_ADD_547_U155 = ~(P3_ADD_547_U122 & P3_ADD_547_U56); 
assign P3_ADD_371_1212_U16 = P3_ADD_371_1212_U178 & P3_ADD_371_1212_U73; 
assign P3_ADD_371_1212_U75 = ~(P3_ADD_371_1212_U173 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_494_U56 = ~(P3_ADD_494_U118 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_494_U148 = ~(P3_ADD_494_U118 & P3_ADD_494_U55); 
assign P3_ADD_536_U56 = ~(P3_ADD_536_U118 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_536_U148 = ~(P3_ADD_536_U118 & P3_ADD_536_U55); 
assign P2_R2099_U87 = ~(P2_R2099_U211 & P2_R2099_U210); 
assign P2_R2099_U132 = ~P2_R2099_U39; 
assign P2_R2099_U208 = ~(P2_U2730 & P2_R2099_U39); 
assign P2_ADD_391_1196_U60 = ~P2_R2182_U87; 
assign P2_ADD_391_1196_U75 = ~P2_R2096_U81; 
assign P2_ADD_391_1196_U86 = ~(P2_ADD_391_1196_U210 & P2_ADD_391_1196_U208 & P2_ADD_391_1196_U209); 
assign P2_ADD_391_1196_U109 = ~(P2_ADD_391_1196_U476 & P2_ADD_391_1196_U475); 
assign P2_ADD_391_1196_U149 = P2_ADD_391_1196_U441 & P2_ADD_391_1196_U440; 
assign P2_ADD_391_1196_U240 = P2_R2182_U87 | P2_R2096_U88; 
assign P2_ADD_391_1196_U242 = ~(P2_R2096_U88 & P2_R2182_U87); 
assign P2_ADD_391_1196_U427 = ~(P2_R2182_U87 & P2_ADD_391_1196_U61); 
assign P2_ADD_391_1196_U429 = ~(P2_R2182_U87 & P2_ADD_391_1196_U61); 
assign P2_ADD_391_1196_U433 = ~(P2_R2096_U89 & P2_ADD_391_1196_U58); 
assign P2_ADD_391_1196_U435 = ~(P2_R2096_U89 & P2_ADD_391_1196_U58); 
assign P2_ADD_391_1196_U444 = ~(P2_ADD_391_1196_U443 & P2_ADD_391_1196_U442); 
assign P2_R2182_U7 = P2_U2690 & P2_R2182_U8; 
assign P2_R2182_U86 = ~(P2_R2182_U278 & P2_R2182_U277); 
assign P2_R2182_U153 = ~P2_R2182_U8; 
assign P2_R2182_U273 = ~(P2_R2182_U37 & P2_R2182_U8); 
assign P2_R2182_U276 = ~(P2_R2182_U152 & P2_U2691); 
assign P2_R2027_U57 = ~(P2_R2027_U122 & P2_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P2_R2027_U155 = ~(P2_R2027_U122 & P2_R2027_U56); 
assign P2_R2337_U57 = ~(P2_R2337_U119 & P2_PHYADDRPOINTER_REG_28__SCAN_IN); 
assign P2_R2337_U146 = ~(P2_R2337_U119 & P2_R2337_U56); 
assign P2_R2096_U22 = P2_U2620 & P2_R2096_U14; 
assign P2_R2096_U80 = ~(P2_R2096_U224 & P2_R2096_U223); 
assign P2_R2096_U164 = ~P2_R2096_U14; 
assign P2_R2096_U219 = ~(P2_R2096_U40 & P2_R2096_U14); 
assign P2_R2096_U222 = ~(P2_R2096_U163 & P2_U2621); 
assign P2_R2256_U17 = ~(P2_R2256_U48 & P2_R2256_U47); 
assign P2_R1957_U40 = ~P2_U3664; 
assign P2_R1957_U66 = P2_R1957_U143 & P2_R1957_U142; 
assign P2_R1957_U110 = ~(P2_U3664 & P2_R1957_U109); 
assign P2_R2278_U27 = ~P2_U3630; 
assign P2_R2278_U49 = ~(P2_U3630 & P2_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P2_R2278_U69 = ~P2_U2798; 
assign P2_R2278_U71 = ~(P2_U2798 & P2_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P2_R2278_U90 = ~(P2_R2278_U394 & P2_R2278_U393); 
assign P2_R2278_U115 = P2_R2278_U217 & P2_R2278_U221; 
assign P2_R2278_U131 = P2_R2278_U334 & P2_R2278_U274; 
assign P2_R2278_U132 = P2_R2278_U276 & P2_R2278_U280; 
assign P2_R2278_U181 = P2_R2278_U473 & P2_R2278_U472; 
assign P2_R2278_U216 = ~P2_R2278_U156; 
assign P2_R2278_U218 = ~(P2_R2278_U217 & P2_R2278_U156); 
assign P2_R2278_U231 = P2_U3630 | P2_INSTADDRPOINTER_REG_8__SCAN_IN; 
assign P2_R2278_U283 = P2_U2798 | P2_INSTADDRPOINTER_REG_23__SCAN_IN; 
assign P2_R2278_U316 = ~(P2_R2278_U219 & P2_R2278_U221); 
assign P2_R2278_U336 = ~(P2_R2278_U278 & P2_R2278_U280); 
assign P2_R2278_U354 = ~(P2_U3630 & P2_R2278_U28); 
assign P2_R2278_U356 = ~(P2_U3630 & P2_R2278_U28); 
assign P2_R2278_U374 = ~(P2_R2278_U9 & P2_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P2_R2278_U376 = ~(P2_R2278_U9 & P2_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P2_R2278_U386 = ~(P2_R2278_U155 & P2_R2278_U156); 
assign P2_R2278_U459 = ~(P2_U2798 & P2_R2278_U70); 
assign P2_R2278_U461 = ~(P2_U2798 & P2_R2278_U70); 
assign P2_R2278_U465 = ~(P2_R2278_U37 & P2_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P2_R2278_U467 = ~(P2_R2278_U37 & P2_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P2_R2278_U476 = ~(P2_R2278_U475 & P2_R2278_U474); 
assign P2_ADD_394_U56 = ~(P2_ADD_394_U121 & P2_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P2_ADD_394_U156 = ~(P2_ADD_394_U121 & P2_ADD_394_U55); 
assign P2_R2267_U13 = P2_R2267_U119 & P2_R2267_U38; 
assign P2_R2267_U39 = ~(P2_R2267_U53 & P2_R2267_U109); 
assign P2_R2267_U116 = ~(P2_R2267_U109 & P2_R2267_U68); 
assign P2_R2267_U148 = ~(P2_R2267_U109 & P2_R2267_U68); 
assign P2_ADD_371_1212_U125 = ~(P2_ADD_371_1212_U151 & P2_ADD_371_1212_U150); 
assign P2_ADD_371_1212_U126 = P2_ADD_371_1212_U250 & P2_ADD_371_1212_U249; 
assign P2_ADD_371_1212_U207 = ~(P2_ADD_371_1212_U40 & P2_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P2_ADD_371_1212_U209 = ~(P2_ADD_371_1212_U40 & P2_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P2_ADD_371_1212_U239 = ~(P2_ADD_371_1212_U148 & P2_ADD_371_1212_U237); 
assign P2_ADD_371_1212_U253 = ~(P2_ADD_371_1212_U252 & P2_ADD_371_1212_U251); 
assign P1_R2278_U98 = ~(P1_R2278_U138 & P1_R2278_U354); 
assign P1_R2278_U257 = ~P1_R2278_U178; 
assign P1_R2278_U260 = ~P1_R2278_U176; 
assign P1_R2278_U268 = ~(P1_R2278_U255 & P1_R2278_U267); 
assign P1_R2278_U274 = ~(P1_R2278_U261 & P1_R2278_U176); 
assign P1_R2278_U430 = ~(P1_R2278_U346 & P1_R2278_U176); 
assign P1_R2278_U437 = ~(P1_R2278_U177 & P1_R2278_U178); 
assign P1_R2358_U14 = P1_R2358_U330 & P1_R2358_U329; 
assign P1_R2358_U15 = P1_R2358_U327 & P1_R2358_U325; 
assign P1_R2358_U42 = ~(P1_U2627 & P1_R2358_U546); 
assign P1_R2358_U72 = ~(P1_R2358_U71 & P1_R2358_U255); 
assign P1_R2358_U117 = ~(P1_R2358_U607 & P1_R2358_U606); 
assign P1_R2358_U194 = ~(P1_R2358_U129 & P1_R2358_U393); 
assign P1_R2358_U195 = ~(P1_R2358_U359 & P1_R2358_U395); 
assign P1_R2358_U196 = ~(P1_R2358_U397 & P1_R2358_U51); 
assign P1_R2358_U312 = ~P1_R2358_U71; 
assign P1_R2358_U530 = ~(P1_U2352 & P1_R2358_U174); 
assign P1_R2358_U541 = ~(P1_U2352 & P1_R2358_U174); 
assign P1_R2358_U605 = ~(P1_R2358_U114 & P1_R2358_U271); 
assign P1_R2099_U23 = ~(P1_R2099_U177 & P1_R2099_U47); 
assign P1_R2099_U304 = ~(P1_R2099_U234 & P1_R2099_U177); 
assign P1_R2337_U56 = ~(P1_R2337_U118 & P1_PHYADDRPOINTER_REG_27__SCAN_IN); 
assign P1_R2337_U148 = ~(P1_R2337_U118 & P1_R2337_U55); 
assign P1_R2096_U56 = ~(P1_R2096_U118 & P1_REIP_REG_27__SCAN_IN); 
assign P1_R2096_U148 = ~(P1_R2096_U118 & P1_R2096_U55); 
assign P1_ADD_405_U56 = ~(P1_ADD_405_U121 & P1_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P1_ADD_405_U156 = ~(P1_ADD_405_U121 & P1_ADD_405_U55); 
assign P1_ADD_515_U56 = ~(P1_ADD_515_U118 & P1_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P1_ADD_515_U154 = ~(P1_ADD_515_U118 & P1_ADD_515_U55); 
assign P3_U2839 = ~(P3_U3873 & P3_U6206); 
assign P3_U3884 = P3_U6236 & P3_U6235; 
assign P3_U3886 = P3_U6238 & P3_U6237 & P3_U6239 & P3_U3885; 
assign P3_U3890 = P3_U6248 & P3_U6247 & P3_U6249; 
assign P3_U3891 = P3_U6251 & P3_U6250; 
assign P3_U3896 = P3_U6265 & P3_U6264; 
assign P3_U3898 = P3_U6267 & P3_U6266 & P3_U6268; 
assign P3_U3899 = P3_U6270 & P3_U6269; 
assign P3_U3980 = P3_U6620 & P3_U6619 & P3_U6618 & P3_U6617; 
assign P3_U4117 = P3_U7318 & P3_U7317; 
assign P3_U6228 = ~(P3_U3882 & P3_U3877); 
assign P3_U6280 = ~(P3_ADD_360_1242_U78 & P3_U2395); 
assign P3_U6323 = ~(P3_ADD_371_1212_U16 & P3_U2360); 
assign P3_U6623 = ~(P3_U2396 & P3_ADD_360_1242_U78); 
assign P3_U6635 = ~(P3_U2387 & P3_ADD_371_1212_U16); 
assign P2_U2796 = P2_U3242 & P2_R2267_U13; 
assign P2_U2910 = ~(P2_U4068 & P2_U6363 & P2_U6364); 
assign P2_U3663 = ~(P2_U8382 & P2_U8381); 
assign P2_U6368 = ~(P2_ADD_391_1196_U109 & P2_U2397); 
assign P2_U6449 = ~(P2_U2380 & P2_R2096_U80); 
assign P2_U6520 = ~(P2_U2379 & P2_R2099_U87); 
assign P2_U6531 = ~(P2_R2182_U86 & P2_U2393); 
assign P2_U6710 = ~(P2_U2392 & P2_R2099_U87); 
assign P2_U6779 = ~(P2_R2267_U13 & P2_U2587); 
assign P2_U6796 = ~(P2_U2588 & P2_R2096_U80); 
assign P2_U8315 = ~(P2_R2256_U17 & P2_U3572); 
assign P1_U3844 = P1_U5753 & P1_U5755; 
assign P1_U3846 = P1_U3845 & P1_U5756; 
assign P1_U3938 = P1_U6559 & P1_U6557; 
assign P1_U4014 = P1_U6793 & P1_U6794 & P1_U6795; 
assign P1_U5852 = ~(P1_R2358_U14 & P1_U2364); 
assign P1_U5857 = ~(P1_R2358_U15 & P1_U2364); 
assign P1_U5867 = ~(P1_R2358_U117 & P1_U2364); 
assign P1_U6185 = ~(P1_U2386 & P1_R2358_U14); 
assign P1_U6188 = ~(P1_U2386 & P1_R2358_U15); 
assign P1_U6194 = ~(P1_U2386 & P1_R2358_U117); 
assign P1_U6295 = ~(P1_U2383 & P1_R2358_U14); 
assign P1_U6298 = ~(P1_U2383 & P1_R2358_U15); 
assign P1_U6304 = ~(P1_U2383 & P1_R2358_U117); 
assign P3_ADD_476_U74 = ~(P3_ADD_476_U148 & P3_ADD_476_U147); 
assign P3_ADD_476_U119 = ~P3_ADD_476_U56; 
assign P3_ADD_476_U145 = ~(P3_ADD_476_U56 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_531_U78 = ~(P3_ADD_531_U155 & P3_ADD_531_U154); 
assign P3_ADD_531_U123 = ~P3_ADD_531_U57; 
assign P3_ADD_531_U152 = ~(P3_ADD_531_U57 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_SUB_320_U36 = ~(P3_SUB_320_U41 & P3_SUB_320_U65 & P3_SUB_320_U100); 
assign P3_ADD_318_U74 = ~(P3_ADD_318_U148 & P3_ADD_318_U147); 
assign P3_ADD_318_U119 = ~P3_ADD_318_U56; 
assign P3_ADD_318_U145 = ~(P3_ADD_318_U56 & P3_PHYADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_315_U70 = ~(P3_ADD_315_U140 & P3_ADD_315_U139); 
assign P3_ADD_315_U116 = ~P3_ADD_315_U56; 
assign P3_ADD_315_U137 = ~(P3_ADD_315_U56 & P3_PHYADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_360_1242_U15 = P3_ADD_360_1242_U168 & P3_ADD_360_1242_U71; 
assign P3_ADD_360_1242_U73 = ~(P3_ADD_360_1242_U164 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_467_U74 = ~(P3_ADD_467_U148 & P3_ADD_467_U147); 
assign P3_ADD_467_U119 = ~P3_ADD_467_U56; 
assign P3_ADD_467_U145 = ~(P3_ADD_467_U56 & P3_REIP_REG_28__SCAN_IN); 
assign P3_ADD_430_U74 = ~(P3_ADD_430_U148 & P3_ADD_430_U147); 
assign P3_ADD_430_U119 = ~P3_ADD_430_U56; 
assign P3_ADD_430_U145 = ~(P3_ADD_430_U56 & P3_REIP_REG_28__SCAN_IN); 
assign P3_ADD_380_U78 = ~(P3_ADD_380_U155 & P3_ADD_380_U154); 
assign P3_ADD_380_U123 = ~P3_ADD_380_U57; 
assign P3_ADD_380_U152 = ~(P3_ADD_380_U57 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_344_U78 = ~(P3_ADD_344_U155 & P3_ADD_344_U154); 
assign P3_ADD_344_U123 = ~P3_ADD_344_U57; 
assign P3_ADD_344_U152 = ~(P3_ADD_344_U57 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_339_U74 = ~(P3_ADD_339_U148 & P3_ADD_339_U147); 
assign P3_ADD_339_U119 = ~P3_ADD_339_U56; 
assign P3_ADD_339_U145 = ~(P3_ADD_339_U56 & P3_PHYADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_541_U74 = ~(P3_ADD_541_U148 & P3_ADD_541_U147); 
assign P3_ADD_541_U119 = ~P3_ADD_541_U56; 
assign P3_ADD_541_U145 = ~(P3_ADD_541_U56 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_515_U74 = ~(P3_ADD_515_U148 & P3_ADD_515_U147); 
assign P3_ADD_515_U119 = ~P3_ADD_515_U56; 
assign P3_ADD_515_U145 = ~(P3_ADD_515_U56 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_394_U73 = ~(P3_ADD_394_U150 & P3_ADD_394_U149); 
assign P3_ADD_394_U122 = ~P3_ADD_394_U56; 
assign P3_ADD_394_U147 = ~(P3_ADD_394_U56 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_441_U74 = ~(P3_ADD_441_U148 & P3_ADD_441_U147); 
assign P3_ADD_441_U119 = ~P3_ADD_441_U56; 
assign P3_ADD_441_U145 = ~(P3_ADD_441_U56 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_349_U78 = ~(P3_ADD_349_U155 & P3_ADD_349_U154); 
assign P3_ADD_349_U123 = ~P3_ADD_349_U57; 
assign P3_ADD_349_U152 = ~(P3_ADD_349_U57 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_405_U73 = ~(P3_ADD_405_U150 & P3_ADD_405_U149); 
assign P3_ADD_405_U122 = ~P3_ADD_405_U56; 
assign P3_ADD_405_U147 = ~(P3_ADD_405_U56 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_553_U78 = ~(P3_ADD_553_U155 & P3_ADD_553_U154); 
assign P3_ADD_553_U123 = ~P3_ADD_553_U57; 
assign P3_ADD_553_U152 = ~(P3_ADD_553_U57 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_558_U78 = ~(P3_ADD_558_U155 & P3_ADD_558_U154); 
assign P3_ADD_558_U123 = ~P3_ADD_558_U57; 
assign P3_ADD_558_U152 = ~(P3_ADD_558_U57 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_385_U78 = ~(P3_ADD_385_U155 & P3_ADD_385_U154); 
assign P3_ADD_385_U123 = ~P3_ADD_385_U57; 
assign P3_ADD_385_U152 = ~(P3_ADD_385_U57 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_547_U78 = ~(P3_ADD_547_U155 & P3_ADD_547_U154); 
assign P3_ADD_547_U123 = ~P3_ADD_547_U57; 
assign P3_ADD_547_U152 = ~(P3_ADD_547_U57 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_371_1212_U17 = P3_ADD_371_1212_U176 & P3_ADD_371_1212_U75; 
assign P3_ADD_371_1212_U174 = ~P3_ADD_371_1212_U75; 
assign P3_ADD_371_1212_U238 = ~(P3_ADD_371_1212_U75 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_494_U74 = ~(P3_ADD_494_U148 & P3_ADD_494_U147); 
assign P3_ADD_494_U119 = ~P3_ADD_494_U56; 
assign P3_ADD_494_U145 = ~(P3_ADD_494_U56 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_536_U74 = ~(P3_ADD_536_U148 & P3_ADD_536_U147); 
assign P3_ADD_536_U119 = ~P3_ADD_536_U56; 
assign P3_ADD_536_U145 = ~(P3_ADD_536_U56 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P2_R2099_U41 = ~(P2_U2730 & P2_R2099_U132); 
assign P2_R2099_U209 = ~(P2_R2099_U132 & P2_R2099_U40); 
assign P2_ADD_391_1196_U62 = ~P2_R2182_U86; 
assign P2_ADD_391_1196_U77 = ~P2_R2096_U80; 
assign P2_ADD_391_1196_U147 = P2_ADD_391_1196_U434 & P2_ADD_391_1196_U433; 
assign P2_ADD_391_1196_U156 = ~(P2_ADD_391_1196_U86 & P2_ADD_391_1196_U212); 
assign P2_ADD_391_1196_U211 = ~P2_ADD_391_1196_U86; 
assign P2_ADD_391_1196_U244 = P2_R2182_U86 | P2_R2096_U87; 
assign P2_ADD_391_1196_U246 = ~(P2_R2096_U87 & P2_R2182_U86); 
assign P2_ADD_391_1196_U415 = ~(P2_R2182_U86 & P2_ADD_391_1196_U63); 
assign P2_ADD_391_1196_U417 = ~(P2_R2182_U86 & P2_ADD_391_1196_U63); 
assign P2_ADD_391_1196_U426 = ~(P2_R2096_U88 & P2_ADD_391_1196_U60); 
assign P2_ADD_391_1196_U428 = ~(P2_R2096_U88 & P2_ADD_391_1196_U60); 
assign P2_ADD_391_1196_U437 = ~(P2_ADD_391_1196_U436 & P2_ADD_391_1196_U435); 
assign P2_R2182_U85 = ~(P2_R2182_U276 & P2_R2182_U275); 
assign P2_R2182_U154 = ~P2_R2182_U7; 
assign P2_R2182_U156 = ~(P2_R2182_U155 & P2_R2182_U7); 
assign P2_R2182_U271 = ~(P2_R2182_U120 & P2_R2182_U7); 
assign P2_R2182_U274 = ~(P2_R2182_U153 & P2_U2690); 
assign P2_R2027_U78 = ~(P2_R2027_U155 & P2_R2027_U154); 
assign P2_R2027_U123 = ~P2_R2027_U57; 
assign P2_R2027_U152 = ~(P2_R2027_U57 & P2_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P2_R2337_U72 = ~(P2_R2337_U146 & P2_R2337_U145); 
assign P2_R2337_U120 = ~P2_R2337_U57; 
assign P2_R2337_U143 = ~(P2_R2337_U57 & P2_PHYADDRPOINTER_REG_29__SCAN_IN); 
assign P2_R2096_U79 = ~(P2_R2096_U222 & P2_R2096_U221); 
assign P2_R2096_U165 = ~P2_R2096_U22; 
assign P2_R2096_U166 = ~(P2_U2619 & P2_R2096_U22); 
assign P2_R2096_U168 = ~(P2_R2096_U98 & P2_R2096_U22); 
assign P2_R2096_U210 = ~(P2_R2096_U30 & P2_R2096_U22); 
assign P2_R2096_U220 = ~(P2_R2096_U164 & P2_U2620); 
assign P2_R1957_U35 = ~(P2_R1957_U100 & P2_R1957_U65 & P2_R1957_U40); 
assign P2_R2278_U24 = ~P2_U3632; 
assign P2_R2278_U26 = ~(P2_U3632 & P2_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P2_R2278_U35 = ~P2_U2797; 
assign P2_R2278_U116 = P2_R2278_U316 & P2_R2278_U222; 
assign P2_R2278_U119 = P2_R2278_U231 & P2_R2278_U235; 
assign P2_R2278_U133 = P2_R2278_U336 & P2_R2278_U281; 
assign P2_R2278_U153 = P2_R2278_U375 & P2_R2278_U374; 
assign P2_R2278_U154 = ~(P2_R2278_U23 & P2_R2278_U218); 
assign P2_R2278_U179 = P2_R2278_U466 & P2_R2278_U465; 
assign P2_R2278_U224 = P2_U3632 | P2_INSTADDRPOINTER_REG_6__SCAN_IN; 
assign P2_R2278_U233 = ~P2_R2278_U49; 
assign P2_R2278_U285 = ~P2_R2278_U71; 
assign P2_R2278_U287 = P2_U2797 | P2_INSTADDRPOINTER_REG_24__SCAN_IN; 
assign P2_R2278_U288 = ~(P2_U2797 & P2_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P2_R2278_U315 = ~(P2_R2278_U115 & P2_R2278_U156); 
assign P2_R2278_U353 = ~(P2_R2278_U27 & P2_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P2_R2278_U355 = ~(P2_R2278_U27 & P2_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P2_R2278_U368 = ~(P2_U3632 & P2_R2278_U25); 
assign P2_R2278_U370 = ~(P2_U3632 & P2_R2278_U25); 
assign P2_R2278_U378 = ~(P2_R2278_U377 & P2_R2278_U376); 
assign P2_R2278_U387 = ~(P2_R2278_U216 & P2_R2278_U385); 
assign P2_R2278_U452 = ~(P2_U2797 & P2_R2278_U36); 
assign P2_R2278_U454 = ~(P2_U2797 & P2_R2278_U36); 
assign P2_R2278_U458 = ~(P2_R2278_U69 & P2_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P2_R2278_U460 = ~(P2_R2278_U69 & P2_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P2_R2278_U469 = ~(P2_R2278_U468 & P2_R2278_U467); 
assign P2_ADD_394_U77 = ~(P2_ADD_394_U156 & P2_ADD_394_U155); 
assign P2_ADD_394_U122 = ~P2_ADD_394_U56; 
assign P2_ADD_394_U175 = ~(P2_ADD_394_U56 & P2_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P2_R2267_U69 = P2_R2267_U148 & P2_R2267_U147; 
assign P2_R2267_U110 = ~P2_R2267_U39; 
assign P2_R2267_U117 = ~(P2_U2770 & P2_R2267_U116); 
assign P2_R2267_U145 = ~(P2_U2769 & P2_R2267_U39); 
assign P2_ADD_371_1212_U43 = ~P2_R2256_U17; 
assign P2_ADD_371_1212_U80 = ~(P2_ADD_371_1212_U239 & P2_ADD_371_1212_U238); 
assign P2_ADD_371_1212_U110 = P2_ADD_371_1212_U208 & P2_ADD_371_1212_U207; 
assign P2_ADD_371_1212_U152 = ~P2_ADD_371_1212_U125; 
assign P2_ADD_371_1212_U154 = ~(P2_ADD_371_1212_U153 & P2_ADD_371_1212_U125); 
assign P2_ADD_371_1212_U161 = P2_R2256_U17 | P2_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P2_ADD_371_1212_U163 = ~(P2_R2256_U17 & P2_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P2_ADD_371_1212_U203 = ~(P2_ADD_371_1212_U165 & P2_R2256_U17 & P2_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P2_ADD_371_1212_U211 = ~(P2_ADD_371_1212_U210 & P2_ADD_371_1212_U209); 
assign P2_ADD_371_1212_U247 = ~(P2_ADD_371_1212_U124 & P2_ADD_371_1212_U125); 
assign P2_ADD_371_1212_U275 = ~(P2_R2256_U17 & P2_ADD_371_1212_U44); 
assign P2_ADD_371_1212_U277 = ~(P2_R2256_U17 & P2_ADD_371_1212_U44); 
assign P1_R2278_U18 = P1_R2278_U268 & P1_R2278_U266; 
assign P1_R2278_U224 = ~(P1_R2278_U98 & P1_R2278_U279); 
assign P1_R2278_U225 = ~(P1_R2278_U274 & P1_R2278_U273); 
assign P1_R2278_U278 = ~P1_R2278_U98; 
assign P1_R2278_U431 = ~(P1_R2278_U100 & P1_R2278_U260); 
assign P1_R2278_U438 = ~(P1_R2278_U257 & P1_R2278_U436); 
assign P1_R2358_U98 = P1_R2358_U42 & P1_R2358_U286; 
assign P1_R2358_U115 = ~(P1_R2358_U605 & P1_R2358_U604); 
assign P1_R2358_U172 = ~P1_U2657; 
assign P1_R2358_U287 = ~P1_R2358_U42; 
assign P1_R2358_U288 = ~(P1_R2358_U531 & P1_R2358_U530 & P1_R2358_U40); 
assign P1_R2358_U313 = ~P1_R2358_U72; 
assign P1_R2358_U314 = ~(P1_R2358_U72 & P1_R2358_U61); 
assign P1_R2358_U317 = ~(P1_R2358_U140 & P1_R2358_U72); 
assign P1_R2358_U319 = ~(P1_R2358_U312 & P1_R2358_U318); 
assign P1_R2358_U342 = ~(P1_R2358_U42 & P1_R2358_U286); 
assign P1_R2358_U385 = ~(P1_R2358_U130 & P1_R2358_U194); 
assign P1_R2358_U387 = ~(P1_R2358_U7 & P1_R2358_U194); 
assign P1_R2358_U389 = ~(P1_R2358_U6 & P1_R2358_U194); 
assign P1_R2358_U391 = ~(P1_R2358_U278 & P1_R2358_U194); 
assign P1_R2358_U394 = ~P1_R2358_U194; 
assign P1_R2358_U396 = ~P1_R2358_U195; 
assign P1_R2358_U398 = ~P1_R2358_U196; 
assign P1_R2358_U527 = ~(P1_U2657 & P1_R2358_U23); 
assign P1_R2358_U539 = ~(P1_U2657 & P1_R2358_U23); 
assign P1_R2358_U543 = ~(P1_R2358_U542 & P1_R2358_U541); 
assign P1_R2358_U598 = ~(P1_R2358_U194 & P1_R2358_U347); 
assign P1_R2358_U600 = ~(P1_R2358_U195 & P1_R2358_U348); 
assign P1_R2358_U602 = ~(P1_R2358_U196 & P1_R2358_U349); 
assign P1_R2099_U69 = ~(P1_R2099_U305 & P1_R2099_U304); 
assign P1_R2099_U178 = ~P1_R2099_U23; 
assign P1_R2099_U303 = ~(P1_R2099_U46 & P1_R2099_U23); 
assign P1_R2337_U74 = ~(P1_R2337_U148 & P1_R2337_U147); 
assign P1_R2337_U119 = ~P1_R2337_U56; 
assign P1_R2337_U145 = ~(P1_R2337_U56 & P1_PHYADDRPOINTER_REG_28__SCAN_IN); 
assign P1_R2096_U74 = ~(P1_R2096_U148 & P1_R2096_U147); 
assign P1_R2096_U119 = ~P1_R2096_U56; 
assign P1_R2096_U145 = ~(P1_R2096_U56 & P1_REIP_REG_28__SCAN_IN); 
assign P1_ADD_405_U77 = ~(P1_ADD_405_U156 & P1_ADD_405_U155); 
assign P1_ADD_405_U122 = ~P1_ADD_405_U56; 
assign P1_ADD_405_U175 = ~(P1_ADD_405_U56 & P1_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P1_ADD_515_U77 = ~(P1_ADD_515_U154 & P1_ADD_515_U153); 
assign P1_ADD_515_U119 = ~P1_ADD_515_U56; 
assign P1_ADD_515_U171 = ~(P1_ADD_515_U56 & P1_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_U2804 = ~(P3_U6614 & P3_U6616 & P3_U6613 & P3_U6615 & P3_U3980); 
assign P3_U3887 = P3_U6233 & P3_U6234 & P3_U6232 & P3_U3884 & P3_U3886; 
assign P3_U3892 = P3_U3889 & P3_U3888 & P3_U3891 & P3_U3890; 
assign P3_U3903 = P3_U6281 & P3_U6280; 
assign P3_U6230 = ~(P3_U4318 & P3_U6228); 
assign P3_U6258 = ~(P3_ADD_558_U78 & P3_U3220); 
assign P3_U6259 = ~(P3_ADD_553_U78 & P3_U4298); 
assign P3_U6260 = ~(P3_ADD_547_U78 & P3_U4299); 
assign P3_U6263 = ~(P3_ADD_531_U78 & P3_U2354); 
assign P3_U6271 = ~(P3_ADD_385_U78 & P3_U2358); 
assign P3_U6272 = ~(P3_ADD_380_U78 & P3_U2359); 
assign P3_U6273 = ~(P3_ADD_349_U78 & P3_U4306); 
assign P3_U6274 = ~(P3_ADD_344_U78 & P3_U2362); 
assign P3_U6285 = ~(P3_ADD_541_U74 & P3_U4300); 
assign P3_U6286 = ~(P3_ADD_536_U74 & P3_U4301); 
assign P3_U6289 = ~(P3_ADD_515_U74 & P3_U4302); 
assign P3_U6290 = ~(P3_ADD_494_U74 & P3_U2356); 
assign P3_U6291 = ~(P3_ADD_476_U74 & P3_U4303); 
assign P3_U6292 = ~(P3_ADD_441_U74 & P3_U4304); 
assign P3_U6293 = ~(P3_ADD_405_U73 & P3_U4305); 
assign P3_U6294 = ~(P3_ADD_394_U73 & P3_U2357); 
assign P3_U6304 = ~(P3_ADD_360_1242_U15 & P3_U2395); 
assign P3_U6347 = ~(P3_ADD_371_1212_U17 & P3_U2360); 
assign P3_U6621 = ~(P3_ADD_318_U74 & P3_U2398); 
assign P3_U6626 = ~(P3_ADD_339_U74 & P3_U2388); 
assign P3_U6630 = ~(P3_ADD_315_U70 & P3_U2397); 
assign P3_U6631 = ~(P3_U2396 & P3_ADD_360_1242_U15); 
assign P3_U6643 = ~(P3_U2387 & P3_ADD_371_1212_U17); 
assign P3_U7326 = ~(P3_ADD_467_U74 & P3_U2601); 
assign P3_U7328 = ~(P3_ADD_430_U74 & P3_U2405); 
assign P2_U2795 = P2_U3242 & P2_R2267_U69; 
assign P2_U2871 = ~(P2_U6520 & P2_U6521 & P2_U6519); 
assign P2_U2909 = ~(P2_U6370 & P2_U6367 & P2_U6369 & P2_U6368); 
assign P2_U3631 = ~(P2_U8316 & P2_U8315); 
assign P2_U6454 = ~(P2_U2380 & P2_R2096_U79); 
assign P2_U6534 = ~(P2_R2182_U85 & P2_U2393); 
assign P2_U6787 = ~(P2_R2267_U69 & P2_U2587); 
assign P2_U6804 = ~(P2_U2588 & P2_R2096_U79); 
assign P2_U8379 = ~(P2_R2337_U72 & P2_U3284); 
assign P1_U2656 = ~(P1_U6792 & P1_U4014); 
assign P1_U2859 = ~(P1_U6305 & P1_U6306 & P1_U6304); 
assign P1_U2861 = ~(P1_U6299 & P1_U6300 & P1_U6298); 
assign P1_U2862 = ~(P1_U6296 & P1_U6297 & P1_U6295); 
assign P1_U2891 = ~(P1_U6195 & P1_U6193 & P1_U6194); 
assign P1_U2893 = ~(P1_U6189 & P1_U6187 & P1_U6188); 
assign P1_U2894 = ~(P1_U6186 & P1_U6184 & P1_U6185); 
assign P1_U5621 = ~(P1_R2278_U18 & P1_U2377); 
assign P1_U5752 = ~(P1_R2099_U69 & P1_U2380); 
assign P1_U5762 = ~(P1_ADD_405_U77 & P1_U2375); 
assign P1_U5763 = ~(P1_ADD_515_U77 & P1_U2374); 
assign P1_U5835 = ~(P1_U2372 & P1_R2278_U18); 
assign P1_U5882 = ~(P1_R2358_U115 & P1_U2364); 
assign P1_U5934 = ~(P1_R2337_U74 & P1_U2376); 
assign P1_U6204 = ~(P1_U2386 & P1_R2358_U115); 
assign P1_U6313 = ~(P1_U2383 & P1_R2358_U115); 
assign P1_U6344 = ~(P1_U2371 & P1_R2099_U69); 
assign P1_U6556 = ~(P1_U2604 & P1_R2099_U69); 
assign P1_U6564 = ~(P1_R2096_U74 & P1_U7485); 
assign P1_U6791 = ~(P1_R2337_U74 & P1_U2352); 
assign P3_ADD_476_U58 = ~(P3_ADD_476_U119 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_476_U146 = ~(P3_ADD_476_U119 & P3_ADD_476_U57); 
assign P3_ADD_531_U59 = ~(P3_ADD_531_U123 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_531_U153 = ~(P3_ADD_531_U123 & P3_ADD_531_U58); 
assign P3_SUB_320_U14 = P3_SUB_320_U110 & P3_SUB_320_U36; 
assign P3_SUB_320_U63 = ~P3_ADD_318_U74; 
assign P3_SUB_320_U101 = ~P3_SUB_320_U36; 
assign P3_SUB_320_U140 = ~(P3_ADD_318_U74 & P3_SUB_320_U36); 
assign P3_ADD_318_U58 = ~(P3_ADD_318_U119 & P3_PHYADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_318_U146 = ~(P3_ADD_318_U119 & P3_ADD_318_U57); 
assign P3_ADD_315_U58 = ~(P3_ADD_315_U116 & P3_PHYADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_315_U138 = ~(P3_ADD_315_U116 & P3_ADD_315_U57); 
assign P3_ADD_360_1242_U16 = P3_ADD_360_1242_U166 & P3_ADD_360_1242_U73; 
assign P3_ADD_360_1242_U165 = ~P3_ADD_360_1242_U73; 
assign P3_ADD_360_1242_U229 = ~(P3_ADD_360_1242_U73 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_467_U58 = ~(P3_ADD_467_U119 & P3_REIP_REG_28__SCAN_IN); 
assign P3_ADD_467_U146 = ~(P3_ADD_467_U119 & P3_ADD_467_U57); 
assign P3_ADD_430_U58 = ~(P3_ADD_430_U119 & P3_REIP_REG_28__SCAN_IN); 
assign P3_ADD_430_U146 = ~(P3_ADD_430_U119 & P3_ADD_430_U57); 
assign P3_ADD_380_U59 = ~(P3_ADD_380_U123 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_380_U153 = ~(P3_ADD_380_U123 & P3_ADD_380_U58); 
assign P3_ADD_344_U59 = ~(P3_ADD_344_U123 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_344_U153 = ~(P3_ADD_344_U123 & P3_ADD_344_U58); 
assign P3_ADD_339_U58 = ~(P3_ADD_339_U119 & P3_PHYADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_339_U146 = ~(P3_ADD_339_U119 & P3_ADD_339_U57); 
assign P3_ADD_541_U58 = ~(P3_ADD_541_U119 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_541_U146 = ~(P3_ADD_541_U119 & P3_ADD_541_U57); 
assign P3_ADD_515_U58 = ~(P3_ADD_515_U119 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_515_U146 = ~(P3_ADD_515_U119 & P3_ADD_515_U57); 
assign P3_ADD_394_U58 = ~(P3_ADD_394_U122 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_394_U148 = ~(P3_ADD_394_U122 & P3_ADD_394_U57); 
assign P3_ADD_441_U58 = ~(P3_ADD_441_U119 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_441_U146 = ~(P3_ADD_441_U119 & P3_ADD_441_U57); 
assign P3_ADD_349_U59 = ~(P3_ADD_349_U123 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_349_U153 = ~(P3_ADD_349_U123 & P3_ADD_349_U58); 
assign P3_ADD_405_U58 = ~(P3_ADD_405_U122 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_405_U148 = ~(P3_ADD_405_U122 & P3_ADD_405_U57); 
assign P3_ADD_553_U59 = ~(P3_ADD_553_U123 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_553_U153 = ~(P3_ADD_553_U123 & P3_ADD_553_U58); 
assign P3_ADD_558_U59 = ~(P3_ADD_558_U123 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_558_U153 = ~(P3_ADD_558_U123 & P3_ADD_558_U58); 
assign P3_ADD_385_U59 = ~(P3_ADD_385_U123 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_385_U153 = ~(P3_ADD_385_U123 & P3_ADD_385_U58); 
assign P3_ADD_547_U59 = ~(P3_ADD_547_U123 & P3_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P3_ADD_547_U153 = ~(P3_ADD_547_U123 & P3_ADD_547_U58); 
assign P3_ADD_371_1212_U198 = ~(P3_ADD_371_1212_U174 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_371_1212_U237 = ~(P3_ADD_371_1212_U174 & P3_ADD_371_1212_U116 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_371_1212_U239 = ~(P3_ADD_371_1212_U174 & P3_ADD_371_1212_U76); 
assign P3_ADD_494_U58 = ~(P3_ADD_494_U119 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_494_U146 = ~(P3_ADD_494_U119 & P3_ADD_494_U57); 
assign P3_ADD_536_U58 = ~(P3_ADD_536_U119 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_536_U146 = ~(P3_ADD_536_U119 & P3_ADD_536_U57); 
assign P2_R2099_U86 = ~(P2_R2099_U209 & P2_R2099_U208); 
assign P2_R2099_U133 = ~P2_R2099_U41; 
assign P2_R2099_U206 = ~(P2_U2729 & P2_R2099_U41); 
assign P2_ADD_391_1196_U64 = ~P2_R2182_U85; 
assign P2_ADD_391_1196_U78 = ~P2_R2096_U79; 
assign P2_ADD_391_1196_U145 = P2_ADD_391_1196_U427 & P2_ADD_391_1196_U426; 
assign P2_ADD_391_1196_U213 = ~P2_ADD_391_1196_U156; 
assign P2_ADD_391_1196_U215 = ~(P2_ADD_391_1196_U214 & P2_ADD_391_1196_U156); 
assign P2_ADD_391_1196_U248 = P2_R2182_U85 | P2_R2096_U86; 
assign P2_ADD_391_1196_U250 = ~(P2_R2096_U86 & P2_R2182_U85); 
assign P2_ADD_391_1196_U301 = ~(P2_ADD_391_1196_U211 & P2_ADD_391_1196_U300); 
assign P2_ADD_391_1196_U408 = ~(P2_R2182_U85 & P2_ADD_391_1196_U65); 
assign P2_ADD_391_1196_U410 = ~(P2_R2182_U85 & P2_ADD_391_1196_U65); 
assign P2_ADD_391_1196_U414 = ~(P2_R2096_U87 & P2_ADD_391_1196_U62); 
assign P2_ADD_391_1196_U416 = ~(P2_R2096_U87 & P2_ADD_391_1196_U62); 
assign P2_ADD_391_1196_U430 = ~(P2_ADD_391_1196_U429 & P2_ADD_391_1196_U428); 
assign P2_ADD_391_1196_U468 = ~(P2_ADD_391_1196_U155 & P2_ADD_391_1196_U156); 
assign P2_R2182_U84 = ~(P2_R2182_U274 & P2_R2182_U273); 
assign P2_R2182_U119 = ~(P2_R2182_U157 & P2_R2182_U156); 
assign P2_R2182_U272 = ~(P2_R2182_U154 & P2_R2182_U270); 
assign P2_R2027_U59 = ~(P2_R2027_U123 & P2_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P2_R2027_U153 = ~(P2_R2027_U123 & P2_R2027_U58); 
assign P2_R2337_U59 = ~(P2_R2337_U120 & P2_PHYADDRPOINTER_REG_29__SCAN_IN); 
assign P2_R2337_U144 = ~(P2_R2337_U120 & P2_R2337_U58); 
assign P2_R2096_U78 = ~(P2_R2096_U220 & P2_R2096_U219); 
assign P2_R2096_U167 = ~(P2_R2096_U29 & P2_R2096_U166); 
assign P2_R2096_U211 = ~(P2_U2619 & P2_R2096_U165); 
assign P2_R1957_U14 = P2_R1957_U110 & P2_R1957_U35; 
assign P2_R1957_U63 = ~P2_U3663; 
assign P2_R1957_U101 = ~P2_R1957_U35; 
assign P2_R1957_U140 = ~(P2_U3663 & P2_R1957_U35); 
assign P2_R2278_U72 = ~P2_U2796; 
assign P2_R2278_U89 = ~(P2_R2278_U387 & P2_R2278_U386); 
assign P2_R2278_U134 = P2_R2278_U283 & P2_R2278_U287; 
assign P2_R2278_U147 = P2_R2278_U354 & P2_R2278_U353; 
assign P2_R2278_U152 = ~(P2_R2278_U116 & P2_R2278_U315); 
assign P2_R2278_U177 = P2_R2278_U459 & P2_R2278_U458; 
assign P2_R2278_U220 = ~P2_R2278_U154; 
assign P2_R2278_U226 = ~P2_R2278_U26; 
assign P2_R2278_U308 = ~(P2_U2796 & P2_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P2_R2278_U320 = ~(P2_R2278_U233 & P2_R2278_U235); 
assign P2_R2278_U338 = ~(P2_R2278_U285 & P2_R2278_U287); 
assign P2_R2278_U357 = ~(P2_R2278_U356 & P2_R2278_U355); 
assign P2_R2278_U367 = ~(P2_R2278_U24 & P2_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P2_R2278_U369 = ~(P2_R2278_U24 & P2_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P2_R2278_U379 = ~(P2_R2278_U153 & P2_R2278_U154); 
assign P2_R2278_U451 = ~(P2_R2278_U35 & P2_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P2_R2278_U453 = ~(P2_R2278_U35 & P2_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P2_R2278_U462 = ~(P2_R2278_U461 & P2_R2278_U460); 
assign P2_ADD_394_U58 = ~(P2_ADD_394_U122 & P2_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P2_ADD_394_U176 = ~(P2_ADD_394_U122 & P2_ADD_394_U57); 
assign P2_R2267_U14 = P2_R2267_U117 & P2_R2267_U39; 
assign P2_R2267_U40 = ~(P2_R2267_U54 & P2_R2267_U110); 
assign P2_R2267_U114 = ~(P2_R2267_U110 & P2_R2267_U66); 
assign P2_R2267_U146 = ~(P2_R2267_U110 & P2_R2267_U66); 
assign P2_ADD_371_1212_U86 = P2_ADD_371_1212_U203 & P2_ADD_371_1212_U166; 
assign P2_ADD_371_1212_U111 = ~(P2_ADD_371_1212_U155 & P2_ADD_371_1212_U154); 
assign P2_ADD_371_1212_U248 = ~(P2_ADD_371_1212_U152 & P2_ADD_371_1212_U246); 
assign P2_ADD_371_1212_U274 = ~(P2_ADD_371_1212_U43 & P2_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P2_ADD_371_1212_U276 = ~(P2_ADD_371_1212_U43 & P2_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P1_R2278_U101 = ~(P1_R2278_U431 & P1_R2278_U430); 
assign P1_R2278_U102 = ~(P1_R2278_U438 & P1_R2278_U437); 
assign P1_R2278_U226 = ~(P1_R2278_U224 & P1_R2278_U139); 
assign P1_R2278_U275 = ~P1_R2278_U225; 
assign P1_R2278_U280 = ~P1_R2278_U224; 
assign P1_R2278_U328 = ~(P1_R2278_U281 & P1_R2278_U224); 
assign P1_R2278_U341 = ~(P1_R2278_U340 & P1_R2278_U225); 
assign P1_R2278_U344 = ~(P1_R2278_U278 & P1_R2278_U343); 
assign P1_R2278_U600 = ~(P1_R2278_U350 & P1_R2278_U224); 
assign P1_R2278_U607 = ~(P1_R2278_U351 & P1_R2278_U225); 
assign P1_R2358_U8 = P1_R2358_U288 & P1_R2358_U286; 
assign P1_R2358_U189 = ~(P1_R2358_U131 & P1_R2358_U385); 
assign P1_R2358_U190 = ~(P1_R2358_U365 & P1_R2358_U387); 
assign P1_R2358_U191 = ~(P1_R2358_U138 & P1_R2358_U389); 
assign P1_R2358_U192 = ~(P1_R2358_U391 & P1_R2358_U47); 
assign P1_R2358_U289 = ~(P1_U2626 & P1_R2358_U543); 
assign P1_R2358_U315 = ~(P1_R2358_U139 & P1_R2358_U314); 
assign P1_R2358_U320 = ~(P1_R2358_U313 & P1_R2358_U61); 
assign P1_R2358_U367 = ~(P1_R2358_U287 & P1_R2358_U288); 
assign P1_R2358_U526 = ~(P1_U2352 & P1_R2358_U172); 
assign P1_R2358_U538 = ~(P1_U2352 & P1_R2358_U172); 
assign P1_R2358_U599 = ~(P1_R2358_U108 & P1_R2358_U394); 
assign P1_R2358_U601 = ~(P1_R2358_U110 & P1_R2358_U396); 
assign P1_R2358_U603 = ~(P1_R2358_U112 & P1_R2358_U398); 
assign P1_R2099_U24 = ~(P1_R2099_U178 & P1_R2099_U46); 
assign P1_R2099_U302 = ~(P1_R2099_U231 & P1_R2099_U178); 
assign P1_R2337_U58 = ~(P1_R2337_U119 & P1_PHYADDRPOINTER_REG_28__SCAN_IN); 
assign P1_R2337_U146 = ~(P1_R2337_U119 & P1_R2337_U57); 
assign P1_R2096_U58 = ~(P1_R2096_U119 & P1_REIP_REG_28__SCAN_IN); 
assign P1_R2096_U146 = ~(P1_R2096_U119 & P1_R2096_U57); 
assign P1_ADD_405_U58 = ~(P1_ADD_405_U122 & P1_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P1_ADD_405_U176 = ~(P1_ADD_405_U122 & P1_ADD_405_U57); 
assign P1_ADD_515_U58 = ~(P1_ADD_515_U119 & P1_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P1_ADD_515_U172 = ~(P1_ADD_515_U119 & P1_ADD_515_U57); 
assign P3_U2838 = ~(P3_U3883 & P3_U6230); 
assign P3_U3895 = P3_U6260 & P3_U6259; 
assign P3_U3897 = P3_U6262 & P3_U6261 & P3_U6263 & P3_U3896; 
assign P3_U3900 = P3_U6272 & P3_U6271 & P3_U6273; 
assign P3_U3901 = P3_U6275 & P3_U6274; 
assign P3_U3905 = P3_U6289 & P3_U6288; 
assign P3_U3907 = P3_U6291 & P3_U6290 & P3_U6292; 
assign P3_U3908 = P3_U6294 & P3_U6293; 
assign P3_U3912 = P3_U6305 & P3_U6304; 
assign P3_U3981 = P3_U6628 & P3_U6627 & P3_U6626 & P3_U6625; 
assign P3_U4120 = P3_U7326 & P3_U7325; 
assign P3_U6252 = ~(P3_U3892 & P3_U3887); 
assign P3_U6328 = ~(P3_ADD_360_1242_U16 & P3_U2395); 
assign P3_U6639 = ~(P3_U2396 & P3_ADD_360_1242_U16); 
assign P2_U2794 = P2_U3242 & P2_R2267_U14; 
assign P2_U3662 = ~(P2_U8380 & P2_U8379); 
assign P2_U6459 = ~(P2_U2380 & P2_R2096_U78); 
assign P2_U6523 = ~(P2_U2379 & P2_R2099_U86); 
assign P2_U6537 = ~(P2_R2182_U84 & P2_U2393); 
assign P2_U6718 = ~(P2_U2392 & P2_R2099_U86); 
assign P2_U6795 = ~(P2_R2267_U14 & P2_U2587); 
assign P2_U6812 = ~(P2_U2588 & P2_R2096_U78); 
assign P1_U2856 = ~(P1_U6314 & P1_U6315 & P1_U6313); 
assign P1_U2888 = ~(P1_U6203 & P1_U6202 & P1_U6205 & P1_U6204); 
assign P1_U2992 = ~(P1_U5836 & P1_U5834 & P1_U5835 & P1_U5838 & P1_U5837); 
assign P1_U3024 = ~(P1_U3787 & P1_U3789 & P1_U5621); 
assign P1_U3847 = P1_U5760 & P1_U5762; 
assign P1_U3849 = P1_U3848 & P1_U5763; 
assign P1_U3940 = P1_U6566 & P1_U6564; 
assign P1_U4013 = P1_U6789 & P1_U6790 & P1_U6791; 
assign P1_U5628 = ~(P1_R2278_U102 & P1_U2377); 
assign P1_U5635 = ~(P1_R2278_U101 & P1_U2377); 
assign P1_U5840 = ~(P1_U2372 & P1_R2278_U102); 
assign P1_U5845 = ~(P1_U2372 & P1_R2278_U101); 
assign P3_ADD_476_U73 = ~(P3_ADD_476_U146 & P3_ADD_476_U145); 
assign P3_ADD_476_U120 = ~P3_ADD_476_U58; 
assign P3_ADD_476_U143 = ~(P3_ADD_476_U58 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_531_U77 = ~(P3_ADD_531_U153 & P3_ADD_531_U152); 
assign P3_ADD_531_U124 = ~P3_ADD_531_U59; 
assign P3_ADD_531_U150 = ~(P3_ADD_531_U59 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_SUB_320_U107 = ~(P3_SUB_320_U101 & P3_SUB_320_U63); 
assign P3_SUB_320_U141 = ~(P3_SUB_320_U101 & P3_SUB_320_U63); 
assign P3_ADD_318_U73 = ~(P3_ADD_318_U146 & P3_ADD_318_U145); 
assign P3_ADD_318_U120 = ~P3_ADD_318_U58; 
assign P3_ADD_318_U143 = ~(P3_ADD_318_U58 & P3_PHYADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_315_U69 = ~(P3_ADD_315_U138 & P3_ADD_315_U137); 
assign P3_ADD_315_U117 = ~P3_ADD_315_U58; 
assign P3_ADD_315_U135 = ~(P3_ADD_315_U58 & P3_PHYADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_360_1242_U187 = ~(P3_ADD_360_1242_U165 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_360_1242_U228 = ~(P3_ADD_360_1242_U165 & P3_ADD_360_1242_U116 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_360_1242_U230 = ~(P3_ADD_360_1242_U165 & P3_ADD_360_1242_U74); 
assign P3_ADD_467_U73 = ~(P3_ADD_467_U146 & P3_ADD_467_U145); 
assign P3_ADD_467_U120 = ~P3_ADD_467_U58; 
assign P3_ADD_467_U143 = ~(P3_ADD_467_U58 & P3_REIP_REG_29__SCAN_IN); 
assign P3_ADD_430_U73 = ~(P3_ADD_430_U146 & P3_ADD_430_U145); 
assign P3_ADD_430_U120 = ~P3_ADD_430_U58; 
assign P3_ADD_430_U143 = ~(P3_ADD_430_U58 & P3_REIP_REG_29__SCAN_IN); 
assign P3_ADD_380_U77 = ~(P3_ADD_380_U153 & P3_ADD_380_U152); 
assign P3_ADD_380_U124 = ~P3_ADD_380_U59; 
assign P3_ADD_380_U150 = ~(P3_ADD_380_U59 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_344_U77 = ~(P3_ADD_344_U153 & P3_ADD_344_U152); 
assign P3_ADD_344_U124 = ~P3_ADD_344_U59; 
assign P3_ADD_344_U150 = ~(P3_ADD_344_U59 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_339_U73 = ~(P3_ADD_339_U146 & P3_ADD_339_U145); 
assign P3_ADD_339_U120 = ~P3_ADD_339_U58; 
assign P3_ADD_339_U143 = ~(P3_ADD_339_U58 & P3_PHYADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_541_U73 = ~(P3_ADD_541_U146 & P3_ADD_541_U145); 
assign P3_ADD_541_U120 = ~P3_ADD_541_U58; 
assign P3_ADD_541_U143 = ~(P3_ADD_541_U58 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_515_U73 = ~(P3_ADD_515_U146 & P3_ADD_515_U145); 
assign P3_ADD_515_U120 = ~P3_ADD_515_U58; 
assign P3_ADD_515_U143 = ~(P3_ADD_515_U58 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_394_U72 = ~(P3_ADD_394_U148 & P3_ADD_394_U147); 
assign P3_ADD_394_U123 = ~P3_ADD_394_U58; 
assign P3_ADD_394_U145 = ~(P3_ADD_394_U58 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_441_U73 = ~(P3_ADD_441_U146 & P3_ADD_441_U145); 
assign P3_ADD_441_U120 = ~P3_ADD_441_U58; 
assign P3_ADD_441_U143 = ~(P3_ADD_441_U58 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_349_U77 = ~(P3_ADD_349_U153 & P3_ADD_349_U152); 
assign P3_ADD_349_U124 = ~P3_ADD_349_U59; 
assign P3_ADD_349_U150 = ~(P3_ADD_349_U59 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_405_U72 = ~(P3_ADD_405_U148 & P3_ADD_405_U147); 
assign P3_ADD_405_U123 = ~P3_ADD_405_U58; 
assign P3_ADD_405_U145 = ~(P3_ADD_405_U58 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_553_U77 = ~(P3_ADD_553_U153 & P3_ADD_553_U152); 
assign P3_ADD_553_U124 = ~P3_ADD_553_U59; 
assign P3_ADD_553_U150 = ~(P3_ADD_553_U59 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_558_U77 = ~(P3_ADD_558_U153 & P3_ADD_558_U152); 
assign P3_ADD_558_U124 = ~P3_ADD_558_U59; 
assign P3_ADD_558_U150 = ~(P3_ADD_558_U59 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_385_U77 = ~(P3_ADD_385_U153 & P3_ADD_385_U152); 
assign P3_ADD_385_U124 = ~P3_ADD_385_U59; 
assign P3_ADD_385_U150 = ~(P3_ADD_385_U59 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_547_U77 = ~(P3_ADD_547_U153 & P3_ADD_547_U152); 
assign P3_ADD_547_U124 = ~P3_ADD_547_U59; 
assign P3_ADD_547_U150 = ~(P3_ADD_547_U59 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_371_1212_U79 = ~(P3_ADD_371_1212_U239 & P3_ADD_371_1212_U238); 
assign P3_ADD_371_1212_U236 = ~(P3_ADD_371_1212_U198 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_494_U73 = ~(P3_ADD_494_U146 & P3_ADD_494_U145); 
assign P3_ADD_494_U120 = ~P3_ADD_494_U58; 
assign P3_ADD_494_U143 = ~(P3_ADD_494_U58 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_536_U73 = ~(P3_ADD_536_U146 & P3_ADD_536_U145); 
assign P3_ADD_536_U120 = ~P3_ADD_536_U58; 
assign P3_ADD_536_U143 = ~(P3_ADD_536_U58 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P2_R2099_U43 = ~(P2_U2729 & P2_R2099_U133); 
assign P2_R2099_U207 = ~(P2_R2099_U133 & P2_R2099_U42); 
assign P2_ADD_391_1196_U5 = P2_ADD_391_1196_U301 & P2_ADD_391_1196_U299; 
assign P2_ADD_391_1196_U66 = ~P2_R2182_U84; 
assign P2_ADD_391_1196_U80 = ~P2_R2096_U78; 
assign P2_ADD_391_1196_U84 = ~(P2_ADD_391_1196_U216 & P2_ADD_391_1196_U215); 
assign P2_ADD_391_1196_U141 = P2_ADD_391_1196_U415 & P2_ADD_391_1196_U414; 
assign P2_ADD_391_1196_U252 = P2_R2182_U84 | P2_R2096_U85; 
assign P2_ADD_391_1196_U254 = ~(P2_R2096_U85 & P2_R2182_U84); 
assign P2_ADD_391_1196_U401 = ~(P2_R2182_U84 & P2_ADD_391_1196_U67); 
assign P2_ADD_391_1196_U403 = ~(P2_R2182_U84 & P2_ADD_391_1196_U67); 
assign P2_ADD_391_1196_U407 = ~(P2_R2096_U86 & P2_ADD_391_1196_U64); 
assign P2_ADD_391_1196_U409 = ~(P2_R2096_U86 & P2_ADD_391_1196_U64); 
assign P2_ADD_391_1196_U418 = ~(P2_ADD_391_1196_U417 & P2_ADD_391_1196_U416); 
assign P2_ADD_391_1196_U469 = ~(P2_ADD_391_1196_U213 & P2_ADD_391_1196_U467); 
assign P2_R2182_U83 = ~(P2_R2182_U272 & P2_R2182_U271); 
assign P2_R2182_U158 = ~P2_R2182_U119; 
assign P2_R2182_U160 = ~(P2_R2182_U159 & P2_R2182_U119); 
assign P2_R2182_U264 = ~(P2_R2182_U118 & P2_R2182_U119); 
assign P2_R2027_U77 = ~(P2_R2027_U153 & P2_R2027_U152); 
assign P2_R2027_U124 = ~P2_R2027_U59; 
assign P2_R2027_U150 = ~(P2_R2027_U59 & P2_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P2_R2337_U71 = ~(P2_R2337_U144 & P2_R2337_U143); 
assign P2_R2337_U121 = ~P2_R2337_U59; 
assign P2_R2337_U139 = ~(P2_R2337_U59 & P2_PHYADDRPOINTER_REG_30__SCAN_IN); 
assign P2_R2096_U50 = P2_R2096_U168 & P2_R2096_U167; 
assign P2_R2096_U76 = ~(P2_R2096_U211 & P2_R2096_U210); 
assign P2_R1957_U107 = ~(P2_R1957_U101 & P2_R1957_U63); 
assign P2_R1957_U141 = ~(P2_R1957_U101 & P2_R1957_U63); 
assign P2_R2278_U7 = ~P2_U3631; 
assign P2_R2278_U76 = ~P2_U2795; 
assign P2_R2278_U78 = ~(P2_U2795 & P2_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P2_R2278_U120 = P2_R2278_U320 & P2_R2278_U236; 
assign P2_R2278_U135 = P2_R2278_U338 & P2_R2278_U288; 
assign P2_R2278_U151 = P2_R2278_U368 & P2_R2278_U367; 
assign P2_R2278_U175 = P2_R2278_U452 & P2_R2278_U451; 
assign P2_R2278_U223 = ~P2_R2278_U152; 
assign P2_R2278_U225 = ~(P2_R2278_U224 & P2_R2278_U152); 
assign P2_R2278_U228 = P2_U3631 | P2_INSTADDRPOINTER_REG_7__SCAN_IN; 
assign P2_R2278_U229 = ~(P2_U3631 & P2_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P2_R2278_U292 = P2_U2795 | P2_INSTADDRPOINTER_REG_26__SCAN_IN; 
assign P2_R2278_U361 = ~(P2_U3631 & P2_R2278_U8); 
assign P2_R2278_U363 = ~(P2_U3631 & P2_R2278_U8); 
assign P2_R2278_U371 = ~(P2_R2278_U370 & P2_R2278_U369); 
assign P2_R2278_U380 = ~(P2_R2278_U220 & P2_R2278_U378); 
assign P2_R2278_U438 = ~(P2_U2795 & P2_R2278_U77); 
assign P2_R2278_U440 = ~(P2_U2795 & P2_R2278_U77); 
assign P2_R2278_U455 = ~(P2_R2278_U454 & P2_R2278_U453); 
assign P2_ADD_394_U86 = ~(P2_ADD_394_U176 & P2_ADD_394_U175); 
assign P2_ADD_394_U123 = ~P2_ADD_394_U58; 
assign P2_ADD_394_U131 = ~(P2_ADD_394_U58 & P2_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P2_R2267_U67 = P2_R2267_U146 & P2_R2267_U145; 
assign P2_R2267_U111 = ~P2_R2267_U40; 
assign P2_R2267_U113 = ~(P2_U2767 & P2_R2267_U40); 
assign P2_R2267_U115 = ~(P2_U2768 & P2_R2267_U114); 
assign P2_ADD_371_1212_U81 = ~(P2_ADD_371_1212_U248 & P2_ADD_371_1212_U247); 
assign P2_ADD_371_1212_U133 = P2_ADD_371_1212_U275 & P2_ADD_371_1212_U274; 
assign P2_ADD_371_1212_U156 = ~P2_ADD_371_1212_U111; 
assign P2_ADD_371_1212_U158 = ~(P2_ADD_371_1212_U157 & P2_ADD_371_1212_U111); 
assign P2_ADD_371_1212_U212 = ~(P2_ADD_371_1212_U110 & P2_ADD_371_1212_U111); 
assign P2_ADD_371_1212_U278 = ~(P2_ADD_371_1212_U277 & P2_ADD_371_1212_U276); 
assign P1_R2278_U222 = ~(P1_R2278_U168 & P1_R2278_U226); 
assign P1_R2278_U223 = ~(P1_R2278_U68 & P1_R2278_U328); 
assign P1_R2278_U342 = ~(P1_R2278_U175 & P1_R2278_U341); 
assign P1_R2278_U411 = ~(P1_R2278_U141 & P1_R2278_U226); 
assign P1_R2278_U413 = ~(P1_R2278_U151 & P1_R2278_U226); 
assign P1_R2278_U418 = ~(P1_R2278_U160 & P1_R2278_U226); 
assign P1_R2278_U601 = ~(P1_R2278_U124 & P1_R2278_U280); 
assign P1_R2278_U608 = ~(P1_R2278_U275 & P1_R2278_U606); 
assign P1_R2358_U16 = P1_R2358_U320 & P1_R2358_U319; 
assign P1_R2358_U17 = P1_R2358_U317 & P1_R2358_U315; 
assign P1_R2358_U96 = P1_R2358_U289 & P1_R2358_U288; 
assign P1_R2358_U109 = ~(P1_R2358_U599 & P1_R2358_U598); 
assign P1_R2358_U111 = ~(P1_R2358_U601 & P1_R2358_U600); 
assign P1_R2358_U113 = ~(P1_R2358_U603 & P1_R2358_U602); 
assign P1_R2358_U137 = P1_R2358_U367 & P1_R2358_U289; 
assign P1_R2358_U171 = ~P1_U2656; 
assign P1_R2358_U290 = ~(P1_R2358_U527 & P1_R2358_U526 & P1_R2358_U39); 
assign P1_R2358_U341 = ~(P1_R2358_U289 & P1_R2358_U288); 
assign P1_R2358_U368 = ~(P1_R2358_U367 & P1_R2358_U289); 
assign P1_R2358_U375 = ~(P1_R2358_U286 & P1_R2358_U189); 
assign P1_R2358_U377 = ~(P1_R2358_U8 & P1_R2358_U189); 
assign P1_R2358_U386 = ~P1_R2358_U189; 
assign P1_R2358_U388 = ~P1_R2358_U190; 
assign P1_R2358_U390 = ~P1_R2358_U191; 
assign P1_R2358_U392 = ~P1_R2358_U192; 
assign P1_R2358_U525 = ~(P1_U2656 & P1_R2358_U23); 
assign P1_R2358_U536 = ~(P1_U2656 & P1_R2358_U23); 
assign P1_R2358_U540 = ~(P1_R2358_U539 & P1_R2358_U538); 
assign P1_R2358_U588 = ~(P1_R2358_U189 & P1_R2358_U342); 
assign P1_R2358_U590 = ~(P1_R2358_U190 & P1_R2358_U343); 
assign P1_R2358_U592 = ~(P1_R2358_U191 & P1_R2358_U344); 
assign P1_R2358_U594 = ~(P1_R2358_U192 & P1_R2358_U345); 
assign P1_R2099_U68 = ~(P1_R2099_U303 & P1_R2099_U302); 
assign P1_R2099_U179 = ~P1_R2099_U24; 
assign P1_R2099_U301 = ~(P1_R2099_U45 & P1_R2099_U24); 
assign P1_R2337_U73 = ~(P1_R2337_U146 & P1_R2337_U145); 
assign P1_R2337_U120 = ~P1_R2337_U58; 
assign P1_R2337_U143 = ~(P1_R2337_U58 & P1_PHYADDRPOINTER_REG_29__SCAN_IN); 
assign P1_R2096_U73 = ~(P1_R2096_U146 & P1_R2096_U145); 
assign P1_R2096_U120 = ~P1_R2096_U58; 
assign P1_R2096_U143 = ~(P1_R2096_U58 & P1_REIP_REG_29__SCAN_IN); 
assign P1_ADD_405_U86 = ~(P1_ADD_405_U176 & P1_ADD_405_U175); 
assign P1_ADD_405_U123 = ~P1_ADD_405_U58; 
assign P1_ADD_405_U131 = ~(P1_ADD_405_U58 & P1_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P1_ADD_515_U86 = ~(P1_ADD_515_U172 & P1_ADD_515_U171); 
assign P1_ADD_515_U120 = ~P1_ADD_515_U58; 
assign P1_ADD_515_U127 = ~(P1_ADD_515_U58 & P1_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_U2803 = ~(P3_U6622 & P3_U6624 & P3_U6621 & P3_U6623 & P3_U3981); 
assign P3_U3902 = P3_U3899 & P3_U3898 & P3_U3901 & P3_U3900; 
assign P3_U3921 = P3_U6329 & P3_U6328; 
assign P3_U6254 = ~(P3_U4318 & P3_U6252); 
assign P3_U6282 = ~(P3_ADD_558_U77 & P3_U3220); 
assign P3_U6283 = ~(P3_ADD_553_U77 & P3_U4298); 
assign P3_U6284 = ~(P3_ADD_547_U77 & P3_U4299); 
assign P3_U6287 = ~(P3_ADD_531_U77 & P3_U2354); 
assign P3_U6295 = ~(P3_ADD_385_U77 & P3_U2358); 
assign P3_U6296 = ~(P3_ADD_380_U77 & P3_U2359); 
assign P3_U6297 = ~(P3_ADD_349_U77 & P3_U4306); 
assign P3_U6298 = ~(P3_ADD_344_U77 & P3_U2362); 
assign P3_U6309 = ~(P3_ADD_541_U73 & P3_U4300); 
assign P3_U6310 = ~(P3_ADD_536_U73 & P3_U4301); 
assign P3_U6313 = ~(P3_ADD_515_U73 & P3_U4302); 
assign P3_U6314 = ~(P3_ADD_494_U73 & P3_U2356); 
assign P3_U6315 = ~(P3_ADD_476_U73 & P3_U4303); 
assign P3_U6316 = ~(P3_ADD_441_U73 & P3_U4304); 
assign P3_U6317 = ~(P3_ADD_405_U72 & P3_U4305); 
assign P3_U6318 = ~(P3_ADD_394_U72 & P3_U2357); 
assign P3_U6371 = ~(P3_ADD_371_1212_U79 & P3_U2360); 
assign P3_U6629 = ~(P3_ADD_318_U73 & P3_U2398); 
assign P3_U6634 = ~(P3_ADD_339_U73 & P3_U2388); 
assign P3_U6638 = ~(P3_ADD_315_U69 & P3_U2397); 
assign P3_U6651 = ~(P3_U2387 & P3_ADD_371_1212_U79); 
assign P3_U7334 = ~(P3_ADD_467_U73 & P3_U2601); 
assign P3_U7336 = ~(P3_ADD_430_U73 & P3_U2405); 
assign P2_U2793 = P2_U3242 & P2_R2267_U67; 
assign P2_U2870 = ~(P2_U6523 & P2_U6524 & P2_U6522); 
assign P2_U6372 = ~(P2_ADD_391_1196_U5 & P2_U2397); 
assign P2_U6464 = ~(P2_U2380 & P2_R2096_U76); 
assign P2_U6467 = ~(P2_U2380 & P2_R2096_U50); 
assign P2_U6540 = ~(P2_R2182_U83 & P2_U2393); 
assign P2_U6803 = ~(P2_R2267_U67 & P2_U2587); 
assign P2_U6820 = ~(P2_U2588 & P2_R2096_U76); 
assign P2_U6828 = ~(P2_U2588 & P2_R2096_U50); 
assign P2_U8377 = ~(P2_R2337_U71 & P2_U3284); 
assign P1_U2655 = ~(P1_U6788 & P1_U4013); 
assign P1_U2990 = ~(P1_U5846 & P1_U5844 & P1_U5848 & P1_U5845 & P1_U5847); 
assign P1_U2991 = ~(P1_U5841 & P1_U5839 & P1_U5843 & P1_U5840 & P1_U5842); 
assign P1_U3022 = ~(P1_U3793 & P1_U3795 & P1_U5635); 
assign P1_U3023 = ~(P1_U3790 & P1_U3792 & P1_U5628); 
assign P1_U5759 = ~(P1_R2099_U68 & P1_U2380); 
assign P1_U5769 = ~(P1_ADD_405_U86 & P1_U2375); 
assign P1_U5770 = ~(P1_ADD_515_U86 & P1_U2374); 
assign P1_U5872 = ~(P1_R2358_U16 & P1_U2364); 
assign P1_U5877 = ~(P1_R2358_U17 & P1_U2364); 
assign P1_U5887 = ~(P1_R2358_U113 & P1_U2364); 
assign P1_U5892 = ~(P1_R2358_U111 & P1_U2364); 
assign P1_U5897 = ~(P1_R2358_U109 & P1_U2364); 
assign P1_U5939 = ~(P1_R2337_U73 & P1_U2376); 
assign P1_U6197 = ~(P1_U2386 & P1_R2358_U16); 
assign P1_U6200 = ~(P1_U2386 & P1_R2358_U17); 
assign P1_U6208 = ~(P1_U2386 & P1_R2358_U113); 
assign P1_U6212 = ~(P1_U2386 & P1_R2358_U111); 
assign P1_U6216 = ~(P1_U2386 & P1_R2358_U109); 
assign P1_U6307 = ~(P1_U2383 & P1_R2358_U16); 
assign P1_U6310 = ~(P1_U2383 & P1_R2358_U17); 
assign P1_U6316 = ~(P1_U2383 & P1_R2358_U113); 
assign P1_U6319 = ~(P1_U2383 & P1_R2358_U111); 
assign P1_U6322 = ~(P1_U2383 & P1_R2358_U109); 
assign P1_U6347 = ~(P1_U2371 & P1_R2099_U68); 
assign P1_U6563 = ~(P1_U2604 & P1_R2099_U68); 
assign P1_U6571 = ~(P1_R2096_U73 & P1_U7485); 
assign P1_U6787 = ~(P1_R2337_U73 & P1_U2352); 
assign P3_ADD_476_U60 = ~(P3_ADD_476_U120 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_476_U144 = ~(P3_ADD_476_U120 & P3_ADD_476_U59); 
assign P3_ADD_531_U61 = ~(P3_ADD_531_U124 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_531_U151 = ~(P3_ADD_531_U124 & P3_ADD_531_U60); 
assign P3_SUB_320_U40 = ~P3_ADD_318_U73; 
assign P3_SUB_320_U64 = P3_SUB_320_U141 & P3_SUB_320_U140; 
assign P3_SUB_320_U108 = ~(P3_ADD_318_U73 & P3_SUB_320_U107); 
assign P3_ADD_318_U60 = ~(P3_ADD_318_U120 & P3_PHYADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_318_U144 = ~(P3_ADD_318_U120 & P3_ADD_318_U59); 
assign P3_ADD_315_U90 = ~(P3_ADD_315_U117 & P3_PHYADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_315_U136 = ~(P3_ADD_315_U117 & P3_ADD_315_U59); 
assign P3_ADD_360_1242_U77 = ~(P3_ADD_360_1242_U230 & P3_ADD_360_1242_U229); 
assign P3_ADD_360_1242_U227 = ~(P3_ADD_360_1242_U187 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_467_U60 = ~(P3_ADD_467_U120 & P3_REIP_REG_29__SCAN_IN); 
assign P3_ADD_467_U144 = ~(P3_ADD_467_U120 & P3_ADD_467_U59); 
assign P3_ADD_430_U60 = ~(P3_ADD_430_U120 & P3_REIP_REG_29__SCAN_IN); 
assign P3_ADD_430_U144 = ~(P3_ADD_430_U120 & P3_ADD_430_U59); 
assign P3_ADD_380_U61 = ~(P3_ADD_380_U124 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_380_U151 = ~(P3_ADD_380_U124 & P3_ADD_380_U60); 
assign P3_ADD_344_U61 = ~(P3_ADD_344_U124 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_344_U151 = ~(P3_ADD_344_U124 & P3_ADD_344_U60); 
assign P3_ADD_339_U60 = ~(P3_ADD_339_U120 & P3_PHYADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_339_U144 = ~(P3_ADD_339_U120 & P3_ADD_339_U59); 
assign P3_ADD_541_U60 = ~(P3_ADD_541_U120 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_541_U144 = ~(P3_ADD_541_U120 & P3_ADD_541_U59); 
assign P3_ADD_515_U60 = ~(P3_ADD_515_U120 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_515_U144 = ~(P3_ADD_515_U120 & P3_ADD_515_U59); 
assign P3_ADD_394_U60 = ~(P3_ADD_394_U123 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_394_U146 = ~(P3_ADD_394_U123 & P3_ADD_394_U59); 
assign P3_ADD_441_U60 = ~(P3_ADD_441_U120 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_441_U144 = ~(P3_ADD_441_U120 & P3_ADD_441_U59); 
assign P3_ADD_349_U61 = ~(P3_ADD_349_U124 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_349_U151 = ~(P3_ADD_349_U124 & P3_ADD_349_U60); 
assign P3_ADD_405_U60 = ~(P3_ADD_405_U123 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_405_U146 = ~(P3_ADD_405_U123 & P3_ADD_405_U59); 
assign P3_ADD_553_U61 = ~(P3_ADD_553_U124 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_553_U151 = ~(P3_ADD_553_U124 & P3_ADD_553_U60); 
assign P3_ADD_558_U61 = ~(P3_ADD_558_U124 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_558_U151 = ~(P3_ADD_558_U124 & P3_ADD_558_U60); 
assign P3_ADD_385_U61 = ~(P3_ADD_385_U124 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_385_U151 = ~(P3_ADD_385_U124 & P3_ADD_385_U60); 
assign P3_ADD_547_U61 = ~(P3_ADD_547_U124 & P3_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P3_ADD_547_U151 = ~(P3_ADD_547_U124 & P3_ADD_547_U60); 
assign P3_ADD_371_1212_U92 = ~(P3_ADD_371_1212_U237 & P3_ADD_371_1212_U236); 
assign P3_ADD_494_U60 = ~(P3_ADD_494_U120 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_494_U144 = ~(P3_ADD_494_U120 & P3_ADD_494_U59); 
assign P3_ADD_536_U60 = ~(P3_ADD_536_U120 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_536_U144 = ~(P3_ADD_536_U120 & P3_ADD_536_U59); 
assign P2_R2099_U85 = ~(P2_R2099_U207 & P2_R2099_U206); 
assign P2_R2099_U134 = ~P2_R2099_U43; 
assign P2_R2099_U204 = ~(P2_U2728 & P2_R2099_U43); 
assign P2_ADD_391_1196_U68 = ~P2_R2182_U83; 
assign P2_ADD_391_1196_U85 = ~(P2_ADD_391_1196_U84 & P2_ADD_391_1196_U218); 
assign P2_ADD_391_1196_U108 = ~(P2_ADD_391_1196_U469 & P2_ADD_391_1196_U468); 
assign P2_ADD_391_1196_U120 = ~P2_R2096_U76; 
assign P2_ADD_391_1196_U139 = P2_ADD_391_1196_U408 & P2_ADD_391_1196_U407; 
assign P2_ADD_391_1196_U217 = ~P2_ADD_391_1196_U84; 
assign P2_ADD_391_1196_U256 = P2_R2182_U83 | P2_R2096_U84; 
assign P2_ADD_391_1196_U258 = ~(P2_R2096_U84 & P2_R2182_U83); 
assign P2_ADD_391_1196_U394 = ~(P2_R2182_U83 & P2_ADD_391_1196_U69); 
assign P2_ADD_391_1196_U396 = ~(P2_R2182_U83 & P2_ADD_391_1196_U69); 
assign P2_ADD_391_1196_U400 = ~(P2_R2096_U85 & P2_ADD_391_1196_U66); 
assign P2_ADD_391_1196_U402 = ~(P2_R2096_U85 & P2_ADD_391_1196_U66); 
assign P2_ADD_391_1196_U411 = ~(P2_ADD_391_1196_U410 & P2_ADD_391_1196_U409); 
assign P2_R2182_U117 = ~(P2_R2182_U161 & P2_R2182_U160); 
assign P2_R2182_U265 = ~(P2_R2182_U158 & P2_R2182_U263); 
assign P2_R2027_U61 = ~(P2_R2027_U124 & P2_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P2_R2027_U151 = ~(P2_R2027_U124 & P2_R2027_U60); 
assign P2_R2337_U93 = ~(P2_R2337_U121 & P2_PHYADDRPOINTER_REG_30__SCAN_IN); 
assign P2_R2337_U140 = ~(P2_R2337_U121 & P2_R2337_U60); 
assign P2_R1957_U39 = ~P2_U3662; 
assign P2_R1957_U64 = P2_R1957_U141 & P2_R1957_U140; 
assign P2_R1957_U108 = ~(P2_U3662 & P2_R1957_U107); 
assign P2_R2278_U74 = ~P2_U2794; 
assign P2_R2278_U88 = ~(P2_R2278_U380 & P2_R2278_U379); 
assign P2_R2278_U117 = P2_R2278_U224 & P2_R2278_U228; 
assign P2_R2278_U150 = ~(P2_R2278_U26 & P2_R2278_U225); 
assign P2_R2278_U294 = ~P2_R2278_U78; 
assign P2_R2278_U296 = P2_U2794 | P2_INSTADDRPOINTER_REG_27__SCAN_IN; 
assign P2_R2278_U297 = ~(P2_U2794 & P2_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P2_R2278_U318 = ~(P2_R2278_U226 & P2_R2278_U228); 
assign P2_R2278_U360 = ~(P2_R2278_U7 & P2_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P2_R2278_U362 = ~(P2_R2278_U7 & P2_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P2_R2278_U372 = ~(P2_R2278_U151 & P2_R2278_U152); 
assign P2_R2278_U373 = ~(P2_R2278_U223 & P2_R2278_U371); 
assign P2_R2278_U431 = ~(P2_U2794 & P2_R2278_U75); 
assign P2_R2278_U433 = ~(P2_U2794 & P2_R2278_U75); 
assign P2_R2278_U437 = ~(P2_R2278_U76 & P2_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P2_R2278_U439 = ~(P2_R2278_U76 & P2_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P2_ADD_394_U61 = ~(P2_ADD_394_U123 & P2_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P2_ADD_394_U132 = ~(P2_ADD_394_U123 & P2_ADD_394_U59); 
assign P2_R2267_U15 = P2_R2267_U115 & P2_R2267_U40; 
assign P2_R2267_U62 = ~(P2_R2267_U111 & P2_R2267_U41); 
assign P2_ADD_371_1212_U134 = ~(P2_ADD_371_1212_U159 & P2_ADD_371_1212_U158); 
assign P2_ADD_371_1212_U213 = ~(P2_ADD_371_1212_U156 & P2_ADD_371_1212_U211); 
assign P1_R2278_U15 = P1_R2278_U344 & P1_R2278_U342; 
assign P1_R2278_U125 = ~(P1_R2278_U601 & P1_R2278_U600); 
assign P1_R2278_U126 = ~(P1_R2278_U608 & P1_R2278_U607); 
assign P1_R2278_U289 = ~(P1_R2278_U288 & P1_R2278_U222); 
assign P1_R2278_U329 = ~P1_R2278_U223; 
assign P1_R2278_U331 = ~(P1_R2278_U330 & P1_R2278_U223); 
assign P1_R2278_U358 = ~(P1_R2278_U6 & P1_R2278_U222); 
assign P1_R2278_U361 = ~(P1_R2278_U7 & P1_R2278_U222); 
assign P1_R2278_U376 = ~(P1_R2278_U161 & P1_R2278_U418); 
assign P1_R2278_U385 = ~(P1_R2278_U11 & P1_R2278_U411 & P1_R2278_U142); 
assign P1_R2278_U397 = ~(P1_R2278_U152 & P1_R2278_U413 & P1_R2278_U153); 
assign P1_R2278_U405 = ~(P1_R2278_U157 & P1_R2278_U411 & P1_R2278_U158); 
assign P1_R2278_U416 = ~P1_R2278_U222; 
assign P1_R2278_U586 = ~(P1_R2278_U221 & P1_R2278_U222); 
assign P1_R2278_U598 = ~(P1_R2278_U349 & P1_R2278_U223); 
assign P1_R2358_U9 = P1_R2358_U8 & P1_R2358_U290; 
assign P1_R2358_U187 = ~(P1_R2358_U137 & P1_R2358_U377); 
assign P1_R2358_U188 = ~(P1_R2358_U375 & P1_R2358_U42); 
assign P1_R2358_U291 = ~(P1_U2625 & P1_R2358_U540); 
assign P1_R2358_U369 = ~(P1_R2358_U368 & P1_R2358_U290); 
assign P1_R2358_U524 = ~(P1_U2352 & P1_R2358_U171); 
assign P1_R2358_U535 = ~(P1_U2352 & P1_R2358_U171); 
assign P1_R2358_U589 = ~(P1_R2358_U98 & P1_R2358_U386); 
assign P1_R2358_U591 = ~(P1_R2358_U100 & P1_R2358_U388); 
assign P1_R2358_U593 = ~(P1_R2358_U102 & P1_R2358_U390); 
assign P1_R2358_U595 = ~(P1_R2358_U104 & P1_R2358_U392); 
assign P1_R2099_U25 = ~(P1_R2099_U179 & P1_R2099_U45); 
assign P1_R2099_U300 = ~(P1_R2099_U228 & P1_R2099_U179); 
assign P1_R2337_U60 = ~(P1_R2337_U120 & P1_PHYADDRPOINTER_REG_29__SCAN_IN); 
assign P1_R2337_U144 = ~(P1_R2337_U120 & P1_R2337_U59); 
assign P1_R2096_U60 = ~(P1_R2096_U120 & P1_REIP_REG_29__SCAN_IN); 
assign P1_R2096_U144 = ~(P1_R2096_U120 & P1_R2096_U59); 
assign P1_ADD_405_U61 = ~(P1_ADD_405_U123 & P1_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P1_ADD_405_U132 = ~(P1_ADD_405_U123 & P1_ADD_405_U59); 
assign P1_ADD_515_U61 = ~(P1_ADD_515_U120 & P1_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P1_ADD_515_U128 = ~(P1_ADD_515_U120 & P1_ADD_515_U59); 
assign P3_U2837 = ~(P3_U3893 & P3_U6254); 
assign P3_U3904 = P3_U6284 & P3_U6283; 
assign P3_U3906 = P3_U6286 & P3_U6285 & P3_U6287 & P3_U3905; 
assign P3_U3909 = P3_U6296 & P3_U6295 & P3_U6297; 
assign P3_U3910 = P3_U6299 & P3_U6298; 
assign P3_U3914 = P3_U6313 & P3_U6312; 
assign P3_U3916 = P3_U6315 & P3_U6314 & P3_U6316; 
assign P3_U3917 = P3_U6318 & P3_U6317; 
assign P3_U3982 = P3_U6636 & P3_U6635 & P3_U6634 & P3_U6633; 
assign P3_U4123 = P3_U7334 & P3_U7333; 
assign P3_U6276 = ~(P3_U3894 & P3_U6258 & P3_U3895 & P3_U3897 & P3_U3902); 
assign P3_U6352 = ~(P3_ADD_360_1242_U77 & P3_U2395); 
assign P3_U6395 = ~(P3_ADD_371_1212_U92 & P3_U2360); 
assign P3_U6647 = ~(P3_U2396 & P3_ADD_360_1242_U77); 
assign P3_U6659 = ~(P3_U2387 & P3_ADD_371_1212_U92); 
assign P2_U2792 = P2_U3242 & P2_R2267_U15; 
assign P2_U2888 = ~(P2_U6468 & P2_U6466 & P2_U6467); 
assign P2_U2908 = ~(P2_U6374 & P2_U6371 & P2_U6373 & P2_U6372); 
assign P2_U3661 = ~(P2_U8378 & P2_U8377); 
assign P2_U6376 = ~(P2_ADD_391_1196_U108 & P2_U2397); 
assign P2_U6526 = ~(P2_U2379 & P2_R2099_U85); 
assign P2_U6726 = ~(P2_U2392 & P2_R2099_U85); 
assign P2_U6811 = ~(P2_R2267_U15 & P2_U2587); 
assign P1_U2853 = ~(P1_U6323 & P1_U6324 & P1_U6322); 
assign P1_U2854 = ~(P1_U6320 & P1_U6321 & P1_U6319); 
assign P1_U2855 = ~(P1_U6317 & P1_U6318 & P1_U6316); 
assign P1_U2857 = ~(P1_U6311 & P1_U6312 & P1_U6310); 
assign P1_U2858 = ~(P1_U6308 & P1_U6309 & P1_U6307); 
assign P1_U2885 = ~(P1_U6215 & P1_U6214 & P1_U6217 & P1_U6216); 
assign P1_U2886 = ~(P1_U6211 & P1_U6210 & P1_U6213 & P1_U6212); 
assign P1_U2887 = ~(P1_U6207 & P1_U6206 & P1_U6209 & P1_U6208); 
assign P1_U2889 = ~(P1_U6201 & P1_U6199 & P1_U6200); 
assign P1_U2890 = ~(P1_U6198 & P1_U6196 & P1_U6197); 
assign P1_U3850 = P1_U5767 & P1_U5769; 
assign P1_U3852 = P1_U3851 & P1_U5770; 
assign P1_U3942 = P1_U6573 & P1_U6571; 
assign P1_U4012 = P1_U6785 & P1_U6786 & P1_U6787; 
assign P1_U5642 = ~(P1_R2278_U126 & P1_U2377); 
assign P1_U5649 = ~(P1_R2278_U15 & P1_U2377); 
assign P1_U5656 = ~(P1_R2278_U125 & P1_U2377); 
assign P1_U5850 = ~(P1_U2372 & P1_R2278_U126); 
assign P1_U5855 = ~(P1_U2372 & P1_R2278_U15); 
assign P1_U5860 = ~(P1_U2372 & P1_R2278_U125); 
assign P3_ADD_476_U72 = ~(P3_ADD_476_U144 & P3_ADD_476_U143); 
assign P3_ADD_476_U121 = ~P3_ADD_476_U60; 
assign P3_ADD_476_U139 = ~(P3_ADD_476_U60 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_531_U76 = ~(P3_ADD_531_U151 & P3_ADD_531_U150); 
assign P3_ADD_531_U125 = ~P3_ADD_531_U61; 
assign P3_ADD_531_U148 = ~(P3_ADD_531_U61 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_SUB_320_U37 = ~(P3_SUB_320_U40 & P3_SUB_320_U63 & P3_SUB_320_U101); 
assign P3_ADD_318_U72 = ~(P3_ADD_318_U144 & P3_ADD_318_U143); 
assign P3_ADD_318_U121 = ~P3_ADD_318_U60; 
assign P3_ADD_318_U139 = ~(P3_ADD_318_U60 & P3_PHYADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_315_U68 = ~(P3_ADD_315_U136 & P3_ADD_315_U135); 
assign P3_ADD_315_U118 = ~P3_ADD_315_U90; 
assign P3_ADD_315_U133 = ~(P3_ADD_315_U90 & P3_PHYADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_360_1242_U90 = ~(P3_ADD_360_1242_U228 & P3_ADD_360_1242_U227); 
assign P3_ADD_467_U72 = ~(P3_ADD_467_U144 & P3_ADD_467_U143); 
assign P3_ADD_467_U121 = ~P3_ADD_467_U60; 
assign P3_ADD_467_U139 = ~(P3_ADD_467_U60 & P3_REIP_REG_30__SCAN_IN); 
assign P3_ADD_430_U72 = ~(P3_ADD_430_U144 & P3_ADD_430_U143); 
assign P3_ADD_430_U121 = ~P3_ADD_430_U60; 
assign P3_ADD_430_U139 = ~(P3_ADD_430_U60 & P3_REIP_REG_30__SCAN_IN); 
assign P3_ADD_380_U76 = ~(P3_ADD_380_U151 & P3_ADD_380_U150); 
assign P3_ADD_380_U125 = ~P3_ADD_380_U61; 
assign P3_ADD_380_U148 = ~(P3_ADD_380_U61 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_344_U76 = ~(P3_ADD_344_U151 & P3_ADD_344_U150); 
assign P3_ADD_344_U125 = ~P3_ADD_344_U61; 
assign P3_ADD_344_U148 = ~(P3_ADD_344_U61 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_339_U72 = ~(P3_ADD_339_U144 & P3_ADD_339_U143); 
assign P3_ADD_339_U121 = ~P3_ADD_339_U60; 
assign P3_ADD_339_U139 = ~(P3_ADD_339_U60 & P3_PHYADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_541_U72 = ~(P3_ADD_541_U144 & P3_ADD_541_U143); 
assign P3_ADD_541_U121 = ~P3_ADD_541_U60; 
assign P3_ADD_541_U139 = ~(P3_ADD_541_U60 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_515_U72 = ~(P3_ADD_515_U144 & P3_ADD_515_U143); 
assign P3_ADD_515_U121 = ~P3_ADD_515_U60; 
assign P3_ADD_515_U139 = ~(P3_ADD_515_U60 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_394_U71 = ~(P3_ADD_394_U146 & P3_ADD_394_U145); 
assign P3_ADD_394_U124 = ~P3_ADD_394_U60; 
assign P3_ADD_394_U143 = ~(P3_ADD_394_U60 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_441_U72 = ~(P3_ADD_441_U144 & P3_ADD_441_U143); 
assign P3_ADD_441_U121 = ~P3_ADD_441_U60; 
assign P3_ADD_441_U139 = ~(P3_ADD_441_U60 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_349_U76 = ~(P3_ADD_349_U151 & P3_ADD_349_U150); 
assign P3_ADD_349_U125 = ~P3_ADD_349_U61; 
assign P3_ADD_349_U148 = ~(P3_ADD_349_U61 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_405_U71 = ~(P3_ADD_405_U146 & P3_ADD_405_U145); 
assign P3_ADD_405_U124 = ~P3_ADD_405_U60; 
assign P3_ADD_405_U143 = ~(P3_ADD_405_U60 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_553_U76 = ~(P3_ADD_553_U151 & P3_ADD_553_U150); 
assign P3_ADD_553_U125 = ~P3_ADD_553_U61; 
assign P3_ADD_553_U148 = ~(P3_ADD_553_U61 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_558_U76 = ~(P3_ADD_558_U151 & P3_ADD_558_U150); 
assign P3_ADD_558_U125 = ~P3_ADD_558_U61; 
assign P3_ADD_558_U148 = ~(P3_ADD_558_U61 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_385_U76 = ~(P3_ADD_385_U151 & P3_ADD_385_U150); 
assign P3_ADD_385_U125 = ~P3_ADD_385_U61; 
assign P3_ADD_385_U148 = ~(P3_ADD_385_U61 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_547_U76 = ~(P3_ADD_547_U151 & P3_ADD_547_U150); 
assign P3_ADD_547_U125 = ~P3_ADD_547_U61; 
assign P3_ADD_547_U148 = ~(P3_ADD_547_U61 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_494_U72 = ~(P3_ADD_494_U144 & P3_ADD_494_U143); 
assign P3_ADD_494_U121 = ~P3_ADD_494_U60; 
assign P3_ADD_494_U139 = ~(P3_ADD_494_U60 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_536_U72 = ~(P3_ADD_536_U144 & P3_ADD_536_U143); 
assign P3_ADD_536_U121 = ~P3_ADD_536_U60; 
assign P3_ADD_536_U139 = ~(P3_ADD_536_U60 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P2_R2099_U45 = ~(P2_U2728 & P2_R2099_U134); 
assign P2_R2099_U205 = ~(P2_R2099_U134 & P2_R2099_U44); 
assign P2_ADD_391_1196_U53 = ~(P2_ADD_391_1196_U85 & P2_ADD_391_1196_U220); 
assign P2_ADD_391_1196_U137 = P2_ADD_391_1196_U401 & P2_ADD_391_1196_U400; 
assign P2_ADD_391_1196_U219 = ~P2_ADD_391_1196_U85; 
assign P2_ADD_391_1196_U294 = ~(P2_ADD_391_1196_U154 & P2_ADD_391_1196_U217); 
assign P2_ADD_391_1196_U393 = ~(P2_R2096_U84 & P2_ADD_391_1196_U68); 
assign P2_ADD_391_1196_U395 = ~(P2_R2096_U84 & P2_ADD_391_1196_U68); 
assign P2_ADD_391_1196_U404 = ~(P2_ADD_391_1196_U403 & P2_ADD_391_1196_U402); 
assign P2_R2182_U82 = ~(P2_R2182_U265 & P2_R2182_U264); 
assign P2_R2182_U162 = ~P2_R2182_U117; 
assign P2_R2182_U164 = ~(P2_R2182_U163 & P2_R2182_U117); 
assign P2_R2182_U257 = ~(P2_R2182_U116 & P2_R2182_U117); 
assign P2_R2027_U76 = ~(P2_R2027_U151 & P2_R2027_U150); 
assign P2_R2027_U125 = ~P2_R2027_U61; 
assign P2_R2027_U148 = ~(P2_R2027_U61 & P2_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P2_R2337_U69 = ~(P2_R2337_U140 & P2_R2337_U139); 
assign P2_R2337_U122 = ~P2_R2337_U93; 
assign P2_R2337_U137 = ~(P2_R2337_U93 & P2_PHYADDRPOINTER_REG_31__SCAN_IN); 
assign P2_R1957_U36 = ~(P2_R1957_U101 & P2_R1957_U63 & P2_R1957_U39); 
assign P2_R2278_U31 = ~P2_U2793; 
assign P2_R2278_U87 = ~(P2_R2278_U373 & P2_R2278_U372); 
assign P2_R2278_U118 = P2_R2278_U318 & P2_R2278_U229; 
assign P2_R2278_U143 = P2_R2278_U292 & P2_R2278_U296; 
assign P2_R2278_U149 = P2_R2278_U361 & P2_R2278_U360; 
assign P2_R2278_U172 = P2_R2278_U438 & P2_R2278_U437; 
assign P2_R2278_U227 = ~P2_R2278_U150; 
assign P2_R2278_U299 = P2_U2793 | P2_INSTADDRPOINTER_REG_28__SCAN_IN; 
assign P2_R2278_U300 = ~(P2_U2793 & P2_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P2_R2278_U317 = ~(P2_R2278_U117 & P2_R2278_U152); 
assign P2_R2278_U340 = ~(P2_R2278_U294 & P2_R2278_U296); 
assign P2_R2278_U364 = ~(P2_R2278_U363 & P2_R2278_U362); 
assign P2_R2278_U424 = ~(P2_U2793 & P2_R2278_U32); 
assign P2_R2278_U426 = ~(P2_U2793 & P2_R2278_U32); 
assign P2_R2278_U430 = ~(P2_R2278_U74 & P2_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P2_R2278_U432 = ~(P2_R2278_U74 & P2_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P2_R2278_U441 = ~(P2_R2278_U440 & P2_R2278_U439); 
assign P2_ADD_394_U65 = ~(P2_ADD_394_U132 & P2_ADD_394_U131); 
assign P2_ADD_394_U124 = ~P2_ADD_394_U61; 
assign P2_ADD_394_U129 = ~(P2_ADD_394_U61 & P2_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P2_R2267_U16 = P2_R2267_U113 & P2_R2267_U62; 
assign P2_R2267_U112 = ~P2_R2267_U62; 
assign P2_R2267_U141 = ~(P2_U2766 & P2_R2267_U62); 
assign P2_ADD_371_1212_U78 = ~(P2_ADD_371_1212_U213 & P2_ADD_371_1212_U212); 
assign P2_ADD_371_1212_U160 = ~P2_ADD_371_1212_U134; 
assign P2_ADD_371_1212_U162 = ~(P2_ADD_371_1212_U161 & P2_ADD_371_1212_U134); 
assign P2_ADD_371_1212_U202 = ~(P2_ADD_371_1212_U165 & P2_ADD_371_1212_U134 & P2_ADD_371_1212_U161); 
assign P2_ADD_371_1212_U279 = ~(P2_ADD_371_1212_U133 & P2_ADD_371_1212_U134); 
assign P1_R2278_U97 = ~(P1_R2278_U229 & P1_R2278_U331); 
assign P1_R2278_U190 = ~(P1_R2278_U406 & P1_R2278_U405 & P1_R2278_U407 & P1_R2278_U159); 
assign P1_R2278_U194 = ~(P1_R2278_U145 & P1_R2278_U385 & P1_R2278_U146); 
assign P1_R2278_U206 = ~(P1_R2278_U163 & P1_R2278_U376 & P1_R2278_U162); 
assign P1_R2278_U216 = ~(P1_R2278_U169 & P1_R2278_U361); 
assign P1_R2278_U218 = ~(P1_R2278_U360 & P1_R2278_U358); 
assign P1_R2278_U220 = ~(P1_R2278_U290 & P1_R2278_U289); 
assign P1_R2278_U467 = ~(P1_R2278_U397 & P1_R2278_U396 & P1_R2278_U155 & P1_R2278_U187); 
assign P1_R2278_U587 = ~(P1_R2278_U416 & P1_R2278_U585); 
assign P1_R2278_U599 = ~(P1_R2278_U329 & P1_R2278_U597); 
assign P1_R2358_U68 = ~(P1_R2358_U369 & P1_R2358_U291); 
assign P1_R2358_U94 = P1_R2358_U291 & P1_R2358_U290; 
assign P1_R2358_U99 = ~(P1_R2358_U589 & P1_R2358_U588); 
assign P1_R2358_U101 = ~(P1_R2358_U591 & P1_R2358_U590); 
assign P1_R2358_U103 = ~(P1_R2358_U593 & P1_R2358_U592); 
assign P1_R2358_U105 = ~(P1_R2358_U595 & P1_R2358_U594); 
assign P1_R2358_U170 = ~P1_U2655; 
assign P1_R2358_U292 = ~(P1_R2358_U525 & P1_R2358_U524 & P1_R2358_U38); 
assign P1_R2358_U340 = ~(P1_R2358_U291 & P1_R2358_U290); 
assign P1_R2358_U376 = ~P1_R2358_U188; 
assign P1_R2358_U378 = ~P1_R2358_U187; 
assign P1_R2358_U379 = ~(P1_R2358_U9 & P1_R2358_U189); 
assign P1_R2358_U523 = ~(P1_U2655 & P1_R2358_U23); 
assign P1_R2358_U533 = ~(P1_U2655 & P1_R2358_U23); 
assign P1_R2358_U537 = ~(P1_R2358_U536 & P1_R2358_U535); 
assign P1_R2358_U586 = ~(P1_R2358_U188 & P1_R2358_U341); 
assign P1_R2099_U67 = ~(P1_R2099_U301 & P1_R2099_U300); 
assign P1_R2099_U180 = ~P1_R2099_U25; 
assign P1_R2099_U299 = ~(P1_R2099_U44 & P1_R2099_U25); 
assign P1_R2337_U72 = ~(P1_R2337_U144 & P1_R2337_U143); 
assign P1_R2337_U121 = ~P1_R2337_U60; 
assign P1_R2337_U139 = ~(P1_R2337_U60 & P1_PHYADDRPOINTER_REG_30__SCAN_IN); 
assign P1_R2096_U72 = ~(P1_R2096_U144 & P1_R2096_U143); 
assign P1_R2096_U121 = ~P1_R2096_U60; 
assign P1_R2096_U139 = ~(P1_R2096_U60 & P1_REIP_REG_30__SCAN_IN); 
assign P1_ADD_405_U65 = ~(P1_ADD_405_U132 & P1_ADD_405_U131); 
assign P1_ADD_405_U124 = ~P1_ADD_405_U61; 
assign P1_ADD_405_U129 = ~(P1_ADD_405_U61 & P1_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P1_ADD_515_U64 = ~(P1_ADD_515_U128 & P1_ADD_515_U127); 
assign P1_ADD_515_U121 = ~P1_ADD_515_U61; 
assign P1_ADD_515_U125 = ~(P1_ADD_515_U61 & P1_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_U2802 = ~(P3_U6632 & P3_U6631 & P3_U6630 & P3_U6629 & P3_U3982); 
assign P3_U3911 = P3_U3908 & P3_U3907 & P3_U3910 & P3_U3909; 
assign P3_U3930 = P3_U6353 & P3_U6352; 
assign P3_U6278 = ~(P3_U4318 & P3_U6276); 
assign P3_U6306 = ~(P3_ADD_558_U76 & P3_U3220); 
assign P3_U6307 = ~(P3_ADD_553_U76 & P3_U4298); 
assign P3_U6308 = ~(P3_ADD_547_U76 & P3_U4299); 
assign P3_U6311 = ~(P3_ADD_531_U76 & P3_U2354); 
assign P3_U6319 = ~(P3_ADD_385_U76 & P3_U2358); 
assign P3_U6320 = ~(P3_ADD_380_U76 & P3_U2359); 
assign P3_U6321 = ~(P3_ADD_349_U76 & P3_U4306); 
assign P3_U6322 = ~(P3_ADD_344_U76 & P3_U2362); 
assign P3_U6333 = ~(P3_ADD_541_U72 & P3_U4300); 
assign P3_U6334 = ~(P3_ADD_536_U72 & P3_U4301); 
assign P3_U6337 = ~(P3_ADD_515_U72 & P3_U4302); 
assign P3_U6338 = ~(P3_ADD_494_U72 & P3_U2356); 
assign P3_U6339 = ~(P3_ADD_476_U72 & P3_U4303); 
assign P3_U6340 = ~(P3_ADD_441_U72 & P3_U4304); 
assign P3_U6341 = ~(P3_ADD_405_U71 & P3_U4305); 
assign P3_U6342 = ~(P3_ADD_394_U71 & P3_U2357); 
assign P3_U6376 = ~(P3_ADD_360_1242_U90 & P3_U2395); 
assign P3_U6637 = ~(P3_ADD_318_U72 & P3_U2398); 
assign P3_U6642 = ~(P3_ADD_339_U72 & P3_U2388); 
assign P3_U6646 = ~(P3_ADD_315_U68 & P3_U2397); 
assign P3_U6655 = ~(P3_U2396 & P3_ADD_360_1242_U90); 
assign P3_U7342 = ~(P3_ADD_467_U72 & P3_U2601); 
assign P3_U7344 = ~(P3_ADD_430_U72 & P3_U2405); 
assign P2_U2791 = P2_U3242 & P2_R2267_U16; 
assign P2_U2869 = ~(P2_U6526 & P2_U6527 & P2_U6525); 
assign P2_U2907 = ~(P2_U6378 & P2_U6375 & P2_U6377 & P2_U6376); 
assign P2_U6543 = ~(P2_R2182_U82 & P2_U2393); 
assign P2_U6819 = ~(P2_R2267_U16 & P2_U2587); 
assign P2_U8373 = ~(P2_R2337_U69 & P2_U3284); 
assign P1_U2654 = ~(P1_U6784 & P1_U4012); 
assign P1_U2987 = ~(P1_U5861 & P1_U5859 & P1_U5863 & P1_U5860 & P1_U5862); 
assign P1_U2988 = ~(P1_U5856 & P1_U5854 & P1_U5858 & P1_U5855 & P1_U5857); 
assign P1_U2989 = ~(P1_U5851 & P1_U5849 & P1_U5853 & P1_U5850 & P1_U5852); 
assign P1_U3019 = ~(P1_U3802 & P1_U3804 & P1_U5656); 
assign P1_U3020 = ~(P1_U3799 & P1_U3801 & P1_U5649); 
assign P1_U3021 = ~(P1_U3796 & P1_U3798 & P1_U5642); 
assign P1_U5766 = ~(P1_R2099_U67 & P1_U2380); 
assign P1_U5776 = ~(P1_ADD_405_U65 & P1_U2375); 
assign P1_U5777 = ~(P1_ADD_515_U64 & P1_U2374); 
assign P1_U5902 = ~(P1_R2358_U105 & P1_U2364); 
assign P1_U5907 = ~(P1_R2358_U103 & P1_U2364); 
assign P1_U5912 = ~(P1_R2358_U101 & P1_U2364); 
assign P1_U5917 = ~(P1_R2358_U99 & P1_U2364); 
assign P1_U5944 = ~(P1_R2337_U72 & P1_U2376); 
assign P1_U6220 = ~(P1_U2386 & P1_R2358_U105); 
assign P1_U6224 = ~(P1_U2386 & P1_R2358_U103); 
assign P1_U6228 = ~(P1_U2386 & P1_R2358_U101); 
assign P1_U6232 = ~(P1_U2386 & P1_R2358_U99); 
assign P1_U6325 = ~(P1_U2383 & P1_R2358_U105); 
assign P1_U6328 = ~(P1_U2383 & P1_R2358_U103); 
assign P1_U6331 = ~(P1_U2383 & P1_R2358_U101); 
assign P1_U6334 = ~(P1_U2383 & P1_R2358_U99); 
assign P1_U6350 = ~(P1_U2371 & P1_R2099_U67); 
assign P1_U6570 = ~(P1_U2604 & P1_R2099_U67); 
assign P1_U6578 = ~(P1_R2096_U72 & P1_U7485); 
assign P1_U6783 = ~(P1_R2337_U72 & P1_U2352); 
assign P3_ADD_476_U93 = ~(P3_ADD_476_U121 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_476_U140 = ~(P3_ADD_476_U121 & P3_ADD_476_U61); 
assign P3_ADD_531_U63 = ~(P3_ADD_531_U125 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_531_U149 = ~(P3_ADD_531_U125 & P3_ADD_531_U62); 
assign P3_SUB_320_U15 = P3_SUB_320_U108 & P3_SUB_320_U37; 
assign P3_SUB_320_U39 = ~P3_ADD_318_U72; 
assign P3_SUB_320_U102 = ~P3_SUB_320_U37; 
assign P3_SUB_320_U106 = ~(P3_ADD_318_U72 & P3_SUB_320_U37); 
assign P3_ADD_318_U93 = ~(P3_ADD_318_U121 & P3_PHYADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_318_U140 = ~(P3_ADD_318_U121 & P3_ADD_318_U61); 
assign P3_ADD_315_U134 = ~(P3_ADD_315_U118 & P3_ADD_315_U89); 
assign P3_ADD_467_U93 = ~(P3_ADD_467_U121 & P3_REIP_REG_30__SCAN_IN); 
assign P3_ADD_467_U140 = ~(P3_ADD_467_U121 & P3_ADD_467_U61); 
assign P3_ADD_430_U93 = ~(P3_ADD_430_U121 & P3_REIP_REG_30__SCAN_IN); 
assign P3_ADD_430_U140 = ~(P3_ADD_430_U121 & P3_ADD_430_U61); 
assign P3_ADD_380_U63 = ~(P3_ADD_380_U125 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_380_U149 = ~(P3_ADD_380_U125 & P3_ADD_380_U62); 
assign P3_ADD_344_U63 = ~(P3_ADD_344_U125 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_344_U149 = ~(P3_ADD_344_U125 & P3_ADD_344_U62); 
assign P3_ADD_339_U93 = ~(P3_ADD_339_U121 & P3_PHYADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_339_U140 = ~(P3_ADD_339_U121 & P3_ADD_339_U61); 
assign P3_ADD_541_U93 = ~(P3_ADD_541_U121 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_541_U140 = ~(P3_ADD_541_U121 & P3_ADD_541_U61); 
assign P3_ADD_515_U93 = ~(P3_ADD_515_U121 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_515_U140 = ~(P3_ADD_515_U121 & P3_ADD_515_U61); 
assign P3_ADD_394_U95 = ~(P3_ADD_394_U124 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_394_U144 = ~(P3_ADD_394_U124 & P3_ADD_394_U61); 
assign P3_ADD_441_U93 = ~(P3_ADD_441_U121 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_441_U140 = ~(P3_ADD_441_U121 & P3_ADD_441_U61); 
assign P3_ADD_349_U63 = ~(P3_ADD_349_U125 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_349_U149 = ~(P3_ADD_349_U125 & P3_ADD_349_U62); 
assign P3_ADD_405_U95 = ~(P3_ADD_405_U124 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_405_U144 = ~(P3_ADD_405_U124 & P3_ADD_405_U61); 
assign P3_ADD_553_U63 = ~(P3_ADD_553_U125 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_553_U149 = ~(P3_ADD_553_U125 & P3_ADD_553_U62); 
assign P3_ADD_558_U63 = ~(P3_ADD_558_U125 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_558_U149 = ~(P3_ADD_558_U125 & P3_ADD_558_U62); 
assign P3_ADD_385_U63 = ~(P3_ADD_385_U125 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_385_U149 = ~(P3_ADD_385_U125 & P3_ADD_385_U62); 
assign P3_ADD_547_U63 = ~(P3_ADD_547_U125 & P3_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P3_ADD_547_U149 = ~(P3_ADD_547_U125 & P3_ADD_547_U62); 
assign P3_ADD_494_U93 = ~(P3_ADD_494_U121 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_494_U140 = ~(P3_ADD_494_U121 & P3_ADD_494_U61); 
assign P3_ADD_536_U93 = ~(P3_ADD_536_U121 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_536_U140 = ~(P3_ADD_536_U121 & P3_ADD_536_U61); 
assign P2_R2099_U84 = ~(P2_R2099_U205 & P2_R2099_U204); 
assign P2_R2099_U135 = ~P2_R2099_U45; 
assign P2_R2099_U197 = ~(P2_U2727 & P2_R2099_U45); 
assign P2_ADD_391_1196_U70 = ~P2_R2182_U82; 
assign P2_ADD_391_1196_U135 = P2_ADD_391_1196_U394 & P2_ADD_391_1196_U393; 
assign P2_ADD_391_1196_U221 = ~P2_ADD_391_1196_U53; 
assign P2_ADD_391_1196_U260 = P2_R2182_U82 | P2_R2096_U83; 
assign P2_ADD_391_1196_U262 = ~(P2_R2096_U83 & P2_R2182_U82); 
assign P2_ADD_391_1196_U289 = ~(P2_ADD_391_1196_U288 & P2_ADD_391_1196_U53); 
assign P2_ADD_391_1196_U296 = ~(P2_ADD_391_1196_U219 & P2_ADD_391_1196_U295); 
assign P2_ADD_391_1196_U387 = ~(P2_R2182_U82 & P2_ADD_391_1196_U71); 
assign P2_ADD_391_1196_U389 = ~(P2_R2182_U82 & P2_ADD_391_1196_U71); 
assign P2_ADD_391_1196_U397 = ~(P2_ADD_391_1196_U396 & P2_ADD_391_1196_U395); 
assign P2_ADD_391_1196_U459 = ~(P2_ADD_391_1196_U304 & P2_ADD_391_1196_U53); 
assign P2_R2182_U115 = ~(P2_R2182_U165 & P2_R2182_U164); 
assign P2_R2182_U258 = ~(P2_R2182_U162 & P2_R2182_U256); 
assign P2_R2027_U63 = ~(P2_R2027_U125 & P2_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P2_R2027_U149 = ~(P2_R2027_U125 & P2_R2027_U62); 
assign P2_R2337_U138 = ~(P2_R2337_U122 & P2_R2337_U92); 
assign P2_R1957_U15 = P2_R1957_U108 & P2_R1957_U36; 
assign P2_R1957_U38 = ~P2_U3661; 
assign P2_R1957_U102 = ~P2_R1957_U36; 
assign P2_R1957_U106 = ~(P2_U3661 & P2_R1957_U36); 
assign P2_R2278_U33 = ~P2_U2792; 
assign P2_R2278_U81 = ~(P2_R2278_U340 & P2_R2278_U297); 
assign P2_R2278_U136 = P2_R2278_U299 & P2_R2278_U296 & P2_R2278_U292; 
assign P2_R2278_U148 = ~(P2_R2278_U118 & P2_R2278_U317); 
assign P2_R2278_U170 = P2_R2278_U431 & P2_R2278_U430; 
assign P2_R2278_U302 = P2_U2792 | P2_INSTADDRPOINTER_REG_29__SCAN_IN; 
assign P2_R2278_U304 = ~(P2_U2792 & P2_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P2_R2278_U365 = ~(P2_R2278_U149 & P2_R2278_U150); 
assign P2_R2278_U366 = ~(P2_R2278_U227 & P2_R2278_U364); 
assign P2_R2278_U417 = ~(P2_U2792 & P2_R2278_U34); 
assign P2_R2278_U419 = ~(P2_U2792 & P2_R2278_U34); 
assign P2_R2278_U423 = ~(P2_R2278_U31 & P2_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P2_R2278_U425 = ~(P2_R2278_U31 & P2_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P2_R2278_U434 = ~(P2_R2278_U433 & P2_R2278_U432); 
assign P2_ADD_394_U93 = ~(P2_ADD_394_U124 & P2_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P2_ADD_394_U130 = ~(P2_ADD_394_U124 & P2_ADD_394_U60); 
assign P2_R2267_U142 = ~(P2_R2267_U112 & P2_R2267_U61); 
assign P2_ADD_371_1212_U117 = ~(P2_ADD_371_1212_U86 & P2_ADD_371_1212_U202); 
assign P2_ADD_371_1212_U127 = ~(P2_ADD_371_1212_U163 & P2_ADD_371_1212_U162); 
assign P2_ADD_371_1212_U280 = ~(P2_ADD_371_1212_U160 & P2_ADD_371_1212_U278); 
assign P1_R2278_U121 = ~(P1_R2278_U587 & P1_R2278_U586); 
assign P1_R2278_U123 = ~(P1_R2278_U599 & P1_R2278_U598); 
assign P1_R2278_U291 = ~P1_R2278_U220; 
assign P1_R2278_U294 = ~P1_R2278_U218; 
assign P1_R2278_U297 = ~P1_R2278_U216; 
assign P1_R2278_U299 = ~(P1_R2278_U298 & P1_R2278_U216); 
assign P1_R2278_U310 = ~P1_R2278_U206; 
assign P1_R2278_U323 = ~P1_R2278_U194; 
assign P1_R2278_U326 = ~P1_R2278_U190; 
assign P1_R2278_U332 = ~P1_R2278_U97; 
assign P1_R2278_U334 = ~(P1_R2278_U333 & P1_R2278_U97); 
assign P1_R2278_U363 = ~(P1_R2278_U171 & P1_R2278_U216); 
assign P1_R2278_U365 = ~(P1_R2278_U8 & P1_R2278_U216); 
assign P1_R2278_U375 = ~(P1_R2278_U147 & P1_R2278_U194); 
assign P1_R2278_U419 = ~(P1_R2278_U11 & P1_R2278_U206); 
assign P1_R2278_U421 = ~(P1_R2278_U311 & P1_R2278_U206); 
assign P1_R2278_U423 = ~(P1_R2278_U10 & P1_R2278_U206); 
assign P1_R2278_U425 = ~(P1_R2278_U164 & P1_R2278_U206); 
assign P1_R2278_U427 = ~(P1_R2278_U166 & P1_R2278_U206); 
assign P1_R2278_U476 = ~(P1_R2278_U189 & P1_R2278_U190); 
assign P1_R2278_U490 = ~(P1_R2278_U193 & P1_R2278_U194); 
assign P1_R2278_U532 = ~(P1_R2278_U205 & P1_R2278_U206); 
assign P1_R2278_U565 = ~(P1_R2278_U215 & P1_R2278_U216); 
assign P1_R2278_U572 = ~(P1_R2278_U217 & P1_R2278_U218); 
assign P1_R2278_U579 = ~(P1_R2278_U219 & P1_R2278_U220); 
assign P1_R2278_U593 = ~(P1_R2278_U348 & P1_R2278_U97); 
assign P1_R2358_U10 = P1_R2358_U9 & P1_R2358_U292; 
assign P1_R2358_U293 = ~(P1_U2624 & P1_R2358_U537); 
assign P1_R2358_U370 = ~P1_R2358_U68; 
assign P1_R2358_U371 = ~(P1_R2358_U68 & P1_R2358_U292); 
assign P1_R2358_U522 = ~(P1_U2352 & P1_R2358_U170); 
assign P1_R2358_U532 = ~(P1_U2352 & P1_R2358_U170); 
assign P1_R2358_U584 = ~(P1_R2358_U187 & P1_R2358_U340); 
assign P1_R2358_U585 = ~(P1_R2358_U94 & P1_R2358_U378); 
assign P1_R2358_U587 = ~(P1_R2358_U96 & P1_R2358_U376); 
assign P1_R2099_U135 = ~(P1_R2099_U96 & P1_R2099_U180); 
assign P1_R2099_U136 = ~(P1_R2099_U180 & P1_R2099_U44); 
assign P1_R2099_U298 = ~(P1_R2099_U288 & P1_R2099_U180); 
assign P1_R2337_U93 = ~(P1_R2337_U121 & P1_PHYADDRPOINTER_REG_30__SCAN_IN); 
assign P1_R2337_U140 = ~(P1_R2337_U121 & P1_R2337_U61); 
assign P1_R2096_U93 = ~(P1_R2096_U121 & P1_REIP_REG_30__SCAN_IN); 
assign P1_R2096_U140 = ~(P1_R2096_U121 & P1_R2096_U61); 
assign P1_ADD_405_U93 = ~(P1_ADD_405_U124 & P1_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P1_ADD_405_U130 = ~(P1_ADD_405_U124 & P1_ADD_405_U60); 
assign P1_ADD_515_U93 = ~(P1_ADD_515_U121 & P1_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P1_ADD_515_U126 = ~(P1_ADD_515_U121 & P1_ADD_515_U60); 
assign P3_U2836 = ~(P3_U6279 & P3_U6277 & P3_U6278); 
assign P3_U3913 = P3_U6308 & P3_U6307; 
assign P3_U3915 = P3_U6310 & P3_U6309 & P3_U6311 & P3_U3914; 
assign P3_U3918 = P3_U6320 & P3_U6319 & P3_U6321; 
assign P3_U3919 = P3_U6323 & P3_U6322; 
assign P3_U3923 = P3_U6337 & P3_U6336; 
assign P3_U3925 = P3_U6339 & P3_U6338 & P3_U6340; 
assign P3_U3926 = P3_U6342 & P3_U6341; 
assign P3_U3940 = P3_U6377 & P3_U6376; 
assign P3_U3983 = P3_U6644 & P3_U6641 & P3_U6643 & P3_U6642; 
assign P3_U4126 = P3_U7342 & P3_U7341; 
assign P3_U6300 = ~(P3_U3903 & P3_U6282 & P3_U3904 & P3_U3906 & P3_U3911); 
assign P2_U3659 = ~(P2_U8374 & P2_U8373); 
assign P2_U6529 = ~(P2_U2379 & P2_R2099_U84); 
assign P2_U6734 = ~(P2_U2392 & P2_R2099_U84); 
assign P1_U2849 = ~(P1_U6335 & P1_U6336 & P1_U6334); 
assign P1_U2850 = ~(P1_U6332 & P1_U6333 & P1_U6331); 
assign P1_U2851 = ~(P1_U6329 & P1_U6330 & P1_U6328); 
assign P1_U2852 = ~(P1_U6326 & P1_U6327 & P1_U6325); 
assign P1_U2881 = ~(P1_U6231 & P1_U6230 & P1_U6233 & P1_U6232); 
assign P1_U2882 = ~(P1_U6227 & P1_U6226 & P1_U6229 & P1_U6228); 
assign P1_U2883 = ~(P1_U6223 & P1_U6222 & P1_U6225 & P1_U6224); 
assign P1_U2884 = ~(P1_U6219 & P1_U6218 & P1_U6221 & P1_U6220); 
assign P1_U3853 = P1_U5774 & P1_U5776; 
assign P1_U3855 = P1_U3854 & P1_U5777; 
assign P1_U3944 = P1_U6580 & P1_U6578; 
assign P1_U4011 = P1_U6781 & P1_U6782 & P1_U6783; 
assign P1_U5663 = ~(P1_R2278_U123 & P1_U2377); 
assign P1_U5684 = ~(P1_R2278_U121 & P1_U2377); 
assign P1_U5865 = ~(P1_U2372 & P1_R2278_U123); 
assign P1_U5880 = ~(P1_U2372 & P1_R2278_U121); 
assign P3_ADD_476_U70 = ~(P3_ADD_476_U140 & P3_ADD_476_U139); 
assign P3_ADD_476_U122 = ~P3_ADD_476_U93; 
assign P3_ADD_476_U137 = ~(P3_ADD_476_U93 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_531_U75 = ~(P3_ADD_531_U149 & P3_ADD_531_U148); 
assign P3_ADD_531_U126 = ~P3_ADD_531_U63; 
assign P3_ADD_531_U144 = ~(P3_ADD_531_U63 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_SUB_320_U38 = ~(P3_SUB_320_U102 & P3_SUB_320_U39); 
assign P3_ADD_318_U70 = ~(P3_ADD_318_U140 & P3_ADD_318_U139); 
assign P3_ADD_318_U122 = ~P3_ADD_318_U93; 
assign P3_ADD_318_U137 = ~(P3_ADD_318_U93 & P3_PHYADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_315_U67 = ~(P3_ADD_315_U134 & P3_ADD_315_U133); 
assign P3_ADD_467_U70 = ~(P3_ADD_467_U140 & P3_ADD_467_U139); 
assign P3_ADD_467_U122 = ~P3_ADD_467_U93; 
assign P3_ADD_467_U137 = ~(P3_ADD_467_U93 & P3_REIP_REG_31__SCAN_IN); 
assign P3_ADD_430_U70 = ~(P3_ADD_430_U140 & P3_ADD_430_U139); 
assign P3_ADD_430_U122 = ~P3_ADD_430_U93; 
assign P3_ADD_430_U137 = ~(P3_ADD_430_U93 & P3_REIP_REG_31__SCAN_IN); 
assign P3_ADD_380_U75 = ~(P3_ADD_380_U149 & P3_ADD_380_U148); 
assign P3_ADD_380_U126 = ~P3_ADD_380_U63; 
assign P3_ADD_380_U144 = ~(P3_ADD_380_U63 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_344_U75 = ~(P3_ADD_344_U149 & P3_ADD_344_U148); 
assign P3_ADD_344_U126 = ~P3_ADD_344_U63; 
assign P3_ADD_344_U144 = ~(P3_ADD_344_U63 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_339_U70 = ~(P3_ADD_339_U140 & P3_ADD_339_U139); 
assign P3_ADD_339_U122 = ~P3_ADD_339_U93; 
assign P3_ADD_339_U137 = ~(P3_ADD_339_U93 & P3_PHYADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_541_U70 = ~(P3_ADD_541_U140 & P3_ADD_541_U139); 
assign P3_ADD_541_U122 = ~P3_ADD_541_U93; 
assign P3_ADD_541_U137 = ~(P3_ADD_541_U93 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_515_U70 = ~(P3_ADD_515_U140 & P3_ADD_515_U139); 
assign P3_ADD_515_U122 = ~P3_ADD_515_U93; 
assign P3_ADD_515_U137 = ~(P3_ADD_515_U93 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_394_U70 = ~(P3_ADD_394_U144 & P3_ADD_394_U143); 
assign P3_ADD_394_U125 = ~P3_ADD_394_U95; 
assign P3_ADD_394_U141 = ~(P3_ADD_394_U95 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_441_U70 = ~(P3_ADD_441_U140 & P3_ADD_441_U139); 
assign P3_ADD_441_U122 = ~P3_ADD_441_U93; 
assign P3_ADD_441_U137 = ~(P3_ADD_441_U93 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_349_U75 = ~(P3_ADD_349_U149 & P3_ADD_349_U148); 
assign P3_ADD_349_U126 = ~P3_ADD_349_U63; 
assign P3_ADD_349_U144 = ~(P3_ADD_349_U63 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_405_U70 = ~(P3_ADD_405_U144 & P3_ADD_405_U143); 
assign P3_ADD_405_U125 = ~P3_ADD_405_U95; 
assign P3_ADD_405_U141 = ~(P3_ADD_405_U95 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_553_U75 = ~(P3_ADD_553_U149 & P3_ADD_553_U148); 
assign P3_ADD_553_U126 = ~P3_ADD_553_U63; 
assign P3_ADD_553_U144 = ~(P3_ADD_553_U63 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_558_U75 = ~(P3_ADD_558_U149 & P3_ADD_558_U148); 
assign P3_ADD_558_U126 = ~P3_ADD_558_U63; 
assign P3_ADD_558_U144 = ~(P3_ADD_558_U63 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_385_U75 = ~(P3_ADD_385_U149 & P3_ADD_385_U148); 
assign P3_ADD_385_U126 = ~P3_ADD_385_U63; 
assign P3_ADD_385_U144 = ~(P3_ADD_385_U63 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_547_U75 = ~(P3_ADD_547_U149 & P3_ADD_547_U148); 
assign P3_ADD_547_U126 = ~P3_ADD_547_U63; 
assign P3_ADD_547_U144 = ~(P3_ADD_547_U63 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_494_U70 = ~(P3_ADD_494_U140 & P3_ADD_494_U139); 
assign P3_ADD_494_U122 = ~P3_ADD_494_U93; 
assign P3_ADD_494_U137 = ~(P3_ADD_494_U93 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_536_U70 = ~(P3_ADD_536_U140 & P3_ADD_536_U139); 
assign P3_ADD_536_U122 = ~P3_ADD_536_U93; 
assign P3_ADD_536_U137 = ~(P3_ADD_536_U93 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P2_R2099_U47 = ~(P2_U2727 & P2_R2099_U135); 
assign P2_R2099_U198 = ~(P2_R2099_U135 & P2_R2099_U46); 
assign P2_ADD_391_1196_U6 = P2_ADD_391_1196_U296 & P2_ADD_391_1196_U294; 
assign P2_ADD_391_1196_U222 = ~(P2_ADD_391_1196_U221 & P2_ADD_391_1196_U159); 
assign P2_ADD_391_1196_U290 = ~(P2_ADD_391_1196_U289 & P2_ADD_391_1196_U159 & P2_ADD_391_1196_U153); 
assign P2_ADD_391_1196_U386 = ~(P2_R2096_U83 & P2_ADD_391_1196_U70); 
assign P2_ADD_391_1196_U388 = ~(P2_R2096_U83 & P2_ADD_391_1196_U70); 
assign P2_ADD_391_1196_U460 = ~(P2_ADD_391_1196_U458 & P2_ADD_391_1196_U221); 
assign P2_R2182_U81 = ~(P2_R2182_U258 & P2_R2182_U257); 
assign P2_R2182_U166 = ~P2_R2182_U115; 
assign P2_R2182_U168 = ~(P2_R2182_U167 & P2_R2182_U115); 
assign P2_R2182_U250 = ~(P2_R2182_U114 & P2_R2182_U115); 
assign P2_R2027_U75 = ~(P2_R2027_U149 & P2_R2027_U148); 
assign P2_R2027_U126 = ~P2_R2027_U63; 
assign P2_R2027_U144 = ~(P2_R2027_U63 & P2_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P2_R2337_U68 = ~(P2_R2337_U138 & P2_R2337_U137); 
assign P2_R1957_U37 = ~(P2_R1957_U102 & P2_R1957_U38); 
assign P2_R2278_U79 = ~P2_U2791; 
assign P2_R2278_U86 = ~(P2_R2278_U366 & P2_R2278_U365); 
assign P2_R2278_U137 = P2_R2278_U304 & P2_R2278_U300; 
assign P2_R2278_U168 = P2_R2278_U424 & P2_R2278_U423; 
assign P2_R2278_U230 = ~P2_R2278_U148; 
assign P2_R2278_U232 = ~(P2_R2278_U231 & P2_R2278_U148); 
assign P2_R2278_U306 = ~(P2_U2791 & P2_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P2_R2278_U307 = P2_U2791 | P2_INSTADDRPOINTER_REG_30__SCAN_IN; 
assign P2_R2278_U319 = ~(P2_R2278_U119 & P2_R2278_U148); 
assign P2_R2278_U341 = ~P2_R2278_U81; 
assign P2_R2278_U343 = ~(P2_R2278_U81 & P2_R2278_U299); 
assign P2_R2278_U358 = ~(P2_R2278_U147 & P2_R2278_U148); 
assign P2_R2278_U403 = ~(P2_U2791 & P2_R2278_U80); 
assign P2_R2278_U405 = ~(P2_U2791 & P2_R2278_U80); 
assign P2_R2278_U416 = ~(P2_R2278_U33 & P2_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P2_R2278_U418 = ~(P2_R2278_U33 & P2_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P2_R2278_U427 = ~(P2_R2278_U426 & P2_R2278_U425); 
assign P2_ADD_394_U64 = ~(P2_ADD_394_U130 & P2_ADD_394_U129); 
assign P2_ADD_394_U126 = ~P2_ADD_394_U93; 
assign P2_ADD_394_U169 = ~(P2_ADD_394_U93 & P2_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P2_R2267_U63 = P2_R2267_U142 & P2_R2267_U141; 
assign P2_ADD_371_1212_U85 = ~(P2_ADD_371_1212_U280 & P2_ADD_371_1212_U279); 
assign P2_ADD_371_1212_U112 = ~(P2_ADD_371_1212_U12 & P2_ADD_371_1212_U117); 
assign P2_ADD_371_1212_U113 = ~(P2_ADD_371_1212_U9 & P2_ADD_371_1212_U117); 
assign P2_ADD_371_1212_U114 = ~(P2_ADD_371_1212_U95 & P2_ADD_371_1212_U117); 
assign P2_ADD_371_1212_U119 = ~(P2_ADD_371_1212_U117 & P2_ADD_371_1212_U100); 
assign P2_ADD_371_1212_U120 = ~(P2_ADD_371_1212_U105 & P2_ADD_371_1212_U117); 
assign P2_ADD_371_1212_U123 = ~(P2_ADD_371_1212_U8 & P2_ADD_371_1212_U117); 
assign P2_ADD_371_1212_U131 = ~(P2_ADD_371_1212_U6 & P2_ADD_371_1212_U117); 
assign P2_ADD_371_1212_U132 = ~(P2_ADD_371_1212_U102 & P2_ADD_371_1212_U117); 
assign P2_ADD_371_1212_U135 = ~(P2_ADD_371_1212_U109 & P2_ADD_371_1212_U117); 
assign P2_ADD_371_1212_U164 = ~P2_ADD_371_1212_U127; 
assign P2_ADD_371_1212_U167 = ~P2_ADD_371_1212_U117; 
assign P2_ADD_371_1212_U168 = ~(P2_ADD_371_1212_U5 & P2_ADD_371_1212_U117); 
assign P2_ADD_371_1212_U170 = ~(P2_ADD_371_1212_U4 & P2_ADD_371_1212_U117); 
assign P2_ADD_371_1212_U174 = ~(P2_ADD_371_1212_U96 & P2_ADD_371_1212_U117); 
assign P2_ADD_371_1212_U176 = ~(P2_ADD_371_1212_U117 & P2_ADD_371_1212_U97); 
assign P2_ADD_371_1212_U180 = ~(P2_ADD_371_1212_U117 & P2_ADD_371_1212_U93); 
assign P2_ADD_371_1212_U184 = ~(P2_ADD_371_1212_U10 & P2_ADD_371_1212_U117); 
assign P2_ADD_371_1212_U186 = ~(P2_ADD_371_1212_U99 & P2_ADD_371_1212_U117); 
assign P2_ADD_371_1212_U189 = ~(P2_ADD_371_1212_U117 & P2_ADD_371_1212_U103); 
assign P2_ADD_371_1212_U193 = ~(P2_ADD_371_1212_U11 & P2_ADD_371_1212_U117); 
assign P2_ADD_371_1212_U195 = ~(P2_ADD_371_1212_U117 & P2_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P2_ADD_371_1212_U197 = ~(P2_ADD_371_1212_U108 & P2_ADD_371_1212_U117); 
assign P2_ADD_371_1212_U199 = ~(P2_ADD_371_1212_U7 & P2_ADD_371_1212_U117); 
assign P2_ADD_371_1212_U201 = ~(P2_ADD_371_1212_U107 & P2_ADD_371_1212_U117); 
assign P2_ADD_371_1212_U227 = ~(P2_ADD_371_1212_U117 & P2_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P2_ADD_371_1212_U254 = ~(P2_ADD_371_1212_U126 & P2_ADD_371_1212_U127); 
assign P2_ADD_371_1212_U257 = ~(P2_ADD_371_1212_U106 & P2_ADD_371_1212_U117 & P2_ADD_371_1212_U128); 
assign P1_R2278_U16 = P1_R2278_U188 & P1_R2278_U375 & P1_R2278_U468 & P1_R2278_U467; 
assign P1_R2278_U196 = ~(P1_R2278_U419 & P1_R2278_U409); 
assign P1_R2278_U198 = ~(P1_R2278_U425 & P1_R2278_U373); 
assign P1_R2278_U200 = ~(P1_R2278_U165 & P1_R2278_U423); 
assign P1_R2278_U202 = ~(P1_R2278_U167 & P1_R2278_U427); 
assign P1_R2278_U204 = ~(P1_R2278_U421 & P1_R2278_U312); 
assign P1_R2278_U208 = ~(P1_R2278_U170 & P1_R2278_U365); 
assign P1_R2278_U210 = ~(P1_R2278_U172 & P1_R2278_U363); 
assign P1_R2278_U212 = ~(P1_R2278_U300 & P1_R2278_U299); 
assign P1_R2278_U335 = ~(P1_R2278_U173 & P1_R2278_U334); 
assign P1_R2278_U336 = ~(P1_R2278_U332 & P1_R2278_U285); 
assign P1_R2278_U477 = ~(P1_R2278_U326 & P1_R2278_U475); 
assign P1_R2278_U491 = ~(P1_R2278_U323 & P1_R2278_U489); 
assign P1_R2278_U533 = ~(P1_R2278_U310 & P1_R2278_U531); 
assign P1_R2278_U566 = ~(P1_R2278_U297 & P1_R2278_U564); 
assign P1_R2278_U573 = ~(P1_R2278_U294 & P1_R2278_U571); 
assign P1_R2278_U580 = ~(P1_R2278_U291 & P1_R2278_U578); 
assign P1_R2278_U594 = ~(P1_R2278_U592 & P1_R2278_U332); 
assign P1_R2358_U67 = ~(P1_R2358_U371 & P1_R2358_U293); 
assign P1_R2358_U92 = P1_R2358_U293 & P1_R2358_U292; 
assign P1_R2358_U95 = ~(P1_R2358_U585 & P1_R2358_U584); 
assign P1_R2358_U97 = ~(P1_R2358_U587 & P1_R2358_U586); 
assign P1_R2358_U175 = ~P1_U2654; 
assign P1_R2358_U186 = ~(P1_R2358_U370 & P1_R2358_U379); 
assign P1_R2358_U294 = ~(P1_R2358_U523 & P1_R2358_U522 & P1_R2358_U37); 
assign P1_R2358_U339 = ~(P1_R2358_U293 & P1_R2358_U292); 
assign P1_R2358_U381 = ~(P1_R2358_U10 & P1_R2358_U189); 
assign P1_R2358_U534 = ~(P1_R2358_U533 & P1_R2358_U532); 
assign P1_R2358_U548 = ~(P1_U2654 & P1_R2358_U23); 
assign P1_R2358_U550 = ~(P1_U2654 & P1_R2358_U23); 
assign P1_R2099_U66 = ~(P1_R2099_U299 & P1_R2099_U298); 
assign P1_R2099_U145 = ~P1_R2099_U135; 
assign P1_R2099_U181 = ~P1_R2099_U136; 
assign P1_R2099_U293 = ~(P1_R2099_U97 & P1_R2099_U135); 
assign P1_R2099_U295 = ~(P1_R2099_U43 & P1_R2099_U136); 
assign P1_R2337_U70 = ~(P1_R2337_U140 & P1_R2337_U139); 
assign P1_R2337_U122 = ~P1_R2337_U93; 
assign P1_R2337_U137 = ~(P1_R2337_U93 & P1_PHYADDRPOINTER_REG_31__SCAN_IN); 
assign P1_R2096_U70 = ~(P1_R2096_U140 & P1_R2096_U139); 
assign P1_R2096_U122 = ~P1_R2096_U93; 
assign P1_R2096_U137 = ~(P1_R2096_U93 & P1_REIP_REG_31__SCAN_IN); 
assign P1_ADD_405_U64 = ~(P1_ADD_405_U130 & P1_ADD_405_U129); 
assign P1_ADD_405_U126 = ~P1_ADD_405_U93; 
assign P1_ADD_405_U169 = ~(P1_ADD_405_U93 & P1_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P1_ADD_515_U63 = ~(P1_ADD_515_U126 & P1_ADD_515_U125); 
assign P1_ADD_515_U122 = ~P1_ADD_515_U93; 
assign P1_ADD_515_U167 = ~(P1_ADD_515_U93 & P1_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_U2801 = ~(P3_U6640 & P3_U6639 & P3_U6638 & P3_U6637 & P3_U3983); 
assign P3_U3920 = P3_U3917 & P3_U3916 & P3_U3919 & P3_U3918; 
assign P3_U6302 = ~(P3_U4318 & P3_U6300); 
assign P3_U6330 = ~(P3_ADD_558_U75 & P3_U3220); 
assign P3_U6331 = ~(P3_ADD_553_U75 & P3_U4298); 
assign P3_U6332 = ~(P3_ADD_547_U75 & P3_U4299); 
assign P3_U6335 = ~(P3_ADD_531_U75 & P3_U2354); 
assign P3_U6343 = ~(P3_ADD_385_U75 & P3_U2358); 
assign P3_U6344 = ~(P3_ADD_380_U75 & P3_U2359); 
assign P3_U6345 = ~(P3_ADD_349_U75 & P3_U4306); 
assign P3_U6346 = ~(P3_ADD_344_U75 & P3_U2362); 
assign P3_U6357 = ~(P3_ADD_541_U70 & P3_U4300); 
assign P3_U6358 = ~(P3_ADD_536_U70 & P3_U4301); 
assign P3_U6361 = ~(P3_ADD_515_U70 & P3_U4302); 
assign P3_U6362 = ~(P3_ADD_494_U70 & P3_U2356); 
assign P3_U6363 = ~(P3_ADD_476_U70 & P3_U4303); 
assign P3_U6364 = ~(P3_ADD_441_U70 & P3_U4304); 
assign P3_U6365 = ~(P3_ADD_405_U70 & P3_U4305); 
assign P3_U6366 = ~(P3_ADD_394_U70 & P3_U2357); 
assign P3_U6645 = ~(P3_ADD_318_U70 & P3_U2398); 
assign P3_U6650 = ~(P3_ADD_339_U70 & P3_U2388); 
assign P3_U6654 = ~(P3_ADD_315_U67 & P3_U2397); 
assign P3_U7350 = ~(P3_ADD_467_U70 & P3_U2601); 
assign P3_U7352 = ~(P3_ADD_430_U70 & P3_U2405); 
assign P2_U2790 = P2_U3242 & P2_R2267_U63; 
assign P2_U2868 = ~(P2_U6529 & P2_U6530 & P2_U6528); 
assign P2_U6380 = ~(P2_ADD_391_1196_U6 & P2_U2397); 
assign P2_U6546 = ~(P2_R2182_U81 & P2_U2393); 
assign P2_U6827 = ~(P2_R2267_U63 & P2_U2587); 
assign P2_U8349 = ~(P2_R2337_U68 & P2_U3284); 
assign P1_U2653 = ~(P1_U6780 & P1_U4011); 
assign P1_U2983 = ~(P1_U5881 & P1_U5879 & P1_U5883 & P1_U5880 & P1_U5882); 
assign P1_U2986 = ~(P1_U5866 & P1_U5864 & P1_U5868 & P1_U5865 & P1_U5867); 
assign P1_U3015 = ~(P1_U3816 & P1_U3814 & P1_U5682 & P1_U5684); 
assign P1_U3018 = ~(P1_U3807 & P1_U3805 & P1_U5661 & P1_U5663); 
assign P1_U5773 = ~(P1_R2099_U66 & P1_U2380); 
assign P1_U5783 = ~(P1_ADD_405_U64 & P1_U2375); 
assign P1_U5784 = ~(P1_ADD_515_U63 & P1_U2374); 
assign P1_U5789 = ~(P1_R2278_U16 & P1_U2377); 
assign P1_U5922 = ~(P1_R2358_U97 & P1_U2364); 
assign P1_U5927 = ~(P1_R2358_U95 & P1_U2364); 
assign P1_U5949 = ~(P1_R2337_U70 & P1_U2376); 
assign P1_U5955 = ~(P1_U2372 & P1_R2278_U16); 
assign P1_U6236 = ~(P1_U2386 & P1_R2358_U97); 
assign P1_U6240 = ~(P1_U2386 & P1_R2358_U95); 
assign P1_U6337 = ~(P1_U2383 & P1_R2358_U97); 
assign P1_U6340 = ~(P1_U2383 & P1_R2358_U95); 
assign P1_U6353 = ~(P1_U2371 & P1_R2099_U66); 
assign P1_U6577 = ~(P1_U2604 & P1_R2099_U66); 
assign P1_U6585 = ~(P1_R2096_U70 & P1_U7485); 
assign P1_U6774 = ~(P1_R2337_U70 & P1_U2352); 
assign P3_ADD_476_U138 = ~(P3_ADD_476_U122 & P3_ADD_476_U92); 
assign P3_ADD_531_U97 = ~(P3_ADD_531_U126 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_531_U145 = ~(P3_ADD_531_U126 & P3_ADD_531_U64); 
assign P3_SUB_320_U16 = P3_SUB_320_U106 & P3_SUB_320_U38; 
assign P3_SUB_320_U61 = ~P3_ADD_318_U70; 
assign P3_SUB_320_U103 = ~P3_SUB_320_U38; 
assign P3_SUB_320_U138 = ~(P3_ADD_318_U70 & P3_SUB_320_U38); 
assign P3_ADD_318_U138 = ~(P3_ADD_318_U122 & P3_ADD_318_U92); 
assign P3_ADD_467_U138 = ~(P3_ADD_467_U122 & P3_ADD_467_U92); 
assign P3_ADD_430_U138 = ~(P3_ADD_430_U122 & P3_ADD_430_U92); 
assign P3_ADD_380_U97 = ~(P3_ADD_380_U126 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_380_U145 = ~(P3_ADD_380_U126 & P3_ADD_380_U64); 
assign P3_ADD_344_U97 = ~(P3_ADD_344_U126 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_344_U145 = ~(P3_ADD_344_U126 & P3_ADD_344_U64); 
assign P3_ADD_339_U138 = ~(P3_ADD_339_U122 & P3_ADD_339_U92); 
assign P3_ADD_541_U138 = ~(P3_ADD_541_U122 & P3_ADD_541_U92); 
assign P3_ADD_515_U138 = ~(P3_ADD_515_U122 & P3_ADD_515_U92); 
assign P3_ADD_394_U142 = ~(P3_ADD_394_U125 & P3_ADD_394_U94); 
assign P3_ADD_441_U138 = ~(P3_ADD_441_U122 & P3_ADD_441_U92); 
assign P3_ADD_349_U97 = ~(P3_ADD_349_U126 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_349_U145 = ~(P3_ADD_349_U126 & P3_ADD_349_U64); 
assign P3_ADD_405_U142 = ~(P3_ADD_405_U125 & P3_ADD_405_U94); 
assign P3_ADD_553_U97 = ~(P3_ADD_553_U126 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_553_U145 = ~(P3_ADD_553_U126 & P3_ADD_553_U64); 
assign P3_ADD_558_U97 = ~(P3_ADD_558_U126 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_558_U145 = ~(P3_ADD_558_U126 & P3_ADD_558_U64); 
assign P3_ADD_385_U97 = ~(P3_ADD_385_U126 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_385_U145 = ~(P3_ADD_385_U126 & P3_ADD_385_U64); 
assign P3_ADD_547_U97 = ~(P3_ADD_547_U126 & P3_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P3_ADD_547_U145 = ~(P3_ADD_547_U126 & P3_ADD_547_U64); 
assign P3_ADD_494_U138 = ~(P3_ADD_494_U122 & P3_ADD_494_U92); 
assign P3_ADD_536_U138 = ~(P3_ADD_536_U122 & P3_ADD_536_U92); 
assign P2_R2099_U83 = ~(P2_R2099_U198 & P2_R2099_U197); 
assign P2_R2099_U136 = ~P2_R2099_U47; 
assign P2_R2099_U195 = ~(P2_U2726 & P2_R2099_U47); 
assign P2_ADD_391_1196_U72 = ~P2_R2182_U81; 
assign P2_ADD_391_1196_U83 = ~(P2_ADD_391_1196_U224 & P2_ADD_391_1196_U222 & P2_ADD_391_1196_U223); 
assign P2_ADD_391_1196_U107 = ~(P2_ADD_391_1196_U460 & P2_ADD_391_1196_U459); 
assign P2_ADD_391_1196_U133 = P2_ADD_391_1196_U387 & P2_ADD_391_1196_U386; 
assign P2_ADD_391_1196_U264 = P2_R2182_U81 | P2_R2096_U82; 
assign P2_ADD_391_1196_U266 = ~(P2_R2096_U82 & P2_R2182_U81); 
assign P2_ADD_391_1196_U380 = ~(P2_R2182_U81 & P2_ADD_391_1196_U73); 
assign P2_ADD_391_1196_U382 = ~(P2_R2182_U81 & P2_ADD_391_1196_U73); 
assign P2_ADD_391_1196_U390 = ~(P2_ADD_391_1196_U389 & P2_ADD_391_1196_U388); 
assign P2_R2182_U113 = ~(P2_R2182_U169 & P2_R2182_U168); 
assign P2_R2182_U251 = ~(P2_R2182_U166 & P2_R2182_U249); 
assign P2_R2027_U97 = ~(P2_R2027_U126 & P2_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P2_R2027_U145 = ~(P2_R2027_U126 & P2_R2027_U64); 
assign P2_R1957_U16 = P2_R1957_U106 & P2_R1957_U37; 
assign P2_R1957_U61 = ~P2_U3659; 
assign P2_R1957_U103 = ~P2_R1957_U37; 
assign P2_R1957_U138 = ~(P2_U3659 & P2_R1957_U37); 
assign P2_R2278_U138 = P2_R2278_U307 & P2_R2278_U302; 
assign P2_R2278_U140 = P2_R2278_U343 & P2_R2278_U300; 
assign P2_R2278_U142 = P2_R2278_U304 & P2_R2278_U306; 
assign P2_R2278_U146 = ~(P2_R2278_U49 & P2_R2278_U232); 
assign P2_R2278_U166 = P2_R2278_U417 & P2_R2278_U416; 
assign P2_R2278_U204 = ~(P2_R2278_U120 & P2_R2278_U319); 
assign P2_R2278_U359 = ~(P2_R2278_U230 & P2_R2278_U357); 
assign P2_R2278_U402 = ~(P2_R2278_U79 & P2_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P2_R2278_U404 = ~(P2_R2278_U79 & P2_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P2_R2278_U420 = ~(P2_R2278_U419 & P2_R2278_U418); 
assign P2_ADD_394_U170 = ~(P2_ADD_394_U126 & P2_ADD_394_U92); 
assign P2_ADD_371_1212_U169 = ~P2_ADD_371_1212_U132; 
assign P2_ADD_371_1212_U171 = ~P2_ADD_371_1212_U120; 
assign P2_ADD_371_1212_U172 = ~P2_ADD_371_1212_U114; 
assign P2_ADD_371_1212_U173 = ~P2_ADD_371_1212_U119; 
assign P2_ADD_371_1212_U175 = ~P2_ADD_371_1212_U131; 
assign P2_ADD_371_1212_U177 = ~P2_ADD_371_1212_U113; 
assign P2_ADD_371_1212_U178 = ~P2_ADD_371_1212_U135; 
assign P2_ADD_371_1212_U179 = ~P2_ADD_371_1212_U123; 
assign P2_ADD_371_1212_U181 = ~P2_ADD_371_1212_U112; 
assign P2_ADD_371_1212_U182 = ~(P2_ADD_371_1212_U65 & P2_ADD_371_1212_U180); 
assign P2_ADD_371_1212_U183 = ~(P2_ADD_371_1212_U56 & P2_ADD_371_1212_U174); 
assign P2_ADD_371_1212_U185 = ~(P2_ADD_371_1212_U49 & P2_ADD_371_1212_U184); 
assign P2_ADD_371_1212_U187 = ~(P2_ADD_371_1212_U58 & P2_ADD_371_1212_U186); 
assign P2_ADD_371_1212_U188 = ~(P2_ADD_371_1212_U47 & P2_ADD_371_1212_U168); 
assign P2_ADD_371_1212_U190 = ~(P2_ADD_371_1212_U61 & P2_ADD_371_1212_U189); 
assign P2_ADD_371_1212_U191 = ~(P2_ADD_371_1212_U50 & P2_ADD_371_1212_U170); 
assign P2_ADD_371_1212_U192 = ~(P2_ADD_371_1212_U59 & P2_ADD_371_1212_U176); 
assign P2_ADD_371_1212_U194 = ~(P2_ADD_371_1212_U55 & P2_ADD_371_1212_U193); 
assign P2_ADD_371_1212_U196 = ~(P2_ADD_371_1212_U46 & P2_ADD_371_1212_U195); 
assign P2_ADD_371_1212_U198 = ~(P2_ADD_371_1212_U64 & P2_ADD_371_1212_U197); 
assign P2_ADD_371_1212_U200 = ~(P2_ADD_371_1212_U52 & P2_ADD_371_1212_U199); 
assign P2_ADD_371_1212_U214 = ~(P2_ADD_371_1212_U112 & P2_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P2_ADD_371_1212_U216 = ~(P2_ADD_371_1212_U113 & P2_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P2_ADD_371_1212_U218 = ~(P2_ADD_371_1212_U114 & P2_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P2_ADD_371_1212_U228 = ~(P2_ADD_371_1212_U167 & P2_ADD_371_1212_U45); 
assign P2_ADD_371_1212_U229 = ~(P2_ADD_371_1212_U119 & P2_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P2_ADD_371_1212_U231 = ~(P2_ADD_371_1212_U120 & P2_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P2_ADD_371_1212_U240 = ~(P2_ADD_371_1212_U123 & P2_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P2_ADD_371_1212_U255 = ~(P2_ADD_371_1212_U164 & P2_ADD_371_1212_U253); 
assign P2_ADD_371_1212_U256 = ~(P2_ADD_371_1212_U201 & P2_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P2_ADD_371_1212_U270 = ~(P2_ADD_371_1212_U131 & P2_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P2_ADD_371_1212_U272 = ~(P2_ADD_371_1212_U132 & P2_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P2_ADD_371_1212_U281 = ~(P2_ADD_371_1212_U135 & P2_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P1_R2278_U106 = ~(P1_R2278_U477 & P1_R2278_U476); 
assign P1_R2278_U108 = ~(P1_R2278_U491 & P1_R2278_U490); 
assign P1_R2278_U114 = ~(P1_R2278_U533 & P1_R2278_U532); 
assign P1_R2278_U118 = ~(P1_R2278_U566 & P1_R2278_U565); 
assign P1_R2278_U119 = ~(P1_R2278_U573 & P1_R2278_U572); 
assign P1_R2278_U120 = ~(P1_R2278_U580 & P1_R2278_U579); 
assign P1_R2278_U122 = ~(P1_R2278_U594 & P1_R2278_U593); 
assign P1_R2278_U301 = ~P1_R2278_U212; 
assign P1_R2278_U304 = ~P1_R2278_U210; 
assign P1_R2278_U307 = ~P1_R2278_U208; 
assign P1_R2278_U414 = ~(P1_R2278_U174 & P1_R2278_U336); 
assign P1_R2278_U420 = ~P1_R2278_U196; 
assign P1_R2278_U422 = ~P1_R2278_U204; 
assign P1_R2278_U424 = ~P1_R2278_U200; 
assign P1_R2278_U426 = ~P1_R2278_U198; 
assign P1_R2278_U428 = ~P1_R2278_U202; 
assign P1_R2278_U497 = ~(P1_R2278_U195 & P1_R2278_U196); 
assign P1_R2278_U504 = ~(P1_R2278_U197 & P1_R2278_U198); 
assign P1_R2278_U511 = ~(P1_R2278_U199 & P1_R2278_U200); 
assign P1_R2278_U518 = ~(P1_R2278_U201 & P1_R2278_U202); 
assign P1_R2278_U525 = ~(P1_R2278_U203 & P1_R2278_U204); 
assign P1_R2278_U539 = ~(P1_R2278_U207 & P1_R2278_U208); 
assign P1_R2278_U546 = ~(P1_R2278_U209 & P1_R2278_U210); 
assign P1_R2278_U553 = ~(P1_R2278_U211 & P1_R2278_U212); 
assign P1_R2358_U132 = P1_R2358_U10 & P1_R2358_U294; 
assign P1_R2358_U295 = ~(P1_U2623 & P1_R2358_U534); 
assign P1_R2358_U372 = ~P1_R2358_U67; 
assign P1_R2358_U373 = ~(P1_R2358_U67 & P1_R2358_U294); 
assign P1_R2358_U380 = ~P1_R2358_U186; 
assign P1_R2358_U547 = ~(P1_U2352 & P1_R2358_U175); 
assign P1_R2358_U549 = ~(P1_U2352 & P1_R2358_U175); 
assign P1_R2358_U582 = ~(P1_R2358_U186 & P1_R2358_U339); 
assign P1_R2099_U292 = ~(P1_R2099_U145 & P1_R2099_U291); 
assign P1_R2099_U294 = ~(P1_R2099_U181 & P1_R2099_U285); 
assign P1_R2337_U138 = ~(P1_R2337_U122 & P1_R2337_U92); 
assign P1_R2096_U138 = ~(P1_R2096_U122 & P1_R2096_U92); 
assign P1_ADD_405_U170 = ~(P1_ADD_405_U126 & P1_ADD_405_U92); 
assign P1_ADD_515_U168 = ~(P1_ADD_515_U122 & P1_ADD_515_U92); 
assign P3_U2835 = ~(P3_U6303 & P3_U6301 & P3_U6302); 
assign P3_U3922 = P3_U6332 & P3_U6331; 
assign P3_U3924 = P3_U6334 & P3_U6333 & P3_U6335 & P3_U3923; 
assign P3_U3927 = P3_U6344 & P3_U6343 & P3_U6345; 
assign P3_U3928 = P3_U6347 & P3_U6346; 
assign P3_U3932 = P3_U6361 & P3_U6360; 
assign P3_U3934 = P3_U6363 & P3_U6362 & P3_U6364; 
assign P3_U3935 = P3_U6366 & P3_U6365; 
assign P3_U3984 = P3_U6652 & P3_U6649 & P3_U6651 & P3_U6650; 
assign P3_U4129 = P3_U7350 & P3_U7349; 
assign P3_U6324 = ~(P3_U3912 & P3_U6306 & P3_U3913 & P3_U3915 & P3_U3920); 
assign P2_U2906 = ~(P2_U6382 & P2_U6379 & P2_U6381 & P2_U6380); 
assign P2_U3647 = ~(P2_U8350 & P2_U8349); 
assign P2_U6384 = ~(P2_ADD_391_1196_U107 & P2_U2397); 
assign P2_U6532 = ~(P2_U2379 & P2_R2099_U83); 
assign P2_U6742 = ~(P2_U2392 & P2_R2099_U83); 
assign P1_U2847 = ~(P1_U6341 & P1_U6342 & P1_U6340); 
assign P1_U2848 = ~(P1_U6338 & P1_U6339 & P1_U6337); 
assign P1_U2879 = ~(P1_U6239 & P1_U6238 & P1_U6241 & P1_U6240); 
assign P1_U2880 = ~(P1_U6235 & P1_U6234 & P1_U6237 & P1_U6236); 
assign P1_U3856 = P1_U5781 & P1_U5783; 
assign P1_U3858 = P1_U3857 & P1_U5784; 
assign P1_U3946 = P1_U6587 & P1_U6585; 
assign P1_U4009 = P1_U6772 & P1_U6773 & P1_U6774; 
assign P1_U5670 = ~(P1_R2278_U122 & P1_U2377); 
assign P1_U5691 = ~(P1_R2278_U120 & P1_U2377); 
assign P1_U5698 = ~(P1_R2278_U119 & P1_U2377); 
assign P1_U5705 = ~(P1_R2278_U118 & P1_U2377); 
assign P1_U5733 = ~(P1_R2278_U114 & P1_U2377); 
assign P1_U5775 = ~(P1_R2278_U108 & P1_U2377); 
assign P1_U5782 = ~(P1_R2278_U106 & P1_U2377); 
assign P1_U5870 = ~(P1_U2372 & P1_R2278_U122); 
assign P1_U5885 = ~(P1_U2372 & P1_R2278_U120); 
assign P1_U5890 = ~(P1_U2372 & P1_R2278_U119); 
assign P1_U5895 = ~(P1_U2372 & P1_R2278_U118); 
assign P1_U5915 = ~(P1_U2372 & P1_R2278_U114); 
assign P1_U5945 = ~(P1_U2372 & P1_R2278_U108); 
assign P1_U5950 = ~(P1_U2372 & P1_R2278_U106); 
assign P3_ADD_476_U69 = ~(P3_ADD_476_U138 & P3_ADD_476_U137); 
assign P3_ADD_531_U73 = ~(P3_ADD_531_U145 & P3_ADD_531_U144); 
assign P3_ADD_531_U127 = ~P3_ADD_531_U97; 
assign P3_ADD_531_U142 = ~(P3_ADD_531_U97 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_SUB_320_U127 = ~(P3_SUB_320_U103 & P3_SUB_320_U61); 
assign P3_SUB_320_U139 = ~(P3_SUB_320_U103 & P3_SUB_320_U61); 
assign P3_ADD_318_U69 = ~(P3_ADD_318_U138 & P3_ADD_318_U137); 
assign P3_ADD_467_U69 = ~(P3_ADD_467_U138 & P3_ADD_467_U137); 
assign P3_ADD_430_U69 = ~(P3_ADD_430_U138 & P3_ADD_430_U137); 
assign P3_ADD_380_U73 = ~(P3_ADD_380_U145 & P3_ADD_380_U144); 
assign P3_ADD_380_U127 = ~P3_ADD_380_U97; 
assign P3_ADD_380_U142 = ~(P3_ADD_380_U97 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_344_U73 = ~(P3_ADD_344_U145 & P3_ADD_344_U144); 
assign P3_ADD_344_U127 = ~P3_ADD_344_U97; 
assign P3_ADD_344_U142 = ~(P3_ADD_344_U97 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_339_U69 = ~(P3_ADD_339_U138 & P3_ADD_339_U137); 
assign P3_ADD_541_U69 = ~(P3_ADD_541_U138 & P3_ADD_541_U137); 
assign P3_ADD_515_U69 = ~(P3_ADD_515_U138 & P3_ADD_515_U137); 
assign P3_ADD_394_U69 = ~(P3_ADD_394_U142 & P3_ADD_394_U141); 
assign P3_ADD_441_U69 = ~(P3_ADD_441_U138 & P3_ADD_441_U137); 
assign P3_ADD_349_U73 = ~(P3_ADD_349_U145 & P3_ADD_349_U144); 
assign P3_ADD_349_U127 = ~P3_ADD_349_U97; 
assign P3_ADD_349_U142 = ~(P3_ADD_349_U97 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_405_U69 = ~(P3_ADD_405_U142 & P3_ADD_405_U141); 
assign P3_ADD_553_U73 = ~(P3_ADD_553_U145 & P3_ADD_553_U144); 
assign P3_ADD_553_U127 = ~P3_ADD_553_U97; 
assign P3_ADD_553_U142 = ~(P3_ADD_553_U97 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_558_U73 = ~(P3_ADD_558_U145 & P3_ADD_558_U144); 
assign P3_ADD_558_U127 = ~P3_ADD_558_U97; 
assign P3_ADD_558_U142 = ~(P3_ADD_558_U97 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_385_U73 = ~(P3_ADD_385_U145 & P3_ADD_385_U144); 
assign P3_ADD_385_U127 = ~P3_ADD_385_U97; 
assign P3_ADD_385_U142 = ~(P3_ADD_385_U97 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_547_U73 = ~(P3_ADD_547_U145 & P3_ADD_547_U144); 
assign P3_ADD_547_U127 = ~P3_ADD_547_U97; 
assign P3_ADD_547_U142 = ~(P3_ADD_547_U97 & P3_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P3_ADD_494_U69 = ~(P3_ADD_494_U138 & P3_ADD_494_U137); 
assign P3_ADD_536_U69 = ~(P3_ADD_536_U138 & P3_ADD_536_U137); 
assign P2_R2099_U49 = ~(P2_U2726 & P2_R2099_U136); 
assign P2_R2099_U196 = ~(P2_R2099_U136 & P2_R2099_U48); 
assign P2_ADD_391_1196_U152 = ~(P2_ADD_391_1196_U83 & P2_ADD_391_1196_U226); 
assign P2_ADD_391_1196_U225 = ~P2_ADD_391_1196_U83; 
assign P2_ADD_391_1196_U379 = ~(P2_R2096_U82 & P2_ADD_391_1196_U72); 
assign P2_ADD_391_1196_U381 = ~(P2_R2096_U82 & P2_ADD_391_1196_U72); 
assign P2_R2182_U80 = ~(P2_R2182_U251 & P2_R2182_U250); 
assign P2_R2182_U170 = ~P2_R2182_U113; 
assign P2_R2182_U172 = ~(P2_R2182_U171 & P2_R2182_U113); 
assign P2_R2182_U243 = ~(P2_R2182_U112 & P2_R2182_U113); 
assign P2_R2027_U73 = ~(P2_R2027_U145 & P2_R2027_U144); 
assign P2_R2027_U127 = ~P2_R2027_U97; 
assign P2_R2027_U142 = ~(P2_R2027_U97 & P2_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P2_R1957_U127 = ~(P2_R1957_U103 & P2_R1957_U61); 
assign P2_R1957_U139 = ~(P2_R1957_U103 & P2_R1957_U61); 
assign P2_R2278_U85 = ~(P2_R2278_U359 & P2_R2278_U358); 
assign P2_R2278_U160 = ~P2_U2790; 
assign P2_R2278_U162 = P2_R2278_U403 & P2_R2278_U402; 
assign P2_R2278_U234 = ~P2_R2278_U146; 
assign P2_R2278_U237 = ~P2_R2278_U204; 
assign P2_R2278_U239 = ~(P2_R2278_U238 & P2_R2278_U204); 
assign P2_R2278_U321 = ~(P2_R2278_U121 & P2_R2278_U204); 
assign P2_R2278_U351 = ~(P2_R2278_U145 & P2_R2278_U146); 
assign P2_R2278_U396 = ~(P2_U2790 & P2_R2278_U159); 
assign P2_R2278_U399 = ~(P2_U2790 & P2_R2278_U159); 
assign P2_R2278_U406 = ~(P2_R2278_U405 & P2_R2278_U404); 
assign P2_R2278_U559 = ~(P2_R2278_U203 & P2_R2278_U204); 
assign P2_ADD_394_U84 = ~(P2_ADD_394_U170 & P2_ADD_394_U169); 
assign P2_ADD_371_1212_U13 = P2_ADD_371_1212_U196 & P2_ADD_371_1212_U168; 
assign P2_ADD_371_1212_U14 = P2_ADD_371_1212_U188 & P2_ADD_371_1212_U132; 
assign P2_ADD_371_1212_U15 = P2_ADD_371_1212_U185 & P2_ADD_371_1212_U170; 
assign P2_ADD_371_1212_U16 = P2_ADD_371_1212_U191 & P2_ADD_371_1212_U120; 
assign P2_ADD_371_1212_U17 = P2_ADD_371_1212_U200 & P2_ADD_371_1212_U114; 
assign P2_ADD_371_1212_U18 = P2_ADD_371_1212_U194 & P2_ADD_371_1212_U174; 
assign P2_ADD_371_1212_U19 = P2_ADD_371_1212_U183 & P2_ADD_371_1212_U131; 
assign P2_ADD_371_1212_U20 = P2_ADD_371_1212_U187 & P2_ADD_371_1212_U176; 
assign P2_ADD_371_1212_U21 = P2_ADD_371_1212_U192 & P2_ADD_371_1212_U113; 
assign P2_ADD_371_1212_U22 = P2_ADD_371_1212_U190 & P2_ADD_371_1212_U123; 
assign P2_ADD_371_1212_U23 = P2_ADD_371_1212_U198 & P2_ADD_371_1212_U180; 
assign P2_ADD_371_1212_U24 = P2_ADD_371_1212_U182 & P2_ADD_371_1212_U112; 
assign P2_ADD_371_1212_U82 = ~(P2_ADD_371_1212_U255 & P2_ADD_371_1212_U254); 
assign P2_ADD_371_1212_U83 = ~(P2_ADD_371_1212_U257 & P2_ADD_371_1212_U256); 
assign P2_ADD_371_1212_U118 = P2_ADD_371_1212_U228 & P2_ADD_371_1212_U227; 
assign P2_ADD_371_1212_U215 = ~(P2_ADD_371_1212_U181 & P2_ADD_371_1212_U66); 
assign P2_ADD_371_1212_U217 = ~(P2_ADD_371_1212_U177 & P2_ADD_371_1212_U60); 
assign P2_ADD_371_1212_U219 = ~(P2_ADD_371_1212_U172 & P2_ADD_371_1212_U54); 
assign P2_ADD_371_1212_U230 = ~(P2_ADD_371_1212_U173 & P2_ADD_371_1212_U53); 
assign P2_ADD_371_1212_U232 = ~(P2_ADD_371_1212_U171 & P2_ADD_371_1212_U51); 
assign P2_ADD_371_1212_U241 = ~(P2_ADD_371_1212_U179 & P2_ADD_371_1212_U63); 
assign P2_ADD_371_1212_U271 = ~(P2_ADD_371_1212_U175 & P2_ADD_371_1212_U57); 
assign P2_ADD_371_1212_U273 = ~(P2_ADD_371_1212_U169 & P2_ADD_371_1212_U48); 
assign P2_ADD_371_1212_U282 = ~(P2_ADD_371_1212_U178 & P2_ADD_371_1212_U62); 
assign P1_R2278_U20 = P1_R2278_U414 & P1_R2278_U335; 
assign P1_R2278_U498 = ~(P1_R2278_U420 & P1_R2278_U496); 
assign P1_R2278_U505 = ~(P1_R2278_U426 & P1_R2278_U503); 
assign P1_R2278_U512 = ~(P1_R2278_U424 & P1_R2278_U510); 
assign P1_R2278_U519 = ~(P1_R2278_U428 & P1_R2278_U517); 
assign P1_R2278_U526 = ~(P1_R2278_U422 & P1_R2278_U524); 
assign P1_R2278_U540 = ~(P1_R2278_U307 & P1_R2278_U538); 
assign P1_R2278_U547 = ~(P1_R2278_U304 & P1_R2278_U545); 
assign P1_R2278_U554 = ~(P1_R2278_U301 & P1_R2278_U552); 
assign P1_R2358_U90 = P1_R2358_U295 & P1_R2358_U294; 
assign P1_R2358_U133 = P1_R2358_U373 & P1_R2358_U295; 
assign P1_R2358_U176 = ~P1_U2653; 
assign P1_R2358_U185 = ~(P1_R2358_U372 & P1_R2358_U381); 
assign P1_R2358_U296 = ~(P1_R2358_U548 & P1_R2358_U547 & P1_R2358_U62); 
assign P1_R2358_U338 = ~(P1_R2358_U295 & P1_R2358_U294); 
assign P1_R2358_U383 = ~(P1_R2358_U132 & P1_R2358_U189); 
assign P1_R2358_U551 = ~(P1_R2358_U550 & P1_R2358_U549); 
assign P1_R2358_U553 = ~(P1_U2653 & P1_R2358_U23); 
assign P1_R2358_U563 = ~(P1_U2653 & P1_R2358_U23); 
assign P1_R2358_U583 = ~(P1_R2358_U92 & P1_R2358_U380); 
assign P1_R2099_U64 = ~(P1_R2099_U293 & P1_R2099_U292); 
assign P1_R2099_U65 = ~(P1_R2099_U295 & P1_R2099_U294); 
assign P1_R2337_U69 = ~(P1_R2337_U138 & P1_R2337_U137); 
assign P1_R2096_U69 = ~(P1_R2096_U138 & P1_R2096_U137); 
assign P1_ADD_405_U84 = ~(P1_ADD_405_U170 & P1_ADD_405_U169); 
assign P1_ADD_515_U84 = ~(P1_ADD_515_U168 & P1_ADD_515_U167); 
assign P3_U2800 = ~(P3_U6648 & P3_U6647 & P3_U6646 & P3_U6645 & P3_U3984); 
assign P3_U3258 = ~P3_ADD_318_U69; 
assign P3_U3259 = ~(P3_ADD_318_U69 & P3_U2385); 
assign P3_U3929 = P3_U3926 & P3_U3925 & P3_U3928 & P3_U3927; 
assign P3_U6326 = ~(P3_U4318 & P3_U6324); 
assign P3_U6354 = ~(P3_ADD_558_U73 & P3_U3220); 
assign P3_U6355 = ~(P3_ADD_553_U73 & P3_U4298); 
assign P3_U6356 = ~(P3_ADD_547_U73 & P3_U4299); 
assign P3_U6359 = ~(P3_ADD_531_U73 & P3_U2354); 
assign P3_U6367 = ~(P3_ADD_385_U73 & P3_U2358); 
assign P3_U6368 = ~(P3_ADD_380_U73 & P3_U2359); 
assign P3_U6369 = ~(P3_ADD_349_U73 & P3_U4306); 
assign P3_U6370 = ~(P3_ADD_344_U73 & P3_U2362); 
assign P3_U6381 = ~(P3_ADD_541_U69 & P3_U4300); 
assign P3_U6382 = ~(P3_ADD_536_U69 & P3_U4301); 
assign P3_U6385 = ~(P3_ADD_515_U69 & P3_U4302); 
assign P3_U6386 = ~(P3_ADD_494_U69 & P3_U2356); 
assign P3_U6387 = ~(P3_ADD_476_U69 & P3_U4303); 
assign P3_U6388 = ~(P3_ADD_441_U69 & P3_U4304); 
assign P3_U6389 = ~(P3_ADD_405_U69 & P3_U4305); 
assign P3_U6390 = ~(P3_ADD_394_U69 & P3_U2357); 
assign P3_U6653 = ~(P3_ADD_318_U69 & P3_U2398); 
assign P3_U6658 = ~(P3_ADD_339_U69 & P3_U2388); 
assign P3_U7359 = ~(P3_ADD_467_U69 & P3_U2601); 
assign P3_U7361 = ~(P3_ADD_430_U69 & P3_U2405); 
assign P2_U2382 = P2_U2366 & P2_U3647; 
assign P2_U2867 = ~(P2_U6532 & P2_U6533 & P2_U6531); 
assign P2_U2905 = ~(P2_U6386 & P2_U6383 & P2_U6385 & P2_U6384); 
assign P2_U3528 = ~P2_U3647; 
assign P2_U6549 = ~(P2_R2182_U80 & P2_U2393); 
assign P2_U8086 = ~(P2_U3647 & P2_U3683); 
assign P2_U8089 = ~(P2_R1957_U49 & P2_U3647); 
assign P1_U2367 = P1_U3431 & P1_R2337_U69 & P1_STATE2_REG_1__SCAN_IN; 
assign P1_U2652 = ~(P1_U6771 & P1_U4009); 
assign P1_U2976 = ~(P1_U5916 & P1_U5914 & P1_U5918 & P1_U5915 & P1_U5917); 
assign P1_U2980 = ~(P1_U5896 & P1_U5894 & P1_U5898 & P1_U5895 & P1_U5897); 
assign P1_U2981 = ~(P1_U5891 & P1_U5889 & P1_U5893 & P1_U5890 & P1_U5892); 
assign P1_U2982 = ~(P1_U5886 & P1_U5884 & P1_U5888 & P1_U5885 & P1_U5887); 
assign P1_U2985 = ~(P1_U5871 & P1_U5869 & P1_U5873 & P1_U5870 & P1_U5872); 
assign P1_U3002 = ~(P1_U3855 & P1_U3853 & P1_U5773 & P1_U5775); 
assign P1_U3008 = ~(P1_U3837 & P1_U3835 & P1_U5731 & P1_U5733); 
assign P1_U3012 = ~(P1_U3825 & P1_U3823 & P1_U5703 & P1_U5705); 
assign P1_U3013 = ~(P1_U3822 & P1_U3820 & P1_U5696 & P1_U5698); 
assign P1_U3014 = ~(P1_U3819 & P1_U3817 & P1_U5689 & P1_U5691); 
assign P1_U3017 = ~(P1_U3810 & P1_U3808 & P1_U5668 & P1_U5670); 
assign P1_U3430 = ~P1_R2337_U69; 
assign P1_U5677 = ~(P1_R2278_U20 & P1_U2377); 
assign P1_U5780 = ~(P1_R2099_U65 & P1_U2380); 
assign P1_U5787 = ~(P1_R2099_U64 & P1_U2380); 
assign P1_U5790 = ~(P1_ADD_405_U84 & P1_U2375); 
assign P1_U5791 = ~(P1_ADD_515_U84 & P1_U2374); 
assign P1_U5875 = ~(P1_U2372 & P1_R2278_U20); 
assign P1_U5954 = ~(P1_R2337_U69 & P1_U2376); 
assign P1_U6356 = ~(P1_U2371 & P1_R2099_U65); 
assign P1_U6358 = ~(P1_U2371 & P1_R2099_U64); 
assign P1_U6365 = ~(P1_R2337_U69 & P1_STATE2_REG_1__SCAN_IN); 
assign P1_U6584 = ~(P1_U2604 & P1_R2099_U65); 
assign P1_U6591 = ~(P1_U2604 & P1_R2099_U64); 
assign P1_U6592 = ~(P1_R2096_U69 & P1_U7485); 
assign P1_U6770 = ~(P1_R2337_U69 & P1_U2352); 
assign P3_ADD_531_U143 = ~(P3_ADD_531_U127 & P3_ADD_531_U96); 
assign P3_SUB_320_U60 = ~P3_ADD_318_U69; 
assign P3_SUB_320_U62 = P3_SUB_320_U139 & P3_SUB_320_U138; 
assign P3_SUB_320_U137 = ~(P3_SUB_320_U103 & P3_SUB_320_U61 & P3_ADD_318_U69); 
assign P3_ADD_380_U143 = ~(P3_ADD_380_U127 & P3_ADD_380_U96); 
assign P3_ADD_344_U143 = ~(P3_ADD_344_U127 & P3_ADD_344_U96); 
assign P3_ADD_349_U143 = ~(P3_ADD_349_U127 & P3_ADD_349_U96); 
assign P3_ADD_553_U143 = ~(P3_ADD_553_U127 & P3_ADD_553_U96); 
assign P3_ADD_558_U143 = ~(P3_ADD_558_U127 & P3_ADD_558_U96); 
assign P3_ADD_385_U143 = ~(P3_ADD_385_U127 & P3_ADD_385_U96); 
assign P3_ADD_547_U143 = ~(P3_ADD_547_U127 & P3_ADD_547_U96); 
assign P2_R2099_U82 = ~(P2_R2099_U196 & P2_R2099_U195); 
assign P2_R2099_U137 = ~P2_R2099_U49; 
assign P2_R2099_U193 = ~(P2_U2725 & P2_R2099_U49); 
assign P2_ADD_391_1196_U74 = ~P2_R2182_U80; 
assign P2_ADD_391_1196_U131 = P2_ADD_391_1196_U380 & P2_ADD_391_1196_U379; 
assign P2_ADD_391_1196_U227 = ~P2_ADD_391_1196_U152; 
assign P2_ADD_391_1196_U229 = ~(P2_ADD_391_1196_U228 & P2_ADD_391_1196_U152); 
assign P2_ADD_391_1196_U268 = P2_R2182_U80 | P2_R2096_U81; 
assign P2_ADD_391_1196_U270 = ~(P2_R2096_U81 & P2_R2182_U80); 
assign P2_ADD_391_1196_U292 = ~(P2_ADD_391_1196_U225 & P2_ADD_391_1196_U291); 
assign P2_ADD_391_1196_U373 = ~(P2_R2182_U80 & P2_ADD_391_1196_U75); 
assign P2_ADD_391_1196_U375 = ~(P2_R2182_U80 & P2_ADD_391_1196_U75); 
assign P2_ADD_391_1196_U383 = ~(P2_ADD_391_1196_U382 & P2_ADD_391_1196_U381); 
assign P2_ADD_391_1196_U452 = ~(P2_ADD_391_1196_U151 & P2_ADD_391_1196_U152); 
assign P2_R2182_U111 = ~(P2_R2182_U173 & P2_R2182_U172); 
assign P2_R2182_U244 = ~(P2_R2182_U170 & P2_R2182_U242); 
assign P2_R2027_U143 = ~(P2_R2027_U127 & P2_R2027_U96); 
assign P2_R1957_U60 = ~P2_U3647; 
assign P2_R1957_U62 = P2_R1957_U139 & P2_R1957_U138; 
assign P2_R1957_U137 = ~(P2_R1957_U103 & P2_R1957_U61 & P2_U3647); 
assign P2_R2278_U200 = ~(P2_R2278_U122 & P2_R2278_U321); 
assign P2_R2278_U202 = ~(P2_R2278_U52 & P2_R2278_U239); 
assign P2_R2278_U352 = ~(P2_R2278_U234 & P2_R2278_U350); 
assign P2_R2278_U395 = ~(P2_R2278_U160 & P2_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P2_R2278_U398 = ~(P2_R2278_U160 & P2_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P2_R2278_U560 = ~(P2_R2278_U237 & P2_R2278_U558); 
assign P2_ADD_371_1212_U69 = ~(P2_ADD_371_1212_U215 & P2_ADD_371_1212_U214); 
assign P2_ADD_371_1212_U70 = ~(P2_ADD_371_1212_U217 & P2_ADD_371_1212_U216); 
assign P2_ADD_371_1212_U71 = ~(P2_ADD_371_1212_U219 & P2_ADD_371_1212_U218); 
assign P2_ADD_371_1212_U72 = ~(P2_ADD_371_1212_U230 & P2_ADD_371_1212_U229); 
assign P2_ADD_371_1212_U73 = ~(P2_ADD_371_1212_U232 & P2_ADD_371_1212_U231); 
assign P2_ADD_371_1212_U74 = ~(P2_ADD_371_1212_U241 & P2_ADD_371_1212_U240); 
assign P2_ADD_371_1212_U75 = ~(P2_ADD_371_1212_U271 & P2_ADD_371_1212_U270); 
assign P2_ADD_371_1212_U76 = ~(P2_ADD_371_1212_U273 & P2_ADD_371_1212_U272); 
assign P2_ADD_371_1212_U77 = ~(P2_ADD_371_1212_U282 & P2_ADD_371_1212_U281); 
assign P1_R2278_U109 = ~(P1_R2278_U498 & P1_R2278_U497); 
assign P1_R2278_U110 = ~(P1_R2278_U505 & P1_R2278_U504); 
assign P1_R2278_U111 = ~(P1_R2278_U512 & P1_R2278_U511); 
assign P1_R2278_U112 = ~(P1_R2278_U519 & P1_R2278_U518); 
assign P1_R2278_U113 = ~(P1_R2278_U526 & P1_R2278_U525); 
assign P1_R2278_U115 = ~(P1_R2278_U540 & P1_R2278_U539); 
assign P1_R2278_U116 = ~(P1_R2278_U547 & P1_R2278_U546); 
assign P1_R2278_U117 = ~(P1_R2278_U554 & P1_R2278_U553); 
assign P1_R2358_U93 = ~(P1_R2358_U583 & P1_R2358_U582); 
assign P1_R2358_U184 = ~(P1_R2358_U133 & P1_R2358_U383); 
assign P1_R2358_U297 = ~(P1_U2622 & P1_R2358_U551); 
assign P1_R2358_U382 = ~P1_R2358_U185; 
assign P1_R2358_U552 = ~(P1_U2352 & P1_R2358_U176); 
assign P1_R2358_U562 = ~(P1_U2352 & P1_R2358_U176); 
assign P1_R2358_U580 = ~(P1_R2358_U185 & P1_R2358_U338); 
assign P3_U2403 = P3_U2385 & P3_U3258; 
assign P3_U2834 = ~(P3_U6327 & P3_U6325 & P3_U6326); 
assign P3_U3931 = P3_U6356 & P3_U6355; 
assign P3_U3933 = P3_U6358 & P3_U6357 & P3_U6359 & P3_U3932; 
assign P3_U3936 = P3_U6368 & P3_U6367 & P3_U6369; 
assign P3_U3937 = P3_U6371 & P3_U6370; 
assign P3_U3943 = P3_U6386 & P3_U6385 & P3_U6384; 
assign P3_U3946 = P3_U6388 & P3_U6387 & P3_U6389; 
assign P3_U3985 = P3_U6660 & P3_U6657 & P3_U6659 & P3_U6658; 
assign P3_U4133 = P3_U4132 & P3_U7361; 
assign P3_U4319 = ~P3_U3259; 
assign P3_U6348 = ~(P3_U3921 & P3_U6330 & P3_U3922 & P3_U3924 & P3_U3929); 
assign P2_U2383 = P2_U2366 & P2_U3528; 
assign P2_U6535 = ~(P2_U2379 & P2_R2099_U82); 
assign P2_U6579 = ~(P2_U2382 & P2_U3683); 
assign P2_U6588 = ~(P2_U2382 & P2_R1957_U49); 
assign P2_U6597 = ~(P2_R1957_U17 & P2_U2382); 
assign P2_U6606 = ~(P2_R1957_U59 & P2_U2382); 
assign P2_U6615 = ~(P2_R1957_U18 & P2_U2382); 
assign P2_U6624 = ~(P2_R1957_U57 & P2_U2382); 
assign P2_U6632 = ~(P2_R1957_U19 & P2_U2382); 
assign P2_U6640 = ~(P2_R1957_U55 & P2_U2382); 
assign P2_U6648 = ~(P2_R1957_U20 & P2_U2382); 
assign P2_U6656 = ~(P2_R1957_U53 & P2_U2382); 
assign P2_U6664 = ~(P2_R1957_U6 & P2_U2382); 
assign P2_U6672 = ~(P2_R1957_U82 & P2_U2382); 
assign P2_U6680 = ~(P2_R1957_U7 & P2_U2382); 
assign P2_U6688 = ~(P2_R1957_U80 & P2_U2382); 
assign P2_U6696 = ~(P2_R1957_U8 & P2_U2382); 
assign P2_U6704 = ~(P2_R1957_U78 & P2_U2382); 
assign P2_U6712 = ~(P2_R1957_U9 & P2_U2382); 
assign P2_U6720 = ~(P2_R1957_U76 & P2_U2382); 
assign P2_U6728 = ~(P2_R1957_U10 & P2_U2382); 
assign P2_U6736 = ~(P2_R1957_U74 & P2_U2382); 
assign P2_U6744 = ~(P2_R1957_U11 & P2_U2382); 
assign P2_U6750 = ~(P2_U2392 & P2_R2099_U82); 
assign P2_U6752 = ~(P2_R1957_U70 & P2_U2382); 
assign P2_U6760 = ~(P2_R1957_U12 & P2_U2382); 
assign P2_U6768 = ~(P2_R1957_U68 & P2_U2382); 
assign P2_U6776 = ~(P2_R1957_U13 & P2_U2382); 
assign P2_U6784 = ~(P2_R1957_U66 & P2_U2382); 
assign P2_U6792 = ~(P2_R1957_U14 & P2_U2382); 
assign P2_U6800 = ~(P2_R1957_U64 & P2_U2382); 
assign P2_U6808 = ~(P2_R1957_U15 & P2_U2382); 
assign P2_U6816 = ~(P2_R1957_U16 & P2_U2382); 
assign P2_U6824 = ~(P2_R1957_U62 & P2_U2382); 
assign P2_U8085 = ~(P2_U3528 & P2_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P2_U8088 = ~(P2_U3528 & P2_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P1_U2366 = P1_U3431 & P1_U3430 & P1_STATE2_REG_1__SCAN_IN; 
assign P1_U2651 = ~(P1_U6769 & P1_U6768 & P1_U6770); 
assign P1_U2841 = ~(P1_U6359 & P1_U6358); 
assign P1_U2984 = ~(P1_U5876 & P1_U5874 & P1_U5878 & P1_U5875 & P1_U5877); 
assign P1_U3001 = ~(P1_U3858 & P1_U3856 & P1_U5780 & P1_U5782); 
assign P1_U3016 = ~(P1_U3813 & P1_U3811 & P1_U5675 & P1_U5677); 
assign P1_U3859 = P1_U5788 & P1_U5790; 
assign P1_U3861 = P1_U3860 & P1_U5791; 
assign P1_U3948 = P1_U6594 & P1_U6592; 
assign P1_U5712 = ~(P1_R2278_U117 & P1_U2377); 
assign P1_U5719 = ~(P1_R2278_U116 & P1_U2377); 
assign P1_U5726 = ~(P1_R2278_U115 & P1_U2377); 
assign P1_U5740 = ~(P1_R2278_U113 & P1_U2377); 
assign P1_U5747 = ~(P1_R2278_U112 & P1_U2377); 
assign P1_U5754 = ~(P1_R2278_U111 & P1_U2377); 
assign P1_U5761 = ~(P1_R2278_U110 & P1_U2377); 
assign P1_U5768 = ~(P1_R2278_U109 & P1_U2377); 
assign P1_U5900 = ~(P1_U2372 & P1_R2278_U117); 
assign P1_U5905 = ~(P1_U2372 & P1_R2278_U116); 
assign P1_U5910 = ~(P1_U2372 & P1_R2278_U115); 
assign P1_U5920 = ~(P1_U2372 & P1_R2278_U113); 
assign P1_U5925 = ~(P1_U2372 & P1_R2278_U112); 
assign P1_U5930 = ~(P1_U2372 & P1_R2278_U111); 
assign P1_U5932 = ~(P1_R2358_U93 & P1_U2364); 
assign P1_U5935 = ~(P1_U2372 & P1_R2278_U110); 
assign P1_U5940 = ~(P1_U2372 & P1_R2278_U109); 
assign P1_U6244 = ~(P1_U2386 & P1_R2358_U93); 
assign P1_U6343 = ~(P1_U2383 & P1_R2358_U93); 
assign P1_U6366 = ~(P1_U6365 & P1_U6364); 
assign P1_U6420 = ~(P1_U2367 & P1_R2358_U20); 
assign P1_U6427 = ~(P1_U2367 & P1_R2358_U21); 
assign P1_U6434 = ~(P1_U2367 & P1_R2358_U80); 
assign P1_U6441 = ~(P1_U2367 & P1_R2358_U78); 
assign P1_U6448 = ~(P1_U2367 & P1_R2358_U14); 
assign P1_U6455 = ~(P1_U2367 & P1_R2358_U15); 
assign P1_U6462 = ~(P1_U2367 & P1_R2358_U119); 
assign P1_U6469 = ~(P1_U2367 & P1_R2358_U117); 
assign P1_U6476 = ~(P1_U2367 & P1_R2358_U16); 
assign P1_U6483 = ~(P1_U2367 & P1_R2358_U17); 
assign P1_U6490 = ~(P1_U2367 & P1_R2358_U115); 
assign P1_U6497 = ~(P1_U2367 & P1_R2358_U113); 
assign P1_U6504 = ~(P1_U2367 & P1_R2358_U111); 
assign P1_U6511 = ~(P1_U2367 & P1_R2358_U109); 
assign P1_U6518 = ~(P1_U2367 & P1_R2358_U105); 
assign P1_U6525 = ~(P1_U2367 & P1_R2358_U103); 
assign P1_U6532 = ~(P1_U2367 & P1_R2358_U101); 
assign P1_U6539 = ~(P1_U2367 & P1_R2358_U99); 
assign P1_U6546 = ~(P1_U2367 & P1_R2358_U97); 
assign P1_U6553 = ~(P1_U2367 & P1_R2358_U95); 
assign P1_U6560 = ~(P1_U2367 & P1_R2358_U93); 
assign P3_ADD_531_U72 = ~(P3_ADD_531_U143 & P3_ADD_531_U142); 
assign P3_SUB_320_U136 = ~(P3_SUB_320_U127 & P3_SUB_320_U60); 
assign P3_ADD_380_U72 = ~(P3_ADD_380_U143 & P3_ADD_380_U142); 
assign P3_ADD_344_U72 = ~(P3_ADD_344_U143 & P3_ADD_344_U142); 
assign P3_ADD_349_U72 = ~(P3_ADD_349_U143 & P3_ADD_349_U142); 
assign P3_ADD_553_U72 = ~(P3_ADD_553_U143 & P3_ADD_553_U142); 
assign P3_ADD_558_U72 = ~(P3_ADD_558_U143 & P3_ADD_558_U142); 
assign P3_ADD_385_U72 = ~(P3_ADD_385_U143 & P3_ADD_385_U142); 
assign P3_ADD_547_U72 = ~(P3_ADD_547_U143 & P3_ADD_547_U142); 
assign P2_R2099_U51 = ~(P2_U2725 & P2_R2099_U137); 
assign P2_R2099_U194 = ~(P2_R2099_U137 & P2_R2099_U50); 
assign P2_ADD_391_1196_U7 = P2_ADD_391_1196_U292 & P2_ADD_391_1196_U290; 
assign P2_ADD_391_1196_U150 = ~(P2_ADD_391_1196_U230 & P2_ADD_391_1196_U229); 
assign P2_ADD_391_1196_U372 = ~(P2_R2096_U81 & P2_ADD_391_1196_U74); 
assign P2_ADD_391_1196_U374 = ~(P2_R2096_U81 & P2_ADD_391_1196_U74); 
assign P2_ADD_391_1196_U453 = ~(P2_ADD_391_1196_U227 & P2_ADD_391_1196_U451); 
assign P2_R2182_U79 = ~(P2_R2182_U244 & P2_R2182_U243); 
assign P2_R2182_U174 = ~P2_R2182_U111; 
assign P2_R2182_U176 = ~(P2_R2182_U175 & P2_R2182_U111); 
assign P2_R2182_U236 = ~(P2_R2182_U110 & P2_R2182_U111); 
assign P2_R2027_U72 = ~(P2_R2027_U143 & P2_R2027_U142); 
assign P2_R1957_U136 = ~(P2_R1957_U127 & P2_R1957_U60); 
assign P2_R2278_U4 = P2_R2278_U399 & P2_R2278_U398; 
assign P2_R2278_U84 = ~(P2_R2278_U352 & P2_R2278_U351); 
assign P2_R2278_U112 = ~(P2_R2278_U560 & P2_R2278_U559); 
assign P2_R2278_U241 = ~P2_R2278_U202; 
assign P2_R2278_U244 = ~P2_R2278_U200; 
assign P2_R2278_U246 = ~(P2_R2278_U245 & P2_R2278_U200); 
assign P2_R2278_U323 = ~(P2_R2278_U123 & P2_R2278_U200); 
assign P2_R2278_U397 = ~(P2_R2278_U396 & P2_R2278_U395); 
assign P2_R2278_U545 = ~(P2_R2278_U199 & P2_R2278_U200); 
assign P2_R2278_U552 = ~(P2_R2278_U201 & P2_R2278_U202); 
assign P1_R2358_U88 = P1_R2358_U297 & P1_R2358_U296; 
assign P1_R2358_U178 = ~P1_U2652; 
assign P1_R2358_U298 = ~(P1_R2358_U296 & P1_R2358_U184); 
assign P1_R2358_U300 = ~(P1_R2358_U553 & P1_R2358_U552 & P1_R2358_U64); 
assign P1_R2358_U337 = ~(P1_R2358_U297 & P1_R2358_U296); 
assign P1_R2358_U384 = ~P1_R2358_U184; 
assign P1_R2358_U557 = ~(P1_U2652 & P1_R2358_U23); 
assign P1_R2358_U564 = ~(P1_R2358_U563 & P1_R2358_U562); 
assign P1_R2358_U581 = ~(P1_R2358_U90 & P1_R2358_U382); 
assign P3_U2603 = P3_U7360 & P3_U7358 & P3_U7359 & P3_U4133; 
assign P3_U2799 = ~(P3_U6656 & P3_U6654 & P3_U6655 & P3_U6653 & P3_U3985); 
assign P3_U3938 = P3_U3935 & P3_U3934 & P3_U3937 & P3_U3936; 
assign P3_U6350 = ~(P3_U4318 & P3_U6348); 
assign P3_U6378 = ~(P3_ADD_558_U72 & P3_U3220); 
assign P3_U6379 = ~(P3_ADD_553_U72 & P3_U4298); 
assign P3_U6380 = ~(P3_ADD_547_U72 & P3_U4299); 
assign P3_U6383 = ~(P3_ADD_531_U72 & P3_U2354); 
assign P3_U6391 = ~(P3_ADD_385_U72 & P3_U2358); 
assign P3_U6392 = ~(P3_ADD_380_U72 & P3_U2359); 
assign P3_U6393 = ~(P3_ADD_349_U72 & P3_U4306); 
assign P3_U6394 = ~(P3_ADD_344_U72 & P3_U2362); 
assign P3_U7103 = ~(P3_U2403 & P3_PHYADDRPOINTER_REG_0__SCAN_IN); 
assign P3_U7104 = ~(P3_U4319 & P3_PHYADDRPOINTER_REG_0__SCAN_IN); 
assign P3_U7113 = ~(P3_U2403 & P3_ADD_318_U4); 
assign P3_U7114 = ~(P3_SUB_320_U50 & P3_U4319); 
assign P3_U7123 = ~(P3_U2403 & P3_ADD_318_U71); 
assign P3_U7124 = ~(P3_SUB_320_U17 & P3_U4319); 
assign P3_U7133 = ~(P3_U2403 & P3_ADD_318_U68); 
assign P3_U7134 = ~(P3_SUB_320_U59 & P3_U4319); 
assign P3_U7143 = ~(P3_U2403 & P3_ADD_318_U67); 
assign P3_U7144 = ~(P3_SUB_320_U18 & P3_U4319); 
assign P3_U7153 = ~(P3_U2403 & P3_ADD_318_U66); 
assign P3_U7154 = ~(P3_SUB_320_U57 & P3_U4319); 
assign P3_U7161 = ~(P3_U2403 & P3_ADD_318_U65); 
assign P3_U7162 = ~(P3_SUB_320_U19 & P3_U4319); 
assign P3_U7169 = ~(P3_U2403 & P3_ADD_318_U64); 
assign P3_U7170 = ~(P3_SUB_320_U55 & P3_U4319); 
assign P3_U7177 = ~(P3_U2403 & P3_ADD_318_U63); 
assign P3_U7178 = ~(P3_SUB_320_U20 & P3_U4319); 
assign P3_U7185 = ~(P3_U2403 & P3_ADD_318_U62); 
assign P3_U7186 = ~(P3_SUB_320_U53 & P3_U4319); 
assign P3_U7193 = ~(P3_U2403 & P3_ADD_318_U91); 
assign P3_U7194 = ~(P3_SUB_320_U6 & P3_U4319); 
assign P3_U7201 = ~(P3_U2403 & P3_ADD_318_U90); 
assign P3_U7202 = ~(P3_SUB_320_U82 & P3_U4319); 
assign P3_U7209 = ~(P3_U2403 & P3_ADD_318_U89); 
assign P3_U7210 = ~(P3_SUB_320_U7 & P3_U4319); 
assign P3_U7217 = ~(P3_U2403 & P3_ADD_318_U88); 
assign P3_U7218 = ~(P3_SUB_320_U80 & P3_U4319); 
assign P3_U7225 = ~(P3_U2403 & P3_ADD_318_U87); 
assign P3_U7226 = ~(P3_SUB_320_U8 & P3_U4319); 
assign P3_U7233 = ~(P3_U2403 & P3_ADD_318_U86); 
assign P3_U7234 = ~(P3_SUB_320_U78 & P3_U4319); 
assign P3_U7241 = ~(P3_U2403 & P3_ADD_318_U85); 
assign P3_U7242 = ~(P3_SUB_320_U9 & P3_U4319); 
assign P3_U7249 = ~(P3_U2403 & P3_ADD_318_U84); 
assign P3_U7250 = ~(P3_SUB_320_U76 & P3_U4319); 
assign P3_U7257 = ~(P3_U2403 & P3_ADD_318_U83); 
assign P3_U7258 = ~(P3_SUB_320_U10 & P3_U4319); 
assign P3_U7265 = ~(P3_U2403 & P3_ADD_318_U82); 
assign P3_U7266 = ~(P3_SUB_320_U74 & P3_U4319); 
assign P3_U7273 = ~(P3_U2403 & P3_ADD_318_U81); 
assign P3_U7274 = ~(P3_SUB_320_U11 & P3_U4319); 
assign P3_U7281 = ~(P3_U2403 & P3_ADD_318_U80); 
assign P3_U7282 = ~(P3_SUB_320_U70 & P3_U4319); 
assign P3_U7289 = ~(P3_U2403 & P3_ADD_318_U79); 
assign P3_U7290 = ~(P3_SUB_320_U12 & P3_U4319); 
assign P3_U7297 = ~(P3_U2403 & P3_ADD_318_U78); 
assign P3_U7298 = ~(P3_SUB_320_U68 & P3_U4319); 
assign P3_U7305 = ~(P3_U2403 & P3_ADD_318_U77); 
assign P3_U7306 = ~(P3_SUB_320_U13 & P3_U4319); 
assign P3_U7313 = ~(P3_U2403 & P3_ADD_318_U76); 
assign P3_U7314 = ~(P3_SUB_320_U66 & P3_U4319); 
assign P3_U7321 = ~(P3_U2403 & P3_ADD_318_U75); 
assign P3_U7322 = ~(P3_SUB_320_U14 & P3_U4319); 
assign P3_U7329 = ~(P3_U2403 & P3_ADD_318_U74); 
assign P3_U7330 = ~(P3_SUB_320_U64 & P3_U4319); 
assign P3_U7337 = ~(P3_U2403 & P3_ADD_318_U73); 
assign P3_U7338 = ~(P3_SUB_320_U15 & P3_U4319); 
assign P3_U7345 = ~(P3_U2403 & P3_ADD_318_U72); 
assign P3_U7346 = ~(P3_SUB_320_U16 & P3_U4319); 
assign P3_U7353 = ~(P3_U2403 & P3_ADD_318_U70); 
assign P3_U7354 = ~(P3_SUB_320_U62 & P3_U4319); 
assign P3_U7362 = ~(P3_U2403 & P3_ADD_318_U69); 
assign P2_U2866 = ~(P2_U6535 & P2_U6536 & P2_U6534); 
assign P2_U3597 = ~(P2_U8086 & P2_U8085); 
assign P2_U3598 = ~(P2_U8089 & P2_U8088); 
assign P2_U4087 = P2_U4088 & P2_U6615; 
assign P2_U4091 = P2_U4092 & P2_U6624; 
assign P2_U4124 = P2_U4121 & P2_U6701 & P2_U6702 & P2_U6700 & P2_U6704; 
assign P2_U4128 = P2_U4125 & P2_U6709 & P2_U6710 & P2_U6708 & P2_U6712; 
assign P2_U4132 = P2_U4129 & P2_U6717 & P2_U6718 & P2_U6716 & P2_U6720; 
assign P2_U4136 = P2_U4133 & P2_U6725 & P2_U6726 & P2_U6724 & P2_U6728; 
assign P2_U4140 = P2_U4137 & P2_U6733 & P2_U6734 & P2_U6732 & P2_U6736; 
assign P2_U4143 = P2_U6739 & P2_U6741 & P2_U6742 & P2_U6740 & P2_U6744; 
assign P2_U4146 = P2_U6747 & P2_U6749 & P2_U6750 & P2_U6748 & P2_U6752; 
assign P2_U6388 = ~(P2_ADD_391_1196_U7 & P2_U2397); 
assign P2_U6552 = ~(P2_R2182_U79 & P2_U2393); 
assign P2_U6578 = ~(P2_U2383 & P2_PHYADDRPOINTER_REG_0__SCAN_IN); 
assign P2_U6587 = ~(P2_U2383 & P2_R2337_U4); 
assign P2_U6596 = ~(P2_U2383 & P2_R2337_U70); 
assign P2_U6605 = ~(P2_U2383 & P2_R2337_U67); 
assign P2_U6614 = ~(P2_U2383 & P2_R2337_U66); 
assign P2_U6623 = ~(P2_U2383 & P2_R2337_U65); 
assign P2_U6631 = ~(P2_U2383 & P2_R2337_U64); 
assign P2_U6639 = ~(P2_U2383 & P2_R2337_U63); 
assign P2_U6647 = ~(P2_U2383 & P2_R2337_U62); 
assign P2_U6655 = ~(P2_U2383 & P2_R2337_U61); 
assign P2_U6663 = ~(P2_U2383 & P2_R2337_U90); 
assign P2_U6671 = ~(P2_U2383 & P2_R2337_U89); 
assign P2_U6679 = ~(P2_U2383 & P2_R2337_U88); 
assign P2_U6687 = ~(P2_U2383 & P2_R2337_U87); 
assign P2_U6695 = ~(P2_U2383 & P2_R2337_U86); 
assign P2_U6703 = ~(P2_U2383 & P2_R2337_U85); 
assign P2_U6711 = ~(P2_U2383 & P2_R2337_U84); 
assign P2_U6719 = ~(P2_U2383 & P2_R2337_U83); 
assign P2_U6727 = ~(P2_U2383 & P2_R2337_U82); 
assign P2_U6735 = ~(P2_U2383 & P2_R2337_U81); 
assign P2_U6743 = ~(P2_U2383 & P2_R2337_U80); 
assign P2_U6751 = ~(P2_U2383 & P2_R2337_U79); 
assign P2_U6759 = ~(P2_U2383 & P2_R2337_U78); 
assign P2_U6767 = ~(P2_U2383 & P2_R2337_U77); 
assign P2_U6775 = ~(P2_U2383 & P2_R2337_U76); 
assign P2_U6783 = ~(P2_U2383 & P2_R2337_U75); 
assign P2_U6791 = ~(P2_U2383 & P2_R2337_U74); 
assign P2_U6799 = ~(P2_U2383 & P2_R2337_U73); 
assign P2_U6807 = ~(P2_U2383 & P2_R2337_U72); 
assign P2_U6815 = ~(P2_U2383 & P2_R2337_U71); 
assign P2_U6823 = ~(P2_U2383 & P2_R2337_U69); 
assign P2_U6831 = ~(P2_U2383 & P2_R2337_U68); 
assign P1_U2429 = P1_U6366 & P1_U3431; 
assign P1_U2846 = ~(P1_U6344 & P1_U6345 & P1_U6343); 
assign P1_U2878 = ~(P1_U6243 & P1_U6242 & P1_U6245 & P1_U6244); 
assign P1_U2973 = ~(P1_U5931 & P1_U5929 & P1_U5933 & P1_U5930 & P1_U5932); 
assign P1_U2974 = ~(P1_U5926 & P1_U5924 & P1_U5928 & P1_U5925 & P1_U5927); 
assign P1_U2975 = ~(P1_U5921 & P1_U5919 & P1_U5923 & P1_U5920 & P1_U5922); 
assign P1_U2977 = ~(P1_U5911 & P1_U5909 & P1_U5913 & P1_U5910 & P1_U5912); 
assign P1_U2978 = ~(P1_U5906 & P1_U5904 & P1_U5908 & P1_U5905 & P1_U5907); 
assign P1_U2979 = ~(P1_U5901 & P1_U5899 & P1_U5903 & P1_U5900 & P1_U5902); 
assign P1_U3000 = ~(P1_U3861 & P1_U3859 & P1_U5787 & P1_U5789); 
assign P1_U3003 = ~(P1_U3852 & P1_U3850 & P1_U5766 & P1_U5768); 
assign P1_U3004 = ~(P1_U3849 & P1_U3847 & P1_U5759 & P1_U5761); 
assign P1_U3005 = ~(P1_U3846 & P1_U3844 & P1_U5752 & P1_U5754); 
assign P1_U3006 = ~(P1_U3843 & P1_U3841 & P1_U5745 & P1_U5747); 
assign P1_U3007 = ~(P1_U3840 & P1_U3838 & P1_U5738 & P1_U5740); 
assign P1_U3009 = ~(P1_U3834 & P1_U3832 & P1_U5724 & P1_U5726); 
assign P1_U3010 = ~(P1_U3831 & P1_U3829 & P1_U5717 & P1_U5719); 
assign P1_U3011 = ~(P1_U3828 & P1_U3826 & P1_U5710 & P1_U5712); 
assign P1_U6374 = ~(P1_U2366 & P1_PHYADDRPOINTER_REG_0__SCAN_IN); 
assign P1_U6382 = ~(P1_U2366 & P1_R2337_U4); 
assign P1_U6390 = ~(P1_U2366 & P1_R2337_U71); 
assign P1_U6398 = ~(P1_U2366 & P1_R2337_U68); 
assign P1_U6406 = ~(P1_U2366 & P1_R2337_U67); 
assign P1_U6414 = ~(P1_U2366 & P1_R2337_U66); 
assign P1_U6421 = ~(P1_U2366 & P1_R2337_U65); 
assign P1_U6428 = ~(P1_U2366 & P1_R2337_U64); 
assign P1_U6435 = ~(P1_U2366 & P1_R2337_U63); 
assign P1_U6442 = ~(P1_U2366 & P1_R2337_U62); 
assign P1_U6449 = ~(P1_U2366 & P1_R2337_U91); 
assign P1_U6456 = ~(P1_U2366 & P1_R2337_U90); 
assign P1_U6463 = ~(P1_U2366 & P1_R2337_U89); 
assign P1_U6470 = ~(P1_U2366 & P1_R2337_U88); 
assign P1_U6477 = ~(P1_U2366 & P1_R2337_U87); 
assign P1_U6484 = ~(P1_U2366 & P1_R2337_U86); 
assign P1_U6491 = ~(P1_U2366 & P1_R2337_U85); 
assign P1_U6498 = ~(P1_U2366 & P1_R2337_U84); 
assign P1_U6505 = ~(P1_U2366 & P1_R2337_U83); 
assign P1_U6512 = ~(P1_U2366 & P1_R2337_U82); 
assign P1_U6519 = ~(P1_U2366 & P1_R2337_U81); 
assign P1_U6526 = ~(P1_U2366 & P1_R2337_U80); 
assign P1_U6533 = ~(P1_U2366 & P1_R2337_U79); 
assign P1_U6540 = ~(P1_U2366 & P1_R2337_U78); 
assign P1_U6547 = ~(P1_U2366 & P1_R2337_U77); 
assign P1_U6554 = ~(P1_U2366 & P1_R2337_U76); 
assign P1_U6561 = ~(P1_U2366 & P1_R2337_U75); 
assign P1_U6568 = ~(P1_U2366 & P1_R2337_U74); 
assign P1_U6575 = ~(P1_U2366 & P1_R2337_U73); 
assign P1_U6582 = ~(P1_U2366 & P1_R2337_U72); 
assign P1_U6589 = ~(P1_U2366 & P1_R2337_U70); 
assign P1_U6596 = ~(P1_U2366 & P1_R2337_U69); 
assign P3_SUB_320_U51 = ~(P3_SUB_320_U137 & P3_SUB_320_U136); 
assign P2_R2099_U81 = ~(P2_R2099_U194 & P2_R2099_U193); 
assign P2_R2099_U138 = ~P2_R2099_U51; 
assign P2_R2099_U191 = ~(P2_U2724 & P2_R2099_U51); 
assign P2_ADD_391_1196_U76 = ~P2_R2182_U79; 
assign P2_ADD_391_1196_U106 = ~(P2_ADD_391_1196_U453 & P2_ADD_391_1196_U452); 
assign P2_ADD_391_1196_U129 = P2_ADD_391_1196_U373 & P2_ADD_391_1196_U372; 
assign P2_ADD_391_1196_U231 = ~P2_ADD_391_1196_U150; 
assign P2_ADD_391_1196_U233 = ~(P2_ADD_391_1196_U232 & P2_ADD_391_1196_U150); 
assign P2_ADD_391_1196_U272 = P2_R2182_U79 | P2_R2096_U80; 
assign P2_ADD_391_1196_U274 = ~(P2_R2096_U80 & P2_R2182_U79); 
assign P2_ADD_391_1196_U366 = ~(P2_R2182_U79 & P2_ADD_391_1196_U77); 
assign P2_ADD_391_1196_U368 = ~(P2_R2182_U79 & P2_ADD_391_1196_U77); 
assign P2_ADD_391_1196_U376 = ~(P2_ADD_391_1196_U375 & P2_ADD_391_1196_U374); 
assign P2_ADD_391_1196_U445 = ~(P2_ADD_391_1196_U149 & P2_ADD_391_1196_U150); 
assign P2_R2182_U66 = ~(P2_R2182_U177 & P2_R2182_U176); 
assign P2_R2182_U237 = ~(P2_R2182_U174 & P2_R2182_U235); 
assign P2_R1957_U50 = ~(P2_R1957_U137 & P2_R1957_U136); 
assign P2_R2278_U139 = P2_R2278_U397 & P2_R2278_U138; 
assign P2_R2278_U141 = P2_R2278_U4 & P2_R2278_U142; 
assign P2_R2278_U196 = ~(P2_R2278_U124 & P2_R2278_U323); 
assign P2_R2278_U198 = ~(P2_R2278_U55 & P2_R2278_U246); 
assign P2_R2278_U400 = ~(P2_R2278_U4 & P2_R2278_U79 & P2_R2278_U80); 
assign P2_R2278_U401 = ~(P2_U2791 & P2_R2278_U397 & P2_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P2_R2278_U546 = ~(P2_R2278_U244 & P2_R2278_U544); 
assign P2_R2278_U553 = ~(P2_R2278_U241 & P2_R2278_U551); 
assign P1_R2358_U91 = ~(P1_R2358_U581 & P1_R2358_U580); 
assign P1_R2358_U177 = ~P1_U2651; 
assign P1_R2358_U179 = ~(P1_U2621 & P1_R2358_U564); 
assign P1_R2358_U183 = ~(P1_R2358_U297 & P1_R2358_U298); 
assign P1_R2358_U555 = ~(P1_U2651 & P1_R2358_U23); 
assign P1_R2358_U556 = ~(P1_U2352 & P1_R2358_U178); 
assign P1_R2358_U560 = ~(P1_U2651 & P1_R2358_U23); 
assign P1_R2358_U578 = ~(P1_R2358_U184 & P1_R2358_U337); 
assign P1_R2358_U579 = ~(P1_R2358_U88 & P1_R2358_U384); 
assign P3_U2833 = ~(P3_U6351 & P3_U6349 & P3_U6350); 
assign P3_U3941 = P3_U6380 & P3_U6379; 
assign P3_U3944 = P3_U6383 & P3_U6382 & P3_U3943; 
assign P3_U3947 = P3_U6391 & P3_U6390; 
assign P3_U3949 = P3_U6394 & P3_U6393; 
assign P3_U4033 = P3_U4034 & P3_U7104; 
assign P3_U4037 = P3_U4038 & P3_U7114; 
assign P3_U4041 = P3_U4042 & P3_U7124; 
assign P3_U4045 = P3_U4046 & P3_U7134; 
assign P3_U4049 = P3_U4050 & P3_U7144; 
assign P3_U4051 = P3_U4048 & P3_U7139 & P3_U4047 & P3_U7142 & P3_U7143; 
assign P3_U4054 = P3_U4055 & P3_U7154; 
assign P3_U4056 = P3_U4053 & P3_U7149 & P3_U4052 & P3_U7152 & P3_U7153; 
assign P3_U4058 = P3_U4059 & P3_U7161; 
assign P3_U4061 = P3_U4062 & P3_U7169; 
assign P3_U4064 = P3_U4065 & P3_U7177; 
assign P3_U4067 = P3_U4068 & P3_U7185; 
assign P3_U4070 = P3_U4071 & P3_U7193; 
assign P3_U4073 = P3_U4074 & P3_U7201; 
assign P3_U4076 = P3_U4077 & P3_U7209; 
assign P3_U4079 = P3_U4080 & P3_U7217; 
assign P3_U4082 = P3_U4083 & P3_U7225; 
assign P3_U4085 = P3_U4086 & P3_U7233; 
assign P3_U4088 = P3_U4089 & P3_U7241; 
assign P3_U4091 = P3_U4092 & P3_U7249; 
assign P3_U4094 = P3_U4095 & P3_U7257; 
assign P3_U4097 = P3_U4098 & P3_U7265; 
assign P3_U4100 = P3_U4101 & P3_U7273; 
assign P3_U4103 = P3_U4104 & P3_U7281; 
assign P3_U4106 = P3_U4107 & P3_U7289; 
assign P3_U4109 = P3_U4110 & P3_U7297; 
assign P3_U4112 = P3_U4113 & P3_U7305; 
assign P3_U4115 = P3_U4116 & P3_U7313; 
assign P3_U4118 = P3_U4119 & P3_U7321; 
assign P3_U4121 = P3_U4122 & P3_U7329; 
assign P3_U4124 = P3_U4125 & P3_U7337; 
assign P3_U4127 = P3_U4128 & P3_U7345; 
assign P3_U4130 = P3_U4131 & P3_U7353; 
assign P3_U4134 = P3_U7362 & P3_U3259; 
assign P3_U6372 = ~(P3_U3930 & P3_U6354 & P3_U3931 & P3_U3933 & P3_U3938); 
assign P3_U7363 = ~P3_U7362; 
assign P2_U2904 = ~(P2_U6390 & P2_U6387 & P2_U6389 & P2_U6388); 
assign P2_U4072 = P2_U4073 & P2_U6578; 
assign P2_U4076 = P2_U4077 & P2_U6587; 
assign P2_U4080 = P2_U4081 & P2_U6596; 
assign P2_U4084 = P2_U4085 & P2_U6605; 
assign P2_U4089 = P2_U6612 & P2_U6611 & P2_U4086 & P2_U6613 & P2_U6614; 
assign P2_U4093 = P2_U6621 & P2_U6620 & P2_U4090 & P2_U6622 & P2_U6623; 
assign P2_U4095 = P2_U4096 & P2_U6631; 
assign P2_U4098 = P2_U4099 & P2_U6639; 
assign P2_U4101 = P2_U4102 & P2_U6647; 
assign P2_U4104 = P2_U4105 & P2_U6655; 
assign P2_U4107 = P2_U4108 & P2_U6663; 
assign P2_U4110 = P2_U4111 & P2_U6671; 
assign P2_U4113 = P2_U4114 & P2_U6679; 
assign P2_U4116 = P2_U4117 & P2_U6687; 
assign P2_U4119 = P2_U4120 & P2_U6695; 
assign P2_U4122 = P2_U4123 & P2_U6703; 
assign P2_U4126 = P2_U4127 & P2_U6711; 
assign P2_U4130 = P2_U4131 & P2_U6719; 
assign P2_U4134 = P2_U4135 & P2_U6727; 
assign P2_U4138 = P2_U4139 & P2_U6735; 
assign P2_U4141 = P2_U4142 & P2_U6743; 
assign P2_U4144 = P2_U4145 & P2_U6751; 
assign P2_U4148 = P2_U4147 & P2_U6759 & P2_U6760; 
assign P2_U4150 = P2_U4151 & P2_U6767; 
assign P2_U4153 = P2_U4154 & P2_U6775; 
assign P2_U4156 = P2_U4155 & P2_U6783 & P2_U6784; 
assign P2_U4158 = P2_U4157 & P2_U6791 & P2_U6792; 
assign P2_U4160 = P2_U4159 & P2_U6799 & P2_U6800; 
assign P2_U4162 = P2_U4161 & P2_U6807 & P2_U6808; 
assign P2_U4164 = P2_U4163 & P2_U6815 & P2_U6816; 
assign P2_U4166 = P2_U4165 & P2_U6823 & P2_U6824; 
assign P2_U5620 = ~(P2_U3598 & P2_U3597 & P2_STATE2_REG_1__SCAN_IN); 
assign P2_U6393 = ~(P2_ADD_391_1196_U106 & P2_U2397); 
assign P2_U6538 = ~(P2_U2379 & P2_R2099_U81); 
assign P2_U6758 = ~(P2_U2392 & P2_R2099_U81); 
assign P2_U6832 = ~(P2_R1957_U50 & P2_U2382); 
assign P2_U8087 = ~P2_U3597; 
assign P2_U8090 = ~P2_U3598; 
assign P2_U8282 = ~(P2_U3598 & P2_U3597 & P2_FLUSH_REG_SCAN_IN); 
assign P1_U3895 = P1_U6405 & P1_U6404 & P1_U6407 & P1_U6406; 
assign P1_U3899 = P1_U6422 & P1_U6419 & P1_U6421; 
assign P1_U3901 = P1_U6429 & P1_U6426 & P1_U6428; 
assign P1_U3903 = P1_U6436 & P1_U6433 & P1_U6435; 
assign P1_U3905 = P1_U6443 & P1_U6440 & P1_U6442; 
assign P1_U3907 = P1_U6450 & P1_U6447 & P1_U6449; 
assign P1_U3909 = P1_U6457 & P1_U6454 & P1_U6456; 
assign P1_U3911 = P1_U6464 & P1_U6461 & P1_U6463; 
assign P1_U3913 = P1_U6471 & P1_U6468 & P1_U6470; 
assign P1_U3915 = P1_U6478 & P1_U6475 & P1_U6477; 
assign P1_U3917 = P1_U6485 & P1_U6482 & P1_U6484; 
assign P1_U3919 = P1_U6492 & P1_U6489 & P1_U6491; 
assign P1_U3921 = P1_U6499 & P1_U6496 & P1_U6498; 
assign P1_U3923 = P1_U6506 & P1_U6503 & P1_U6505; 
assign P1_U3925 = P1_U6513 & P1_U6510 & P1_U6512; 
assign P1_U3927 = P1_U6519 & P1_U6520; 
assign P1_U3929 = P1_U6526 & P1_U6527; 
assign P1_U3931 = P1_U6533 & P1_U6534; 
assign P1_U3933 = P1_U6540 & P1_U6541; 
assign P1_U3935 = P1_U6547 & P1_U6548; 
assign P1_U3937 = P1_U6554 & P1_U6555; 
assign P1_U3939 = P1_U6561 & P1_U6562; 
assign P1_U3941 = P1_U6568 & P1_U6569; 
assign P1_U3943 = P1_U6575 & P1_U6576; 
assign P1_U3945 = P1_U6582 & P1_U6583; 
assign P1_U3947 = P1_U6589 & P1_U6590; 
assign P1_U3949 = P1_U6596 & P1_U6597; 
assign P1_U5937 = ~(P1_R2358_U91 & P1_U2364); 
assign P1_U6248 = ~(P1_U2386 & P1_R2358_U91); 
assign P1_U6346 = ~(P1_U2383 & P1_R2358_U91); 
assign P1_U6371 = ~(P1_U2429 & P1_R2358_U76); 
assign P1_U6379 = ~(P1_U2429 & P1_R2358_U107); 
assign P1_U6387 = ~(P1_U2429 & P1_R2358_U18); 
assign P1_U6395 = ~(P1_U2429 & P1_R2358_U19); 
assign P1_U6403 = ~(P1_U2429 & P1_R2358_U84); 
assign P1_U6411 = ~(P1_U2429 & P1_R2358_U82); 
assign P1_U6567 = ~(P1_U2367 & P1_R2358_U91); 
assign P2_R2099_U53 = ~(P2_U2724 & P2_R2099_U138); 
assign P2_R2099_U192 = ~(P2_R2099_U138 & P2_R2099_U52); 
assign P2_ADD_391_1196_U148 = ~(P2_ADD_391_1196_U234 & P2_ADD_391_1196_U233); 
assign P2_ADD_391_1196_U365 = ~(P2_R2096_U80 & P2_ADD_391_1196_U76); 
assign P2_ADD_391_1196_U367 = ~(P2_R2096_U80 & P2_ADD_391_1196_U76); 
assign P2_ADD_391_1196_U446 = ~(P2_ADD_391_1196_U231 & P2_ADD_391_1196_U444); 
assign P2_R2182_U78 = ~(P2_R2182_U237 & P2_R2182_U236); 
assign P2_R2182_U178 = ~P2_R2182_U66; 
assign P2_R2182_U180 = ~(P2_R2182_U179 & P2_R2182_U66); 
assign P2_R2182_U229 = ~(P2_R2182_U109 & P2_R2182_U66); 
assign P2_R2278_U110 = ~(P2_R2278_U546 & P2_R2278_U545); 
assign P2_R2278_U111 = ~(P2_R2278_U553 & P2_R2278_U552); 
assign P2_R2278_U161 = P2_R2278_U401 & P2_R2278_U400; 
assign P2_R2278_U248 = ~P2_R2278_U198; 
assign P2_R2278_U251 = ~P2_R2278_U196; 
assign P2_R2278_U253 = ~(P2_R2278_U252 & P2_R2278_U196); 
assign P2_R2278_U325 = ~(P2_R2278_U125 & P2_R2278_U196); 
assign P2_R2278_U531 = ~(P2_R2278_U195 & P2_R2278_U196); 
assign P2_R2278_U538 = ~(P2_R2278_U197 & P2_R2278_U198); 
assign P1_R2358_U75 = ~(P1_R2358_U557 & P1_R2358_U556); 
assign P1_R2358_U86 = P1_R2358_U179 & P1_R2358_U300; 
assign P1_R2358_U89 = ~(P1_R2358_U579 & P1_R2358_U578); 
assign P1_R2358_U299 = ~P1_R2358_U183; 
assign P1_R2358_U301 = ~P1_R2358_U179; 
assign P1_R2358_U302 = ~(P1_R2358_U300 & P1_R2358_U183); 
assign P1_R2358_U336 = ~(P1_R2358_U179 & P1_R2358_U300); 
assign P1_R2358_U554 = ~(P1_U2352 & P1_R2358_U177); 
assign P1_R2358_U559 = ~(P1_U2352 & P1_R2358_U177); 
assign P3_U2641 = ~(P3_U7352 & P3_U7351 & P3_U4129 & P3_U7354 & P3_U4130); 
assign P3_U2642 = ~(P3_U7344 & P3_U7343 & P3_U4126 & P3_U7346 & P3_U4127); 
assign P3_U2643 = ~(P3_U7336 & P3_U7335 & P3_U4123 & P3_U7338 & P3_U4124); 
assign P3_U2644 = ~(P3_U7328 & P3_U7327 & P3_U4120 & P3_U7330 & P3_U4121); 
assign P3_U2645 = ~(P3_U7320 & P3_U7319 & P3_U4117 & P3_U7322 & P3_U4118); 
assign P3_U2646 = ~(P3_U7312 & P3_U7311 & P3_U4114 & P3_U7314 & P3_U4115); 
assign P3_U2647 = ~(P3_U7304 & P3_U7303 & P3_U4111 & P3_U7306 & P3_U4112); 
assign P3_U2648 = ~(P3_U7296 & P3_U7295 & P3_U4108 & P3_U7298 & P3_U4109); 
assign P3_U2649 = ~(P3_U7288 & P3_U7287 & P3_U4105 & P3_U7290 & P3_U4106); 
assign P3_U2650 = ~(P3_U7280 & P3_U7279 & P3_U4102 & P3_U7282 & P3_U4103); 
assign P3_U2651 = ~(P3_U7272 & P3_U7271 & P3_U4099 & P3_U7274 & P3_U4100); 
assign P3_U2652 = ~(P3_U7264 & P3_U7263 & P3_U4096 & P3_U7266 & P3_U4097); 
assign P3_U2653 = ~(P3_U7256 & P3_U7255 & P3_U4093 & P3_U7258 & P3_U4094); 
assign P3_U2654 = ~(P3_U7248 & P3_U7247 & P3_U4090 & P3_U7250 & P3_U4091); 
assign P3_U2655 = ~(P3_U7240 & P3_U7239 & P3_U4087 & P3_U7242 & P3_U4088); 
assign P3_U2656 = ~(P3_U7232 & P3_U7231 & P3_U4084 & P3_U7234 & P3_U4085); 
assign P3_U2657 = ~(P3_U7224 & P3_U7223 & P3_U4081 & P3_U7226 & P3_U4082); 
assign P3_U2658 = ~(P3_U7216 & P3_U7215 & P3_U4078 & P3_U7218 & P3_U4079); 
assign P3_U2659 = ~(P3_U7208 & P3_U7207 & P3_U4075 & P3_U7210 & P3_U4076); 
assign P3_U2660 = ~(P3_U7200 & P3_U7199 & P3_U4072 & P3_U7202 & P3_U4073); 
assign P3_U2661 = ~(P3_U7192 & P3_U7191 & P3_U4069 & P3_U7194 & P3_U4070); 
assign P3_U2662 = ~(P3_U7184 & P3_U7183 & P3_U4066 & P3_U7186 & P3_U4067); 
assign P3_U2663 = ~(P3_U7176 & P3_U7175 & P3_U4063 & P3_U7178 & P3_U4064); 
assign P3_U2664 = ~(P3_U7168 & P3_U7167 & P3_U4060 & P3_U7170 & P3_U4061); 
assign P3_U2665 = ~(P3_U7160 & P3_U7159 & P3_U4057 & P3_U7162 & P3_U4058); 
assign P3_U2666 = ~(P3_U4056 & P3_U4054); 
assign P3_U2667 = ~(P3_U4051 & P3_U4049); 
assign P3_U2668 = ~(P3_U7129 & P3_U4043 & P3_U7132 & P3_U7133 & P3_U4045); 
assign P3_U2669 = ~(P3_U7119 & P3_U4039 & P3_U7122 & P3_U7123 & P3_U4041); 
assign P3_U2670 = ~(P3_U7109 & P3_U4035 & P3_U7112 & P3_U7113 & P3_U4037); 
assign P3_U2671 = ~(P3_U7099 & P3_U4031 & P3_U7102 & P3_U7103 & P3_U4033); 
assign P3_U3942 = P3_U3941 & P3_U6381; 
assign P3_U3948 = P3_U3946 & P3_U6392 & P3_U3947; 
assign P3_U4135 = ~(P3_SUB_320_U51 | P3_U7363); 
assign P3_U6374 = ~(P3_U4318 & P3_U6372); 
assign P3_U7907 = ~(P3_U4134 & P3_U2603); 
assign P2_U2833 = ~(P2_U6755 & P2_U6757 & P2_U6758 & P2_U6756 & P2_U4148); 
assign P2_U2834 = ~(P2_U4146 & P2_U4144); 
assign P2_U2835 = ~(P2_U4143 & P2_U4141); 
assign P2_U2836 = ~(P2_U4140 & P2_U4138); 
assign P2_U2837 = ~(P2_U4136 & P2_U4134); 
assign P2_U2838 = ~(P2_U4132 & P2_U4130); 
assign P2_U2839 = ~(P2_U4128 & P2_U4126); 
assign P2_U2840 = ~(P2_U4124 & P2_U4122); 
assign P2_U2841 = ~(P2_U6693 & P2_U4118 & P2_U6692 & P2_U6696 & P2_U4119); 
assign P2_U2842 = ~(P2_U6685 & P2_U4115 & P2_U6684 & P2_U6688 & P2_U4116); 
assign P2_U2843 = ~(P2_U6677 & P2_U4112 & P2_U6676 & P2_U6680 & P2_U4113); 
assign P2_U2844 = ~(P2_U6670 & P2_U6669 & P2_U4109 & P2_U6672 & P2_U4110); 
assign P2_U2845 = ~(P2_U6662 & P2_U6661 & P2_U4106 & P2_U6664 & P2_U4107); 
assign P2_U2846 = ~(P2_U6654 & P2_U6653 & P2_U4103 & P2_U6656 & P2_U4104); 
assign P2_U2847 = ~(P2_U6646 & P2_U6645 & P2_U4100 & P2_U6648 & P2_U4101); 
assign P2_U2848 = ~(P2_U6638 & P2_U6637 & P2_U4097 & P2_U6640 & P2_U4098); 
assign P2_U2849 = ~(P2_U6630 & P2_U6629 & P2_U4094 & P2_U6632 & P2_U4095); 
assign P2_U2850 = ~(P2_U4093 & P2_U4091); 
assign P2_U2851 = ~(P2_U4089 & P2_U4087); 
assign P2_U2852 = ~(P2_U6602 & P2_U4082 & P2_U6606 & P2_U4084); 
assign P2_U2853 = ~(P2_U6593 & P2_U4078 & P2_U6597 & P2_U4080); 
assign P2_U2854 = ~(P2_U6584 & P2_U4074 & P2_U6588 & P2_U4076); 
assign P2_U2855 = ~(P2_U6575 & P2_U4070 & P2_U6579 & P2_U4072); 
assign P2_U2865 = ~(P2_U6538 & P2_U6539 & P2_U6537); 
assign P2_U2903 = ~(P2_U6392 & P2_U6391 & P2_U6395 & P2_U6394 & P2_U6393); 
assign P2_U3613 = ~(P2_U8282 & P2_U8281); 
assign P2_U4168 = P2_U4167 & P2_U6831 & P2_U6832; 
assign P2_U5623 = ~(P2_U5621 & P2_U5622 & P2_U5620); 
assign P2_U5630 = ~(P2_U8090 & P2_U3597 & P2_STATE2_REG_1__SCAN_IN); 
assign P2_U5640 = ~(P2_U8087 & P2_STATE2_REG_1__SCAN_IN); 
assign P2_U6555 = ~(P2_R2182_U78 & P2_U2393); 
assign P2_U8284 = ~(P2_U3597 & P2_U8090 & P2_FLUSH_REG_SCAN_IN); 
assign P2_U8286 = ~(P2_U8087 & P2_FLUSH_REG_SCAN_IN); 
assign P1_U2813 = ~(P1_U6565 & P1_U3940 & P1_U3941 & P1_U6563 & P1_U6567); 
assign P1_U2814 = ~(P1_U6558 & P1_U3938 & P1_U3939 & P1_U6556 & P1_U6560); 
assign P1_U2815 = ~(P1_U6551 & P1_U3936 & P1_U3937 & P1_U6549 & P1_U6553); 
assign P1_U2816 = ~(P1_U6544 & P1_U3934 & P1_U3935 & P1_U6542 & P1_U6546); 
assign P1_U2817 = ~(P1_U6537 & P1_U3932 & P1_U3933 & P1_U6535 & P1_U6539); 
assign P1_U2818 = ~(P1_U6530 & P1_U3930 & P1_U3931 & P1_U6528 & P1_U6532); 
assign P1_U2819 = ~(P1_U6523 & P1_U3928 & P1_U3929 & P1_U6521 & P1_U6525); 
assign P1_U2820 = ~(P1_U6516 & P1_U3926 & P1_U3927 & P1_U6514 & P1_U6518); 
assign P1_U2821 = ~(P1_U3924 & P1_U6509 & P1_U3925 & P1_U6507 & P1_U6511); 
assign P1_U2822 = ~(P1_U3922 & P1_U6502 & P1_U3923 & P1_U6500 & P1_U6504); 
assign P1_U2823 = ~(P1_U3920 & P1_U6495 & P1_U3921 & P1_U6493 & P1_U6497); 
assign P1_U2824 = ~(P1_U6488 & P1_U6487 & P1_U3919 & P1_U3918 & P1_U6490); 
assign P1_U2825 = ~(P1_U6481 & P1_U6480 & P1_U3917 & P1_U3916 & P1_U6483); 
assign P1_U2826 = ~(P1_U3915 & P1_U6474 & P1_U3914 & P1_U6473 & P1_U6476); 
assign P1_U2827 = ~(P1_U3913 & P1_U6467 & P1_U3912 & P1_U6466 & P1_U6469); 
assign P1_U2828 = ~(P1_U3911 & P1_U6460 & P1_U3910 & P1_U6459 & P1_U6462); 
assign P1_U2829 = ~(P1_U3909 & P1_U6453 & P1_U3908 & P1_U6452 & P1_U6455); 
assign P1_U2830 = ~(P1_U3907 & P1_U6446 & P1_U3906 & P1_U6445 & P1_U6448); 
assign P1_U2831 = ~(P1_U3905 & P1_U6439 & P1_U3904 & P1_U6438 & P1_U6441); 
assign P1_U2832 = ~(P1_U3903 & P1_U6432 & P1_U3902 & P1_U6431 & P1_U6434); 
assign P1_U2833 = ~(P1_U3901 & P1_U6425 & P1_U3900 & P1_U6424 & P1_U6427); 
assign P1_U2834 = ~(P1_U3899 & P1_U6418 & P1_U3898 & P1_U6417 & P1_U6420); 
assign P1_U2836 = ~(P1_U3894 & P1_U6401 & P1_U3895 & P1_U6403 & P1_U6402); 
assign P1_U2845 = ~(P1_U6347 & P1_U6348 & P1_U6346); 
assign P1_U2877 = ~(P1_U6247 & P1_U6246 & P1_U6249 & P1_U6248); 
assign P1_U2972 = ~(P1_U5936 & P1_U5934 & P1_U5938 & P1_U5935 & P1_U5937); 
assign P1_U3890 = P1_U6373 & P1_U6372 & P1_U6375 & P1_U6374 & P1_U6371; 
assign P1_U3891 = P1_U6381 & P1_U6380 & P1_U6383 & P1_U6382 & P1_U6379; 
assign P1_U3892 = P1_U6389 & P1_U6388 & P1_U6391 & P1_U6390 & P1_U6387; 
assign P1_U3893 = P1_U6397 & P1_U6396 & P1_U6399 & P1_U6398 & P1_U6395; 
assign P1_U3897 = P1_U6413 & P1_U6412 & P1_U6415 & P1_U6414 & P1_U6411; 
assign P1_U5942 = ~(P1_R2358_U89 & P1_U2364); 
assign P1_U6252 = ~(P1_U2386 & P1_R2358_U89); 
assign P1_U6349 = ~(P1_U2383 & P1_R2358_U89); 
assign P1_U6574 = ~(P1_U2367 & P1_R2358_U89); 
assign P2_R2099_U80 = ~(P2_R2099_U192 & P2_R2099_U191); 
assign P2_R2099_U139 = ~P2_R2099_U53; 
assign P2_R2099_U189 = ~(P2_U2723 & P2_R2099_U53); 
assign P2_ADD_391_1196_U79 = ~P2_R2182_U78; 
assign P2_ADD_391_1196_U105 = ~(P2_ADD_391_1196_U446 & P2_ADD_391_1196_U445); 
assign P2_ADD_391_1196_U127 = P2_ADD_391_1196_U366 & P2_ADD_391_1196_U365; 
assign P2_ADD_391_1196_U235 = ~P2_ADD_391_1196_U148; 
assign P2_ADD_391_1196_U237 = ~(P2_ADD_391_1196_U236 & P2_ADD_391_1196_U148); 
assign P2_ADD_391_1196_U276 = P2_R2096_U79 | P2_R2182_U78; 
assign P2_ADD_391_1196_U278 = ~(P2_R2182_U78 & P2_R2096_U79); 
assign P2_ADD_391_1196_U358 = ~(P2_R2182_U78 & P2_ADD_391_1196_U78); 
assign P2_ADD_391_1196_U360 = ~(P2_R2182_U78 & P2_ADD_391_1196_U78); 
assign P2_ADD_391_1196_U369 = ~(P2_ADD_391_1196_U368 & P2_ADD_391_1196_U367); 
assign P2_ADD_391_1196_U438 = ~(P2_ADD_391_1196_U147 & P2_ADD_391_1196_U148); 
assign P2_R2182_U182 = ~(P2_R2182_U97 & P2_R2182_U180); 
assign P2_R2182_U184 = ~(P2_R2182_U178 & P2_R2182_U183); 
assign P2_R2182_U230 = ~(P2_R2182_U228 & P2_R2182_U178); 
assign P2_R2278_U192 = ~(P2_R2278_U126 & P2_R2278_U325); 
assign P2_R2278_U194 = ~(P2_R2278_U58 & P2_R2278_U253); 
assign P2_R2278_U532 = ~(P2_R2278_U251 & P2_R2278_U530); 
assign P2_R2278_U539 = ~(P2_R2278_U248 & P2_R2278_U537); 
assign P1_R2358_U13 = P1_R2358_U555 & P1_R2358_U554; 
assign P1_R2358_U182 = ~(P1_R2358_U179 & P1_R2358_U302); 
assign P1_R2358_U304 = ~(P1_U2620 & P1_R2358_U75); 
assign P1_R2358_U558 = ~P1_R2358_U75; 
assign P1_R2358_U561 = ~(P1_R2358_U560 & P1_R2358_U559); 
assign P1_R2358_U570 = ~(P1_R2358_U75 & P1_R2358_U63); 
assign P1_R2358_U572 = ~(P1_R2358_U75 & P1_R2358_U63); 
assign P1_R2358_U576 = ~(P1_R2358_U336 & P1_R2358_U183); 
assign P1_R2358_U577 = ~(P1_R2358_U86 & P1_R2358_U299); 
assign P3_U2832 = ~(P3_U6375 & P3_U6373 & P3_U6374); 
assign P3_U3945 = P3_U3940 & P3_U6378 & P3_U3942 & P3_U3944; 
assign P3_U3950 = P3_U6398 & P3_U6397 & P3_U6395 & P3_U3949 & P3_U3948; 
assign P3_U7357 = ~(P3_U4135 & P3_U2603); 
assign P2_U3614 = ~(P2_U8284 & P2_U8283); 
assign P2_U3615 = ~(P2_U8286 & P2_U8285); 
assign P2_U5633 = ~(P2_U5631 & P2_U5632 & P2_U5630); 
assign P2_U5641 = ~(P2_U5639 & P2_U5638 & P2_U5640); 
assign P2_U6398 = ~(P2_ADD_391_1196_U105 & P2_U2397); 
assign P2_U6541 = ~(P2_U2379 & P2_R2099_U80); 
assign P2_U6766 = ~(P2_U2392 & P2_R2099_U80); 
assign P2_U8094 = ~(P2_U5623 & P2_U4394); 
assign P1_U2812 = ~(P1_U6572 & P1_U3942 & P1_U3943 & P1_U6570 & P1_U6574); 
assign P1_U2835 = ~(P1_U3896 & P1_U6409 & P1_U6410 & P1_U3897); 
assign P1_U2837 = ~(P1_U6393 & P1_U6392 & P1_U6394 & P1_U3893); 
assign P1_U2838 = ~(P1_U6385 & P1_U6384 & P1_U6386 & P1_U3892); 
assign P1_U2839 = ~(P1_U6377 & P1_U6376 & P1_U6378 & P1_U3891); 
assign P1_U2840 = ~(P1_U6369 & P1_U6368 & P1_U6370 & P1_U3890); 
assign P1_U2844 = ~(P1_U6350 & P1_U6351 & P1_U6349); 
assign P1_U2876 = ~(P1_U6251 & P1_U6250 & P1_U6253 & P1_U6252); 
assign P1_U2971 = ~(P1_U5941 & P1_U5939 & P1_U5943 & P1_U5940 & P1_U5942); 
assign P2_R2099_U55 = ~(P2_U2723 & P2_R2099_U139); 
assign P2_R2099_U190 = ~(P2_R2099_U139 & P2_R2099_U54); 
assign P2_ADD_391_1196_U146 = ~(P2_ADD_391_1196_U238 & P2_ADD_391_1196_U237); 
assign P2_ADD_391_1196_U359 = ~(P2_R2096_U79 & P2_ADD_391_1196_U79); 
assign P2_ADD_391_1196_U361 = ~(P2_R2096_U79 & P2_ADD_391_1196_U79); 
assign P2_ADD_391_1196_U439 = ~(P2_ADD_391_1196_U235 & P2_ADD_391_1196_U437); 
assign P2_R2182_U77 = ~(P2_R2182_U230 & P2_R2182_U229); 
assign P2_R2182_U186 = ~(P2_R2182_U98 & P2_R2182_U184); 
assign P2_SUB_589_U9 = ~P2_U3613; 
assign P2_R2278_U108 = ~(P2_R2278_U532 & P2_R2278_U531); 
assign P2_R2278_U109 = ~(P2_R2278_U539 & P2_R2278_U538); 
assign P2_R2278_U255 = ~P2_R2278_U194; 
assign P2_R2278_U258 = ~P2_R2278_U192; 
assign P2_R2278_U260 = ~(P2_R2278_U259 & P2_R2278_U192); 
assign P2_R2278_U327 = ~(P2_R2278_U127 & P2_R2278_U192); 
assign P2_R2278_U517 = ~(P2_R2278_U191 & P2_R2278_U192); 
assign P2_R2278_U524 = ~(P2_R2278_U193 & P2_R2278_U194); 
assign P1_R2358_U87 = ~(P1_R2358_U577 & P1_R2358_U576); 
assign P1_R2358_U135 = P1_R2358_U304 & P1_R2358_U13; 
assign P1_R2358_U303 = ~P1_R2358_U182; 
assign P1_R2358_U305 = ~(P1_R2358_U558 & P1_R2358_U63); 
assign P1_R2358_U567 = ~(P1_R2358_U13 & P1_R2358_U558 & P1_R2358_U63); 
assign P1_R2358_U568 = ~(P1_R2358_U561 & P1_R2358_U75 & P1_U2620); 
assign P1_R2358_U569 = ~(P1_R2358_U558 & P1_U2620); 
assign P1_R2358_U571 = ~(P1_R2358_U558 & P1_U2620); 
assign P3_U2640 = P3_U7357 & P3_U7907; 
assign P3_U6396 = ~(P3_U3950 & P3_U3945); 
assign P2_U2864 = ~(P2_U6541 & P2_U6542 & P2_U6540); 
assign P2_U2902 = ~(P2_U6397 & P2_U6396 & P2_U6400 & P2_U6399 & P2_U6398); 
assign P2_U3599 = ~(P2_U8094 & P2_U8093); 
assign P2_U4149 = P2_U6763 & P2_U6765 & P2_U6766 & P2_U6768 & P2_U4150; 
assign P2_U6558 = ~(P2_R2182_U77 & P2_U2393); 
assign P2_U8102 = ~(P2_U5633 & P2_U4394); 
assign P2_U8104 = ~(P2_U5641 & P2_U4394); 
assign P2_U8430 = ~(P2_SUB_589_U9 & P2_STATE2_REG_1__SCAN_IN); 
assign P1_U5947 = ~(P1_R2358_U87 & P1_U2364); 
assign P1_U6256 = ~(P1_U2386 & P1_R2358_U87); 
assign P1_U6352 = ~(P1_U2383 & P1_R2358_U87); 
assign P1_U6581 = ~(P1_U2367 & P1_R2358_U87); 
assign P2_R2099_U79 = ~(P2_R2099_U190 & P2_R2099_U189); 
assign P2_R2099_U140 = ~P2_R2099_U55; 
assign P2_R2099_U187 = ~(P2_U2722 & P2_R2099_U55); 
assign P2_ADD_391_1196_U81 = ~P2_R2182_U77; 
assign P2_ADD_391_1196_U104 = ~(P2_ADD_391_1196_U439 & P2_ADD_391_1196_U438); 
assign P2_ADD_391_1196_U125 = P2_ADD_391_1196_U359 & P2_ADD_391_1196_U358; 
assign P2_ADD_391_1196_U239 = ~P2_ADD_391_1196_U146; 
assign P2_ADD_391_1196_U241 = ~(P2_ADD_391_1196_U240 & P2_ADD_391_1196_U146); 
assign P2_ADD_391_1196_U280 = P2_R2096_U78 | P2_R2182_U77; 
assign P2_ADD_391_1196_U282 = ~(P2_R2182_U77 & P2_R2096_U78); 
assign P2_ADD_391_1196_U284 = ~(P2_R2182_U77 & P2_R2096_U78); 
assign P2_ADD_391_1196_U286 = P2_R2182_U77 | P2_R2096_U78; 
assign P2_ADD_391_1196_U351 = ~(P2_R2182_U77 & P2_ADD_391_1196_U80); 
assign P2_ADD_391_1196_U353 = ~(P2_R2182_U77 & P2_ADD_391_1196_U80); 
assign P2_ADD_391_1196_U362 = ~(P2_ADD_391_1196_U361 & P2_ADD_391_1196_U360); 
assign P2_ADD_391_1196_U431 = ~(P2_ADD_391_1196_U145 & P2_ADD_391_1196_U146); 
assign P2_R2182_U41 = P2_R2182_U186 & P2_R2182_U182; 
assign P2_SUB_589_U6 = ~P2_U3614; 
assign P2_SUB_589_U7 = ~P2_U3615; 
assign P2_R2278_U188 = ~(P2_R2278_U128 & P2_R2278_U327); 
assign P2_R2278_U190 = ~(P2_R2278_U61 & P2_R2278_U260); 
assign P2_R2278_U518 = ~(P2_R2278_U258 & P2_R2278_U516); 
assign P2_R2278_U525 = ~(P2_R2278_U255 & P2_R2278_U523); 
assign P1_R2358_U134 = P1_R2358_U561 & P1_R2358_U305; 
assign P1_R2358_U180 = P1_R2358_U568 & P1_R2358_U567; 
assign P1_R2358_U181 = P1_R2358_U570 & P1_R2358_U569; 
assign P1_R2358_U565 = ~(P1_R2358_U135 & P1_R2358_U302 & P1_R2358_U179); 
assign P1_R2358_U566 = ~(P1_R2358_U561 & P1_R2358_U305 & P1_R2358_U301); 
assign P1_R2358_U573 = ~(P1_R2358_U572 & P1_R2358_U571); 
assign P3_U2831 = P3_U6396 & P3_U7906; 
assign P2_U2832 = ~(P2_U6764 & P2_U4149); 
assign P2_U3600 = ~(P2_U8102 & P2_U8101); 
assign P2_U3601 = ~(P2_U8104 & P2_U8103); 
assign P2_U3687 = ~(P2_U8430 & P2_U8429); 
assign P2_U6403 = ~(P2_ADD_391_1196_U104 & P2_U2397); 
assign P2_U6544 = ~(P2_U2379 & P2_R2099_U79); 
assign P2_U6561 = ~(P2_R2182_U41 & P2_U2393); 
assign P2_U6774 = ~(P2_U2392 & P2_R2099_U79); 
assign P2_U8432 = ~(P2_SUB_589_U6 & P2_STATE2_REG_1__SCAN_IN); 
assign P2_U8434 = ~(P2_SUB_589_U7 & P2_STATE2_REG_1__SCAN_IN); 
assign P1_U2811 = ~(P1_U6579 & P1_U3944 & P1_U3945 & P1_U6577 & P1_U6581); 
assign P1_U2843 = ~(P1_U6353 & P1_U6354 & P1_U6352); 
assign P1_U2875 = ~(P1_U6255 & P1_U6254 & P1_U6257 & P1_U6256); 
assign P1_U2970 = ~(P1_U5946 & P1_U5944 & P1_U5948 & P1_U5945 & P1_U5947); 
assign P2_R2099_U57 = ~(P2_U2722 & P2_R2099_U140); 
assign P2_R2099_U188 = ~(P2_R2099_U140 & P2_R2099_U56); 
assign P2_ADD_391_1196_U119 = ~P2_R2182_U41; 
assign P2_ADD_391_1196_U142 = ~(P2_ADD_391_1196_U242 & P2_ADD_391_1196_U241); 
assign P2_ADD_391_1196_U339 = ~(P2_R2182_U41 & P2_ADD_391_1196_U120); 
assign P2_ADD_391_1196_U341 = ~(P2_R2182_U41 & P2_ADD_391_1196_U120); 
assign P2_ADD_391_1196_U352 = ~(P2_R2096_U78 & P2_ADD_391_1196_U81); 
assign P2_ADD_391_1196_U354 = ~(P2_R2096_U78 & P2_ADD_391_1196_U81); 
assign P2_ADD_391_1196_U432 = ~(P2_ADD_391_1196_U239 & P2_ADD_391_1196_U430); 
assign P2_R2278_U106 = ~(P2_R2278_U518 & P2_R2278_U517); 
assign P2_R2278_U107 = ~(P2_R2278_U525 & P2_R2278_U524); 
assign P2_R2278_U262 = ~P2_R2278_U190; 
assign P2_R2278_U265 = ~P2_R2278_U188; 
assign P2_R2278_U267 = ~(P2_R2278_U266 & P2_R2278_U188); 
assign P2_R2278_U329 = ~(P2_R2278_U144 & P2_R2278_U188); 
assign P2_R2278_U333 = ~(P2_R2278_U266 & P2_R2278_U188 & P2_R2278_U129); 
assign P2_R2278_U503 = ~(P2_R2278_U187 & P2_R2278_U188); 
assign P2_R2278_U510 = ~(P2_R2278_U189 & P2_R2278_U190); 
assign P1_R2358_U374 = ~(P1_R2358_U300 & P1_R2358_U183 & P1_R2358_U134); 
assign P1_R2358_U574 = ~(P1_R2358_U181 & P1_R2358_U182); 
assign P1_R2358_U575 = ~(P1_R2358_U303 & P1_R2358_U573); 
assign P2_U2863 = ~(P2_U6544 & P2_U6545 & P2_U6543); 
assign P2_U2901 = ~(P2_U6402 & P2_U6401 & P2_U6405 & P2_U6404 & P2_U6403); 
assign P2_U3688 = ~(P2_U8432 & P2_U8431); 
assign P2_U3689 = ~(P2_U8434 & P2_U8433); 
assign P2_U4152 = P2_U6771 & P2_U6773 & P2_U6774 & P2_U6776 & P2_U4153; 
assign P2_R2099_U78 = ~(P2_R2099_U188 & P2_R2099_U187); 
assign P2_R2099_U141 = ~P2_R2099_U57; 
assign P2_R2099_U185 = ~(P2_U2721 & P2_R2099_U57); 
assign P2_ADD_391_1196_U103 = ~(P2_ADD_391_1196_U432 & P2_ADD_391_1196_U431); 
assign P2_ADD_391_1196_U124 = P2_ADD_391_1196_U352 & P2_ADD_391_1196_U351; 
assign P2_ADD_391_1196_U243 = ~P2_ADD_391_1196_U142; 
assign P2_ADD_391_1196_U245 = ~(P2_ADD_391_1196_U244 & P2_ADD_391_1196_U142); 
assign P2_ADD_391_1196_U340 = ~(P2_R2096_U76 & P2_ADD_391_1196_U119); 
assign P2_ADD_391_1196_U342 = ~(P2_R2096_U76 & P2_ADD_391_1196_U119); 
assign P2_ADD_391_1196_U355 = ~(P2_ADD_391_1196_U354 & P2_ADD_391_1196_U353); 
assign P2_ADD_391_1196_U419 = ~(P2_ADD_391_1196_U141 & P2_ADD_391_1196_U142); 
assign P2_R2243_U6 = ~(P2_U3686 | P2_U3685 | P2_U3684 | P2_U3687); 
assign P2_R2278_U182 = ~(P2_R2278_U131 & P2_R2278_U333); 
assign P2_R2278_U184 = ~(P2_R2278_U330 & P2_R2278_U329); 
assign P2_R2278_U186 = ~(P2_R2278_U268 & P2_R2278_U267); 
assign P2_R2278_U504 = ~(P2_R2278_U265 & P2_R2278_U502); 
assign P2_R2278_U511 = ~(P2_R2278_U262 & P2_R2278_U509); 
assign P1_R2358_U85 = ~(P1_R2358_U575 & P1_R2358_U574); 
assign P1_R2358_U136 = P1_R2358_U180 & P1_R2358_U374; 
assign P2_U2831 = ~(P2_U6772 & P2_U4152); 
assign P2_U6408 = ~(P2_ADD_391_1196_U103 & P2_U2397); 
assign P2_U6547 = ~(P2_U2379 & P2_R2099_U78); 
assign P2_U6782 = ~(P2_U2392 & P2_R2099_U78); 
assign P1_U5952 = ~(P1_R2358_U85 & P1_U2364); 
assign P1_U6260 = ~(P1_U2386 & P1_R2358_U85); 
assign P1_U6355 = ~(P1_U2383 & P1_R2358_U85); 
assign P1_U6588 = ~(P1_U2367 & P1_R2358_U85); 
assign P2_R2099_U59 = ~(P2_U2721 & P2_R2099_U141); 
assign P2_R2099_U186 = ~(P2_R2099_U141 & P2_R2099_U58); 
assign P2_ADD_391_1196_U121 = P2_ADD_391_1196_U340 & P2_ADD_391_1196_U339; 
assign P2_ADD_391_1196_U140 = ~(P2_ADD_391_1196_U246 & P2_ADD_391_1196_U245); 
assign P2_ADD_391_1196_U343 = ~(P2_ADD_391_1196_U342 & P2_ADD_391_1196_U341); 
assign P2_ADD_391_1196_U420 = ~(P2_ADD_391_1196_U243 & P2_ADD_391_1196_U418); 
assign P2_R2243_U9 = ~(P2_U3689 | P2_U3687 | P2_U3684 | P2_U3686 | P2_U3685); 
assign P2_R2243_U10 = ~P2_U3688; 
assign P2_R2278_U104 = ~(P2_R2278_U504 & P2_R2278_U503); 
assign P2_R2278_U105 = ~(P2_R2278_U511 & P2_R2278_U510); 
assign P2_R2278_U269 = ~P2_R2278_U186; 
assign P2_R2278_U272 = ~P2_R2278_U184; 
assign P2_R2278_U275 = ~P2_R2278_U182; 
assign P2_R2278_U277 = ~(P2_R2278_U276 & P2_R2278_U182); 
assign P2_R2278_U335 = ~(P2_R2278_U132 & P2_R2278_U182); 
assign P2_R2278_U477 = ~(P2_R2278_U181 & P2_R2278_U182); 
assign P2_R2278_U484 = ~(P2_R2278_U183 & P2_R2278_U184); 
assign P2_R2278_U496 = ~(P2_R2278_U185 & P2_R2278_U186); 
assign P1_R2358_U22 = P1_R2358_U566 & P1_R2358_U565 & P1_R2358_U136; 
assign P2_U2830 = ~(P2_U6779 & P2_U6781 & P2_U6782 & P2_U4156 & P2_U6780); 
assign P2_U2862 = ~(P2_U6547 & P2_U6548 & P2_U6546); 
assign P2_U2900 = ~(P2_U6407 & P2_U6406 & P2_U6410 & P2_U6409 & P2_U6408); 
assign P1_U2810 = ~(P1_U6586 & P1_U3946 & P1_U3947 & P1_U6584 & P1_U6588); 
assign P1_U2842 = ~(P1_U6356 & P1_U6357 & P1_U6355); 
assign P1_U2874 = ~(P1_U6259 & P1_U6258 & P1_U6261 & P1_U6260); 
assign P1_U2969 = ~(P1_U5951 & P1_U5949 & P1_U5953 & P1_U5950 & P1_U5952); 
assign P1_U3479 = P1_R2358_U22 & P1_U4449; 
assign P1_U5957 = ~(P1_R2358_U22 & P1_U2364); 
assign P1_U6595 = ~(P1_U2367 & P1_R2358_U22); 
assign P2_R2099_U77 = ~(P2_R2099_U186 & P2_R2099_U185); 
assign P2_R2099_U142 = ~P2_R2099_U59; 
assign P2_R2099_U183 = ~(P2_U2720 & P2_R2099_U59); 
assign P2_ADD_391_1196_U102 = ~(P2_ADD_391_1196_U420 & P2_ADD_391_1196_U419); 
assign P2_ADD_391_1196_U247 = ~P2_ADD_391_1196_U140; 
assign P2_ADD_391_1196_U249 = ~(P2_ADD_391_1196_U248 & P2_ADD_391_1196_U140); 
assign P2_ADD_391_1196_U412 = ~(P2_ADD_391_1196_U139 & P2_ADD_391_1196_U140); 
assign P2_R2243_U7 = ~(P2_U3684 | P2_R2243_U9); 
assign P2_R2243_U11 = ~(P2_R2243_U6 & P2_R2243_U10); 
assign P2_R2278_U178 = ~(P2_R2278_U133 & P2_R2278_U335); 
assign P2_R2278_U180 = ~(P2_R2278_U68 & P2_R2278_U277); 
assign P2_R2278_U478 = ~(P2_R2278_U275 & P2_R2278_U476); 
assign P2_R2278_U485 = ~(P2_R2278_U272 & P2_R2278_U483); 
assign P2_R2278_U497 = ~(P2_R2278_U269 & P2_R2278_U495); 
assign P2_U6413 = ~(P2_ADD_391_1196_U102 & P2_U2397); 
assign P2_U6550 = ~(P2_U2379 & P2_R2099_U77); 
assign P2_U6790 = ~(P2_U2392 & P2_R2099_U77); 
assign P1_U2809 = ~(P1_U6593 & P1_U3948 & P1_U3949 & P1_U6591 & P1_U6595); 
assign P1_U2968 = ~(P1_U5956 & P1_U5954 & P1_U5958 & P1_U5955 & P1_U5957); 
assign P1_U7745 = ~(P1_U3479 & P1_U4223); 
assign P2_R2099_U61 = ~(P2_U2720 & P2_R2099_U142); 
assign P2_R2099_U184 = ~(P2_R2099_U142 & P2_R2099_U60); 
assign P2_ADD_391_1196_U138 = ~(P2_ADD_391_1196_U250 & P2_ADD_391_1196_U249); 
assign P2_ADD_391_1196_U413 = ~(P2_ADD_391_1196_U247 & P2_ADD_391_1196_U411); 
assign P2_R2243_U8 = ~(P2_R2243_U7 & P2_R2243_U11); 
assign P2_R2278_U101 = ~(P2_R2278_U478 & P2_R2278_U477); 
assign P2_R2278_U102 = ~(P2_R2278_U485 & P2_R2278_U484); 
assign P2_R2278_U103 = ~(P2_R2278_U497 & P2_R2278_U496); 
assign P2_R2278_U279 = ~P2_R2278_U180; 
assign P2_R2278_U282 = ~P2_R2278_U178; 
assign P2_R2278_U284 = ~(P2_R2278_U283 & P2_R2278_U178); 
assign P2_R2278_U337 = ~(P2_R2278_U134 & P2_R2278_U178); 
assign P2_R2278_U463 = ~(P2_R2278_U177 & P2_R2278_U178); 
assign P2_R2278_U470 = ~(P2_R2278_U179 & P2_R2278_U180); 
assign P2_U2829 = ~(P2_U6787 & P2_U6789 & P2_U4158 & P2_U6790 & P2_U6788); 
assign P2_U2861 = ~(P2_U6550 & P2_U6551 & P2_U6549); 
assign P2_U2899 = ~(P2_U6412 & P2_U6411 & P2_U6415 & P2_U6414 & P2_U6413); 
assign P2_U3292 = ~P2_R2243_U8; 
assign P2_U4605 = ~(P2_R2243_U8 & P2_U4428); 
assign P2_U5642 = ~(P2_U2448 & P2_R2243_U8 & P2_STATE2_REG_0__SCAN_IN); 
assign P2_U8132 = ~(P2_R2243_U8 & P2_U2616); 
assign P1_U4176 = P1_U7745 & P1_U7744; 
assign P2_R2099_U76 = ~(P2_R2099_U184 & P2_R2099_U183); 
assign P2_R2099_U143 = ~P2_R2099_U61; 
assign P2_R2099_U181 = ~(P2_U2719 & P2_R2099_U61); 
assign P2_ADD_391_1196_U101 = ~(P2_ADD_391_1196_U413 & P2_ADD_391_1196_U412); 
assign P2_ADD_391_1196_U251 = ~P2_ADD_391_1196_U138; 
assign P2_ADD_391_1196_U253 = ~(P2_ADD_391_1196_U252 & P2_ADD_391_1196_U138); 
assign P2_ADD_391_1196_U405 = ~(P2_ADD_391_1196_U137 & P2_ADD_391_1196_U138); 
assign P2_R2278_U174 = ~(P2_R2278_U135 & P2_R2278_U337); 
assign P2_R2278_U176 = ~(P2_R2278_U71 & P2_R2278_U284); 
assign P2_R2278_U464 = ~(P2_R2278_U282 & P2_R2278_U462); 
assign P2_R2278_U471 = ~(P2_R2278_U279 & P2_R2278_U469); 
assign P2_U3533 = ~(P2_U4455 & P2_U3306 & P2_U5642); 
assign P2_U4399 = P2_U8132 & P2_U8131; 
assign P2_U4464 = ~(P2_U2448 & P2_U3292); 
assign P2_U4607 = ~(P2_U4606 & P2_U4605); 
assign P2_U4611 = ~(P2_U4428 & P2_U3292); 
assign P2_U5665 = ~(P2_U2616 & P2_U3292); 
assign P2_U6418 = ~(P2_ADD_391_1196_U101 & P2_U2397); 
assign P2_U6553 = ~(P2_U2379 & P2_R2099_U76); 
assign P2_U6798 = ~(P2_U2392 & P2_R2099_U76); 
assign P1_U2873 = ~(P1_U4176 & P1_U6262); 
assign P2_R2099_U63 = ~(P2_U2719 & P2_R2099_U143); 
assign P2_R2099_U182 = ~(P2_R2099_U143 & P2_R2099_U62); 
assign P2_ADD_391_1196_U136 = ~(P2_ADD_391_1196_U254 & P2_ADD_391_1196_U253); 
assign P2_ADD_391_1196_U406 = ~(P2_ADD_391_1196_U251 & P2_ADD_391_1196_U404); 
assign P2_R2278_U99 = ~(P2_R2278_U464 & P2_R2278_U463); 
assign P2_R2278_U100 = ~(P2_R2278_U471 & P2_R2278_U470); 
assign P2_R2278_U205 = ~(P2_U2796 & P2_R2278_U174); 
assign P2_R2278_U286 = ~P2_R2278_U176; 
assign P2_R2278_U289 = ~P2_R2278_U174; 
assign P2_R2278_U290 = ~(P2_R2278_U174 & P2_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P2_R2278_U444 = ~(P2_R2278_U174 & P2_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P2_R2278_U446 = ~(P2_R2278_U174 & P2_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P2_R2278_U456 = ~(P2_R2278_U175 & P2_R2278_U176); 
assign P2_U2828 = ~(P2_U6795 & P2_U6797 & P2_U4160 & P2_U6798 & P2_U6796); 
assign P2_U2860 = ~(P2_U6553 & P2_U6554 & P2_U6552); 
assign P2_U2898 = ~(P2_U6417 & P2_U6416 & P2_U6420 & P2_U6419 & P2_U6418); 
assign P2_U4608 = ~(P2_U4420 & P2_U4607); 
assign P2_U4613 = ~(P2_U4612 & P2_U4611); 
assign P2_U5643 = ~P2_U3533; 
assign P2_U5664 = ~(P2_U5662 & P2_U5663 & P2_U4464); 
assign P2_U5667 = ~(P2_U5666 & P2_U5665); 
assign P2_U6839 = ~(P2_U4426 & P2_U4468 & P2_U4399); 
assign P2_U8106 = ~(P2_U5651 & P2_U3533); 
assign P2_U8111 = ~(P2_U5655 & P2_U3533); 
assign P2_U8113 = ~(P2_U5660 & P2_U3533); 
assign P2_R2099_U75 = ~(P2_R2099_U182 & P2_R2099_U181); 
assign P2_R2099_U144 = ~P2_R2099_U63; 
assign P2_R2099_U179 = ~(P2_U2718 & P2_R2099_U63); 
assign P2_ADD_391_1196_U100 = ~(P2_ADD_391_1196_U406 & P2_ADD_391_1196_U405); 
assign P2_ADD_391_1196_U255 = ~P2_ADD_391_1196_U136; 
assign P2_ADD_391_1196_U257 = ~(P2_ADD_391_1196_U256 & P2_ADD_391_1196_U136); 
assign P2_ADD_391_1196_U398 = ~(P2_ADD_391_1196_U135 & P2_ADD_391_1196_U136); 
assign P2_R2278_U173 = ~(P2_R2278_U290 & P2_R2278_U205 & P2_R2278_U308); 
assign P2_R2278_U445 = ~(P2_R2278_U289 & P2_R2278_U73); 
assign P2_R2278_U447 = ~(P2_R2278_U289 & P2_R2278_U73); 
assign P2_R2278_U457 = ~(P2_R2278_U286 & P2_R2278_U455); 
assign P2_U2819 = ~(P2_U6840 & P2_U6839); 
assign P2_U3047 = P2_U5643 & P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign P2_U3257 = ~(P2_U8051 & P2_U8050 & P2_U4609 & P2_U4608); 
assign P2_U4614 = ~(P2_U4420 & P2_U4613); 
assign P2_U5669 = ~(P2_U4420 & P2_U5667); 
assign P2_U5936 = ~(P2_U4420 & P2_U2374 & P2_U4613); 
assign P2_U6423 = ~(P2_ADD_391_1196_U100 & P2_U2397); 
assign P2_U6556 = ~(P2_U2379 & P2_R2099_U75); 
assign P2_U6806 = ~(P2_U2392 & P2_R2099_U75); 
assign P2_U8105 = ~(P2_U5643 & P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign P2_U8110 = ~(P2_U5643 & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign P2_U8112 = ~(P2_U5643 & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign P2_U8114 = ~(P2_U5643 & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign P2_U8115 = ~(P2_U5664 & P2_U3533); 
assign P2_R2099_U65 = ~(P2_U2718 & P2_R2099_U144); 
assign P2_R2099_U180 = ~(P2_R2099_U144 & P2_R2099_U64); 
assign P2_ADD_391_1196_U134 = ~(P2_ADD_391_1196_U258 & P2_ADD_391_1196_U257); 
assign P2_ADD_391_1196_U399 = ~(P2_ADD_391_1196_U255 & P2_ADD_391_1196_U397); 
assign P2_R2278_U98 = ~(P2_R2278_U457 & P2_R2278_U456); 
assign P2_R2278_U291 = ~P2_R2278_U173; 
assign P2_R2278_U293 = ~(P2_R2278_U292 & P2_R2278_U173); 
assign P2_R2278_U339 = ~(P2_R2278_U143 & P2_R2278_U173); 
assign P2_R2278_U342 = ~(P2_R2278_U173 & P2_R2278_U136); 
assign P2_R2278_U442 = ~(P2_R2278_U172 & P2_R2278_U173); 
assign P2_R2278_U448 = ~(P2_R2278_U447 & P2_R2278_U446); 
assign P2_R2278_U449 = ~(P2_R2278_U445 & P2_R2278_U444 & P2_R2278_U72); 
assign P2_U2827 = ~(P2_U6803 & P2_U6805 & P2_U4162 & P2_U6806 & P2_U6804); 
assign P2_U2859 = ~(P2_U6556 & P2_U6557 & P2_U6555); 
assign P2_U2897 = ~(P2_U6422 & P2_U6421 & P2_U6425 & P2_U6424 & P2_U6423); 
assign P2_U3537 = ~(P2_U5937 & P2_U5936); 
assign P2_U3602 = ~(P2_U8106 & P2_U8105); 
assign P2_U3603 = ~(P2_U8111 & P2_U8110); 
assign P2_U3604 = ~(P2_U8113 & P2_U8112); 
assign P2_U3605 = ~(P2_U8115 & P2_U8114); 
assign P2_U4610 = ~P2_U3257; 
assign P2_U5670 = ~(P2_U2512 & P2_U3894 & P2_U4397 & P2_U5669); 
assign P2_U8133 = ~(P2_U6838 & P2_U3257); 
assign P2_R2099_U74 = ~(P2_R2099_U180 & P2_R2099_U179); 
assign P2_R2099_U145 = ~P2_R2099_U65; 
assign P2_R2099_U170 = ~(P2_U2717 & P2_R2099_U65); 
assign P2_ADD_391_1196_U99 = ~(P2_ADD_391_1196_U399 & P2_ADD_391_1196_U398); 
assign P2_ADD_391_1196_U259 = ~P2_ADD_391_1196_U134; 
assign P2_ADD_391_1196_U261 = ~(P2_ADD_391_1196_U260 & P2_ADD_391_1196_U134); 
assign P2_ADD_391_1196_U391 = ~(P2_ADD_391_1196_U133 & P2_ADD_391_1196_U134); 
assign P2_R2278_U167 = ~(P2_R2278_U140 & P2_R2278_U342); 
assign P2_R2278_U169 = ~(P2_R2278_U341 & P2_R2278_U339); 
assign P2_R2278_U171 = ~(P2_R2278_U78 & P2_R2278_U293); 
assign P2_R2278_U344 = ~(P2_R2278_U343 & P2_R2278_U342 & P2_R2278_U137); 
assign P2_R2278_U443 = ~(P2_R2278_U291 & P2_R2278_U441); 
assign P2_R2278_U450 = ~(P2_R2278_U448 & P2_U2796); 
assign P2_U2370 = P2_U2447 & P2_U3537; 
assign P2_U2371 = P2_U3990 & P2_U3537; 
assign P2_U2372 = P2_U3989 & P2_U3537; 
assign P2_U2373 = P2_U4419 & P2_U3537; 
assign P2_U2387 = P2_U5940 & P2_U3537; 
assign P2_U3298 = ~(P2_U7894 & P2_U4444 & P2_LT_563_U6 & P2_U4614 & P2_U4610); 
assign P2_U3609 = ~(P2_U8134 & P2_U8133); 
assign P2_U5671 = ~(P2_U2374 & P2_U5670); 
assign P2_U5938 = ~P2_U3537; 
assign P2_U6428 = ~(P2_ADD_391_1196_U99 & P2_U2397); 
assign P2_U6559 = ~(P2_U2379 & P2_R2099_U74); 
assign P2_U6814 = ~(P2_U2392 & P2_R2099_U74); 
assign P2_R2099_U102 = ~(P2_U2717 & P2_R2099_U145); 
assign P2_R2099_U171 = ~(P2_R2099_U145 & P2_R2099_U66); 
assign P2_ADD_391_1196_U132 = ~(P2_ADD_391_1196_U262 & P2_ADD_391_1196_U261); 
assign P2_ADD_391_1196_U392 = ~(P2_ADD_391_1196_U259 & P2_ADD_391_1196_U390); 
assign P2_R2278_U96 = ~(P2_R2278_U443 & P2_R2278_U442); 
assign P2_R2278_U97 = ~(P2_R2278_U450 & P2_R2278_U449); 
assign P2_R2278_U206 = ~(P2_R2278_U139 & P2_R2278_U344); 
assign P2_R2278_U295 = ~P2_R2278_U171; 
assign P2_R2278_U298 = ~P2_R2278_U169; 
assign P2_R2278_U301 = ~P2_R2278_U167; 
assign P2_R2278_U303 = ~(P2_R2278_U302 & P2_R2278_U167); 
assign P2_R2278_U421 = ~(P2_R2278_U166 & P2_R2278_U167); 
assign P2_R2278_U428 = ~(P2_R2278_U168 & P2_R2278_U169); 
assign P2_R2278_U435 = ~(P2_R2278_U170 & P2_R2278_U171); 
assign P2_U2826 = ~(P2_U6811 & P2_U6813 & P2_U4164 & P2_U6814 & P2_U6812); 
assign P2_U2858 = ~(P2_U6559 & P2_U6560 & P2_U6558); 
assign P2_U2896 = ~(P2_U6427 & P2_U6426 & P2_U6430 & P2_U6429 & P2_U6428); 
assign P2_U3535 = ~(P2_U5672 & P2_U5671); 
assign P2_U4616 = ~P2_U3298; 
assign P2_U4632 = ~(P2_U2374 & P2_U3298); 
assign P2_U5941 = ~(P2_U2387 & P2_PHYADDRPOINTER_REG_0__SCAN_IN); 
assign P2_U5942 = ~(P2_U2373 & P2_ADD_371_1212_U68); 
assign P2_U5943 = ~(P2_U2372 & P2_R2099_U94); 
assign P2_U5944 = ~(P2_U2371 & P2_REIP_REG_0__SCAN_IN); 
assign P2_U5945 = ~(P2_U2370 & P2_R2278_U83); 
assign P2_U5946 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_0__SCAN_IN); 
assign P2_U5947 = ~(P2_R2337_U4 & P2_U2387); 
assign P2_U5948 = ~(P2_U2373 & P2_ADD_371_1212_U25); 
assign P2_U5949 = ~(P2_U2372 & P2_R2099_U5); 
assign P2_U5950 = ~(P2_U2371 & P2_REIP_REG_1__SCAN_IN); 
assign P2_U5951 = ~(P2_U2370 & P2_R2278_U6); 
assign P2_U5952 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_1__SCAN_IN); 
assign P2_U5953 = ~(P2_R2337_U70 & P2_U2387); 
assign P2_U5954 = ~(P2_U2373 & P2_ADD_371_1212_U79); 
assign P2_U5955 = ~(P2_U2372 & P2_R2099_U96); 
assign P2_U5956 = ~(P2_U2371 & P2_REIP_REG_2__SCAN_IN); 
assign P2_U5957 = ~(P2_U2370 & P2_R2278_U92); 
assign P2_U5958 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_2__SCAN_IN); 
assign P2_U5959 = ~(P2_R2337_U67 & P2_U2387); 
assign P2_U5960 = ~(P2_U2373 & P2_ADD_371_1212_U84); 
assign P2_U5961 = ~(P2_U2372 & P2_R2099_U95); 
assign P2_U5962 = ~(P2_U2371 & P2_REIP_REG_3__SCAN_IN); 
assign P2_U5963 = ~(P2_U2370 & P2_R2278_U90); 
assign P2_U5964 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_3__SCAN_IN); 
assign P2_U5965 = ~(P2_R2337_U66 & P2_U2387); 
assign P2_U5966 = ~(P2_U2373 & P2_ADD_371_1212_U80); 
assign P2_U5967 = ~(P2_U2372 & P2_R2099_U98); 
assign P2_U5968 = ~(P2_U2371 & P2_REIP_REG_4__SCAN_IN); 
assign P2_U5969 = ~(P2_U2370 & P2_R2278_U89); 
assign P2_U5970 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_4__SCAN_IN); 
assign P2_U5971 = ~(P2_R2337_U65 & P2_U2387); 
assign P2_U5972 = ~(P2_U2373 & P2_ADD_371_1212_U81); 
assign P2_U5973 = ~(P2_U2372 & P2_R2099_U71); 
assign P2_U5974 = ~(P2_U2371 & P2_REIP_REG_5__SCAN_IN); 
assign P2_U5975 = ~(P2_U2370 & P2_R2278_U88); 
assign P2_U5976 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_5__SCAN_IN); 
assign P2_U5977 = ~(P2_R2337_U64 & P2_U2387); 
assign P2_U5978 = ~(P2_U2373 & P2_ADD_371_1212_U78); 
assign P2_U5979 = ~(P2_U2372 & P2_R2099_U70); 
assign P2_U5980 = ~(P2_U2371 & P2_REIP_REG_6__SCAN_IN); 
assign P2_U5981 = ~(P2_U2370 & P2_R2278_U87); 
assign P2_U5982 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_6__SCAN_IN); 
assign P2_U5983 = ~(P2_R2337_U63 & P2_U2387); 
assign P2_U5984 = ~(P2_U2373 & P2_ADD_371_1212_U85); 
assign P2_U5985 = ~(P2_U2372 & P2_R2099_U69); 
assign P2_U5986 = ~(P2_U2371 & P2_REIP_REG_7__SCAN_IN); 
assign P2_U5987 = ~(P2_U2370 & P2_R2278_U86); 
assign P2_U5988 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_7__SCAN_IN); 
assign P2_U5989 = ~(P2_R2337_U62 & P2_U2387); 
assign P2_U5990 = ~(P2_U2373 & P2_ADD_371_1212_U82); 
assign P2_U5991 = ~(P2_U2372 & P2_R2099_U68); 
assign P2_U5992 = ~(P2_U2371 & P2_REIP_REG_8__SCAN_IN); 
assign P2_U5993 = ~(P2_U2370 & P2_R2278_U85); 
assign P2_U5994 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_8__SCAN_IN); 
assign P2_U5995 = ~(P2_R2337_U61 & P2_U2387); 
assign P2_U5996 = ~(P2_U2373 & P2_ADD_371_1212_U118); 
assign P2_U5997 = ~(P2_U2372 & P2_R2099_U67); 
assign P2_U5998 = ~(P2_U2371 & P2_REIP_REG_9__SCAN_IN); 
assign P2_U5999 = ~(P2_U2370 & P2_R2278_U84); 
assign P2_U6000 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_9__SCAN_IN); 
assign P2_U6001 = ~(P2_R2337_U90 & P2_U2387); 
assign P2_U6002 = ~(P2_U2373 & P2_ADD_371_1212_U13); 
assign P2_U6003 = ~(P2_U2372 & P2_R2099_U93); 
assign P2_U6004 = ~(P2_U2371 & P2_REIP_REG_10__SCAN_IN); 
assign P2_U6005 = ~(P2_U2370 & P2_R2278_U112); 
assign P2_U6006 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_10__SCAN_IN); 
assign P2_U6007 = ~(P2_R2337_U89 & P2_U2387); 
assign P2_U6008 = ~(P2_U2373 & P2_ADD_371_1212_U14); 
assign P2_U6009 = ~(P2_U2372 & P2_R2099_U92); 
assign P2_U6010 = ~(P2_U2371 & P2_REIP_REG_11__SCAN_IN); 
assign P2_U6011 = ~(P2_U2370 & P2_R2278_U111); 
assign P2_U6012 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_11__SCAN_IN); 
assign P2_U6013 = ~(P2_R2337_U88 & P2_U2387); 
assign P2_U6014 = ~(P2_U2373 & P2_ADD_371_1212_U76); 
assign P2_U6015 = ~(P2_U2372 & P2_R2099_U91); 
assign P2_U6016 = ~(P2_U2371 & P2_REIP_REG_12__SCAN_IN); 
assign P2_U6017 = ~(P2_U2370 & P2_R2278_U110); 
assign P2_U6018 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_12__SCAN_IN); 
assign P2_U6019 = ~(P2_R2337_U87 & P2_U2387); 
assign P2_U6020 = ~(P2_U2373 & P2_ADD_371_1212_U15); 
assign P2_U6021 = ~(P2_U2372 & P2_R2099_U90); 
assign P2_U6022 = ~(P2_U2371 & P2_REIP_REG_13__SCAN_IN); 
assign P2_U6023 = ~(P2_U2370 & P2_R2278_U109); 
assign P2_U6024 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_13__SCAN_IN); 
assign P2_U6025 = ~(P2_R2337_U86 & P2_U2387); 
assign P2_U6026 = ~(P2_U2373 & P2_ADD_371_1212_U16); 
assign P2_U6027 = ~(P2_U2372 & P2_R2099_U89); 
assign P2_U6028 = ~(P2_U2371 & P2_REIP_REG_14__SCAN_IN); 
assign P2_U6029 = ~(P2_U2370 & P2_R2278_U108); 
assign P2_U6030 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_14__SCAN_IN); 
assign P2_U6031 = ~(P2_R2337_U85 & P2_U2387); 
assign P2_U6032 = ~(P2_U2373 & P2_ADD_371_1212_U73); 
assign P2_U6033 = ~(P2_U2372 & P2_R2099_U88); 
assign P2_U6034 = ~(P2_U2371 & P2_REIP_REG_15__SCAN_IN); 
assign P2_U6035 = ~(P2_U2370 & P2_R2278_U107); 
assign P2_U6036 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_15__SCAN_IN); 
assign P2_U6037 = ~(P2_R2337_U84 & P2_U2387); 
assign P2_U6038 = ~(P2_U2373 & P2_ADD_371_1212_U17); 
assign P2_U6039 = ~(P2_U2372 & P2_R2099_U87); 
assign P2_U6040 = ~(P2_U2371 & P2_REIP_REG_16__SCAN_IN); 
assign P2_U6041 = ~(P2_U2370 & P2_R2278_U106); 
assign P2_U6042 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_16__SCAN_IN); 
assign P2_U6043 = ~(P2_R2337_U83 & P2_U2387); 
assign P2_U6044 = ~(P2_U2373 & P2_ADD_371_1212_U71); 
assign P2_U6045 = ~(P2_U2372 & P2_R2099_U86); 
assign P2_U6046 = ~(P2_U2371 & P2_REIP_REG_17__SCAN_IN); 
assign P2_U6047 = ~(P2_U2370 & P2_R2278_U105); 
assign P2_U6048 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_17__SCAN_IN); 
assign P2_U6049 = ~(P2_R2337_U82 & P2_U2387); 
assign P2_U6050 = ~(P2_U2373 & P2_ADD_371_1212_U72); 
assign P2_U6051 = ~(P2_U2372 & P2_R2099_U85); 
assign P2_U6052 = ~(P2_U2371 & P2_REIP_REG_18__SCAN_IN); 
assign P2_U6053 = ~(P2_U2370 & P2_R2278_U104); 
assign P2_U6054 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_18__SCAN_IN); 
assign P2_U6055 = ~(P2_R2337_U81 & P2_U2387); 
assign P2_U6056 = ~(P2_U2373 & P2_ADD_371_1212_U18); 
assign P2_U6057 = ~(P2_U2372 & P2_R2099_U84); 
assign P2_U6058 = ~(P2_U2371 & P2_REIP_REG_19__SCAN_IN); 
assign P2_U6059 = ~(P2_U2370 & P2_R2278_U103); 
assign P2_U6060 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_19__SCAN_IN); 
assign P2_U6061 = ~(P2_R2337_U80 & P2_U2387); 
assign P2_U6062 = ~(P2_U2373 & P2_ADD_371_1212_U19); 
assign P2_U6063 = ~(P2_U2372 & P2_R2099_U83); 
assign P2_U6064 = ~(P2_U2371 & P2_REIP_REG_20__SCAN_IN); 
assign P2_U6065 = ~(P2_U2370 & P2_R2278_U102); 
assign P2_U6066 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_20__SCAN_IN); 
assign P2_U6067 = ~(P2_R2337_U79 & P2_U2387); 
assign P2_U6068 = ~(P2_U2373 & P2_ADD_371_1212_U75); 
assign P2_U6069 = ~(P2_U2372 & P2_R2099_U82); 
assign P2_U6070 = ~(P2_U2371 & P2_REIP_REG_21__SCAN_IN); 
assign P2_U6071 = ~(P2_U2370 & P2_R2278_U101); 
assign P2_U6072 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_21__SCAN_IN); 
assign P2_U6073 = ~(P2_R2337_U78 & P2_U2387); 
assign P2_U6074 = ~(P2_U2373 & P2_ADD_371_1212_U20); 
assign P2_U6075 = ~(P2_U2372 & P2_R2099_U81); 
assign P2_U6076 = ~(P2_U2371 & P2_REIP_REG_22__SCAN_IN); 
assign P2_U6077 = ~(P2_U2370 & P2_R2278_U100); 
assign P2_U6078 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_22__SCAN_IN); 
assign P2_U6079 = ~(P2_R2337_U77 & P2_U2387); 
assign P2_U6080 = ~(P2_U2373 & P2_ADD_371_1212_U21); 
assign P2_U6081 = ~(P2_U2372 & P2_R2099_U80); 
assign P2_U6082 = ~(P2_U2371 & P2_REIP_REG_23__SCAN_IN); 
assign P2_U6083 = ~(P2_U2370 & P2_R2278_U99); 
assign P2_U6084 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_23__SCAN_IN); 
assign P2_U6085 = ~(P2_R2337_U76 & P2_U2387); 
assign P2_U6086 = ~(P2_U2373 & P2_ADD_371_1212_U70); 
assign P2_U6087 = ~(P2_U2372 & P2_R2099_U79); 
assign P2_U6088 = ~(P2_U2371 & P2_REIP_REG_24__SCAN_IN); 
assign P2_U6089 = ~(P2_U2370 & P2_R2278_U98); 
assign P2_U6090 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_24__SCAN_IN); 
assign P2_U6091 = ~(P2_R2337_U75 & P2_U2387); 
assign P2_U6092 = ~(P2_U2373 & P2_ADD_371_1212_U77); 
assign P2_U6093 = ~(P2_U2372 & P2_R2099_U78); 
assign P2_U6094 = ~(P2_U2371 & P2_REIP_REG_25__SCAN_IN); 
assign P2_U6095 = ~(P2_U2370 & P2_R2278_U97); 
assign P2_U6096 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_25__SCAN_IN); 
assign P2_U6097 = ~(P2_R2337_U74 & P2_U2387); 
assign P2_U6098 = ~(P2_U2373 & P2_ADD_371_1212_U22); 
assign P2_U6099 = ~(P2_U2372 & P2_R2099_U77); 
assign P2_U6100 = ~(P2_U2371 & P2_REIP_REG_26__SCAN_IN); 
assign P2_U6101 = ~(P2_U2370 & P2_R2278_U96); 
assign P2_U6102 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_26__SCAN_IN); 
assign P2_U6103 = ~(P2_R2337_U73 & P2_U2387); 
assign P2_U6104 = ~(P2_U2373 & P2_ADD_371_1212_U74); 
assign P2_U6105 = ~(P2_U2372 & P2_R2099_U76); 
assign P2_U6106 = ~(P2_U2371 & P2_REIP_REG_27__SCAN_IN); 
assign P2_U6108 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_27__SCAN_IN); 
assign P2_U6109 = ~(P2_R2337_U72 & P2_U2387); 
assign P2_U6110 = ~(P2_U2373 & P2_ADD_371_1212_U23); 
assign P2_U6111 = ~(P2_U2372 & P2_R2099_U75); 
assign P2_U6112 = ~(P2_U2371 & P2_REIP_REG_28__SCAN_IN); 
assign P2_U6114 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_28__SCAN_IN); 
assign P2_U6115 = ~(P2_R2337_U71 & P2_U2387); 
assign P2_U6116 = ~(P2_U2373 & P2_ADD_371_1212_U24); 
assign P2_U6117 = ~(P2_U2372 & P2_R2099_U74); 
assign P2_U6118 = ~(P2_U2371 & P2_REIP_REG_29__SCAN_IN); 
assign P2_U6120 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_29__SCAN_IN); 
assign P2_U6121 = ~(P2_R2337_U69 & P2_U2387); 
assign P2_U6122 = ~(P2_U2373 & P2_ADD_371_1212_U69); 
assign P2_U6124 = ~(P2_U2371 & P2_REIP_REG_30__SCAN_IN); 
assign P2_U6126 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_30__SCAN_IN); 
assign P2_U6127 = ~(P2_R2337_U68 & P2_U2387); 
assign P2_U6128 = ~(P2_U2373 & P2_ADD_371_1212_U83); 
assign P2_U6130 = ~(P2_U2371 & P2_REIP_REG_31__SCAN_IN); 
assign P2_U6132 = ~(P2_U5938 & P2_PHYADDRPOINTER_REG_31__SCAN_IN); 
assign P2_R2099_U73 = ~(P2_R2099_U171 & P2_R2099_U170); 
assign P2_R2099_U146 = ~P2_R2099_U102; 
assign P2_R2099_U168 = ~(P2_U2716 & P2_R2099_U102); 
assign P2_ADD_391_1196_U98 = ~(P2_ADD_391_1196_U392 & P2_ADD_391_1196_U391); 
assign P2_ADD_391_1196_U263 = ~P2_ADD_391_1196_U132; 
assign P2_ADD_391_1196_U265 = ~(P2_ADD_391_1196_U264 & P2_ADD_391_1196_U132); 
assign P2_ADD_391_1196_U384 = ~(P2_ADD_391_1196_U131 & P2_ADD_391_1196_U132); 
assign P2_R2278_U163 = ~(P2_R2278_U304 & P2_R2278_U303); 
assign P2_R2278_U309 = ~(P2_R2278_U303 & P2_R2278_U141); 
assign P2_R2278_U422 = ~(P2_R2278_U301 & P2_R2278_U420); 
assign P2_R2278_U429 = ~(P2_R2278_U298 & P2_R2278_U427); 
assign P2_R2278_U436 = ~(P2_R2278_U295 & P2_R2278_U434); 
assign P2_U2363 = P2_U3535 & P2_STATE2_REG_2__SCAN_IN; 
assign P2_U2381 = P2_U3535 & P2_U3270; 
assign P2_U3721 = P2_U3720 & P2_U4632; 
assign P2_U3991 = P2_U5942 & P2_U5941 & P2_U5943; 
assign P2_U3992 = P2_U5945 & P2_U5944 & P2_U5946; 
assign P2_U3993 = P2_U5948 & P2_U5947 & P2_U5949; 
assign P2_U3994 = P2_U5951 & P2_U5950 & P2_U5952; 
assign P2_U3995 = P2_U5954 & P2_U5953 & P2_U5955; 
assign P2_U3996 = P2_U5957 & P2_U5956 & P2_U5958; 
assign P2_U3997 = P2_U5960 & P2_U5959 & P2_U5961; 
assign P2_U3998 = P2_U5963 & P2_U5962 & P2_U5964; 
assign P2_U3999 = P2_U5966 & P2_U5965 & P2_U5967; 
assign P2_U4000 = P2_U5969 & P2_U5968 & P2_U5970; 
assign P2_U4001 = P2_U5972 & P2_U5971 & P2_U5973; 
assign P2_U4002 = P2_U5975 & P2_U5974 & P2_U5976; 
assign P2_U4003 = P2_U5978 & P2_U5977 & P2_U5979; 
assign P2_U4004 = P2_U5981 & P2_U5980 & P2_U5982; 
assign P2_U4005 = P2_U5984 & P2_U5983 & P2_U5985; 
assign P2_U4006 = P2_U5987 & P2_U5986 & P2_U5988; 
assign P2_U4007 = P2_U5990 & P2_U5989 & P2_U5991; 
assign P2_U4008 = P2_U5993 & P2_U5992 & P2_U5994; 
assign P2_U4009 = P2_U5996 & P2_U5995 & P2_U5997; 
assign P2_U4010 = P2_U5999 & P2_U5998 & P2_U6000; 
assign P2_U4011 = P2_U6002 & P2_U6001 & P2_U6003; 
assign P2_U4012 = P2_U6005 & P2_U6004 & P2_U6006; 
assign P2_U4013 = P2_U6008 & P2_U6007 & P2_U6009; 
assign P2_U4014 = P2_U6011 & P2_U6010 & P2_U6012; 
assign P2_U4015 = P2_U6014 & P2_U6013 & P2_U6015; 
assign P2_U4016 = P2_U6017 & P2_U6016 & P2_U6018; 
assign P2_U4017 = P2_U6020 & P2_U6019 & P2_U6021; 
assign P2_U4018 = P2_U6023 & P2_U6022 & P2_U6024; 
assign P2_U4019 = P2_U6026 & P2_U6025 & P2_U6027; 
assign P2_U4020 = P2_U6029 & P2_U6028 & P2_U6030; 
assign P2_U4021 = P2_U6032 & P2_U6031 & P2_U6033; 
assign P2_U4022 = P2_U6035 & P2_U6034 & P2_U6036; 
assign P2_U4023 = P2_U6038 & P2_U6037 & P2_U6039; 
assign P2_U4024 = P2_U6041 & P2_U6040 & P2_U6042; 
assign P2_U4025 = P2_U6044 & P2_U6043 & P2_U6045; 
assign P2_U4026 = P2_U6047 & P2_U6046 & P2_U6048; 
assign P2_U4027 = P2_U6050 & P2_U6049 & P2_U6051; 
assign P2_U4028 = P2_U6053 & P2_U6052 & P2_U6054; 
assign P2_U4029 = P2_U6056 & P2_U6055 & P2_U6057; 
assign P2_U4030 = P2_U6059 & P2_U6058 & P2_U6060; 
assign P2_U4031 = P2_U6062 & P2_U6061 & P2_U6063; 
assign P2_U4032 = P2_U6065 & P2_U6064 & P2_U6066; 
assign P2_U4033 = P2_U6068 & P2_U6067 & P2_U6069; 
assign P2_U4034 = P2_U6071 & P2_U6070 & P2_U6072; 
assign P2_U4035 = P2_U6074 & P2_U6073 & P2_U6075; 
assign P2_U4036 = P2_U6077 & P2_U6076 & P2_U6078; 
assign P2_U4037 = P2_U6080 & P2_U6079 & P2_U6081; 
assign P2_U4038 = P2_U6083 & P2_U6082 & P2_U6084; 
assign P2_U4039 = P2_U6086 & P2_U6085 & P2_U6087; 
assign P2_U4040 = P2_U6089 & P2_U6088 & P2_U6090; 
assign P2_U4041 = P2_U6092 & P2_U6091 & P2_U6093; 
assign P2_U4042 = P2_U6095 & P2_U6094 & P2_U6096; 
assign P2_U4043 = P2_U6098 & P2_U6097 & P2_U6099; 
assign P2_U4044 = P2_U6101 & P2_U6100 & P2_U6102; 
assign P2_U4045 = P2_U6104 & P2_U6103 & P2_U6105; 
assign P2_U4047 = P2_U6110 & P2_U6109 & P2_U6111; 
assign P2_U4049 = P2_U6116 & P2_U6115 & P2_U6117; 
assign P2_U4617 = ~(P2_U4616 & P2_U3269); 
assign P2_U5673 = ~P2_U3535; 
assign P2_U6123 = ~(P2_U2372 & P2_R2099_U73); 
assign P2_U6433 = ~(P2_ADD_391_1196_U98 & P2_U2397); 
assign P2_U6562 = ~(P2_U2379 & P2_R2099_U73); 
assign P2_U6822 = ~(P2_U2392 & P2_R2099_U73); 
assign P2_R2099_U169 = ~(P2_R2099_U146 & P2_R2099_U101); 
assign P2_ADD_391_1196_U130 = ~(P2_ADD_391_1196_U266 & P2_ADD_391_1196_U265); 
assign P2_ADD_391_1196_U385 = ~(P2_ADD_391_1196_U263 & P2_ADD_391_1196_U383); 
assign P2_R2278_U5 = P2_R2278_U161 & P2_R2278_U309 & P2_R2278_U206; 
assign P2_R2278_U93 = ~(P2_R2278_U422 & P2_R2278_U421); 
assign P2_R2278_U94 = ~(P2_R2278_U429 & P2_R2278_U428); 
assign P2_R2278_U95 = ~(P2_R2278_U436 & P2_R2278_U435); 
assign P2_R2278_U305 = ~P2_R2278_U163; 
assign P2_R2278_U407 = ~(P2_R2278_U162 & P2_R2278_U163); 
assign P2_U2368 = P2_U2363 & P2_U4420; 
assign P2_U2386 = P2_U2363 & P2_U4436; 
assign P2_U2388 = P2_U2363 & P2_U5675; 
assign P2_U2389 = P2_U2363 & P2_U5677; 
assign P2_U2390 = P2_U2363 & P2_U5679; 
assign P2_U2825 = ~(P2_U6819 & P2_U6821 & P2_U4166 & P2_U6822 & P2_U6820); 
assign P2_U2857 = ~(P2_U6562 & P2_U6563 & P2_U6561); 
assign P2_U2895 = ~(P2_U6432 & P2_U6431 & P2_U6435 & P2_U6434 & P2_U6433); 
assign P2_U2988 = ~(P2_U4044 & P2_U4043); 
assign P2_U2989 = ~(P2_U4042 & P2_U4041); 
assign P2_U2990 = ~(P2_U4040 & P2_U4039); 
assign P2_U2991 = ~(P2_U4038 & P2_U4037); 
assign P2_U2992 = ~(P2_U4036 & P2_U4035); 
assign P2_U2993 = ~(P2_U4034 & P2_U4033); 
assign P2_U2994 = ~(P2_U4032 & P2_U4031); 
assign P2_U2995 = ~(P2_U4030 & P2_U4029); 
assign P2_U2996 = ~(P2_U4028 & P2_U4027); 
assign P2_U2997 = ~(P2_U4026 & P2_U4025); 
assign P2_U2998 = ~(P2_U4024 & P2_U4023); 
assign P2_U2999 = ~(P2_U4022 & P2_U4021); 
assign P2_U3000 = ~(P2_U4020 & P2_U4019); 
assign P2_U3001 = ~(P2_U4018 & P2_U4017); 
assign P2_U3002 = ~(P2_U4016 & P2_U4015); 
assign P2_U3003 = ~(P2_U4014 & P2_U4013); 
assign P2_U3004 = ~(P2_U4012 & P2_U4011); 
assign P2_U3005 = ~(P2_U4010 & P2_U4009); 
assign P2_U3006 = ~(P2_U4008 & P2_U4007); 
assign P2_U3007 = ~(P2_U4006 & P2_U4005); 
assign P2_U3008 = ~(P2_U4004 & P2_U4003); 
assign P2_U3009 = ~(P2_U4002 & P2_U4001); 
assign P2_U3010 = ~(P2_U4000 & P2_U3999); 
assign P2_U3011 = ~(P2_U3998 & P2_U3997); 
assign P2_U3012 = ~(P2_U3996 & P2_U3995); 
assign P2_U3013 = ~(P2_U3994 & P2_U3993); 
assign P2_U3014 = ~(P2_U3992 & P2_U3991); 
assign P2_U4051 = P2_U6122 & P2_U6121 & P2_U6123; 
assign P2_U5686 = ~(P2_U2381 & P2_REIP_REG_0__SCAN_IN); 
assign P2_U5687 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_0__SCAN_IN); 
assign P2_U5694 = ~(P2_U2381 & P2_REIP_REG_1__SCAN_IN); 
assign P2_U5695 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_1__SCAN_IN); 
assign P2_U5702 = ~(P2_U2381 & P2_REIP_REG_2__SCAN_IN); 
assign P2_U5703 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_2__SCAN_IN); 
assign P2_U5710 = ~(P2_U2381 & P2_REIP_REG_3__SCAN_IN); 
assign P2_U5711 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_3__SCAN_IN); 
assign P2_U5718 = ~(P2_U2381 & P2_REIP_REG_4__SCAN_IN); 
assign P2_U5719 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_4__SCAN_IN); 
assign P2_U5726 = ~(P2_U2381 & P2_REIP_REG_5__SCAN_IN); 
assign P2_U5727 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_5__SCAN_IN); 
assign P2_U5734 = ~(P2_U2381 & P2_REIP_REG_6__SCAN_IN); 
assign P2_U5735 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_6__SCAN_IN); 
assign P2_U5742 = ~(P2_U2381 & P2_REIP_REG_7__SCAN_IN); 
assign P2_U5743 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_7__SCAN_IN); 
assign P2_U5750 = ~(P2_U2381 & P2_REIP_REG_8__SCAN_IN); 
assign P2_U5751 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_8__SCAN_IN); 
assign P2_U5758 = ~(P2_U2381 & P2_REIP_REG_9__SCAN_IN); 
assign P2_U5759 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_9__SCAN_IN); 
assign P2_U5766 = ~(P2_U2381 & P2_REIP_REG_10__SCAN_IN); 
assign P2_U5767 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_10__SCAN_IN); 
assign P2_U5774 = ~(P2_U2381 & P2_REIP_REG_11__SCAN_IN); 
assign P2_U5775 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_11__SCAN_IN); 
assign P2_U5782 = ~(P2_U2381 & P2_REIP_REG_12__SCAN_IN); 
assign P2_U5783 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_12__SCAN_IN); 
assign P2_U5790 = ~(P2_U2381 & P2_REIP_REG_13__SCAN_IN); 
assign P2_U5791 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_13__SCAN_IN); 
assign P2_U5798 = ~(P2_U2381 & P2_REIP_REG_14__SCAN_IN); 
assign P2_U5799 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_14__SCAN_IN); 
assign P2_U5806 = ~(P2_U2381 & P2_REIP_REG_15__SCAN_IN); 
assign P2_U5807 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_15__SCAN_IN); 
assign P2_U5814 = ~(P2_U2381 & P2_REIP_REG_16__SCAN_IN); 
assign P2_U5815 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_16__SCAN_IN); 
assign P2_U5822 = ~(P2_U2381 & P2_REIP_REG_17__SCAN_IN); 
assign P2_U5823 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_17__SCAN_IN); 
assign P2_U5830 = ~(P2_U2381 & P2_REIP_REG_18__SCAN_IN); 
assign P2_U5831 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_18__SCAN_IN); 
assign P2_U5838 = ~(P2_U2381 & P2_REIP_REG_19__SCAN_IN); 
assign P2_U5839 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_19__SCAN_IN); 
assign P2_U5846 = ~(P2_U2381 & P2_REIP_REG_20__SCAN_IN); 
assign P2_U5847 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_20__SCAN_IN); 
assign P2_U5854 = ~(P2_U2381 & P2_REIP_REG_21__SCAN_IN); 
assign P2_U5855 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_21__SCAN_IN); 
assign P2_U5862 = ~(P2_U2381 & P2_REIP_REG_22__SCAN_IN); 
assign P2_U5863 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_22__SCAN_IN); 
assign P2_U5870 = ~(P2_U2381 & P2_REIP_REG_23__SCAN_IN); 
assign P2_U5871 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_23__SCAN_IN); 
assign P2_U5878 = ~(P2_U2381 & P2_REIP_REG_24__SCAN_IN); 
assign P2_U5879 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_24__SCAN_IN); 
assign P2_U5886 = ~(P2_U2381 & P2_REIP_REG_25__SCAN_IN); 
assign P2_U5887 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_25__SCAN_IN); 
assign P2_U5894 = ~(P2_U2381 & P2_REIP_REG_26__SCAN_IN); 
assign P2_U5895 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_26__SCAN_IN); 
assign P2_U5902 = ~(P2_U2381 & P2_REIP_REG_27__SCAN_IN); 
assign P2_U5903 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_27__SCAN_IN); 
assign P2_U5910 = ~(P2_U2381 & P2_REIP_REG_28__SCAN_IN); 
assign P2_U5911 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_28__SCAN_IN); 
assign P2_U5918 = ~(P2_U2381 & P2_REIP_REG_29__SCAN_IN); 
assign P2_U5919 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_29__SCAN_IN); 
assign P2_U5926 = ~(P2_U2381 & P2_REIP_REG_30__SCAN_IN); 
assign P2_U5927 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_30__SCAN_IN); 
assign P2_U5934 = ~(P2_U2381 & P2_REIP_REG_31__SCAN_IN); 
assign P2_U5935 = ~(P2_U5673 & P2_INSTADDRPOINTER_REG_31__SCAN_IN); 
assign P2_U6107 = ~(P2_U2370 & P2_R2278_U95); 
assign P2_U6113 = ~(P2_U2370 & P2_R2278_U94); 
assign P2_U6119 = ~(P2_U2370 & P2_R2278_U93); 
assign P2_U6131 = ~(P2_U2370 & P2_R2278_U5); 
assign P2_U8057 = ~(P2_U4617 & P2_STATE2_REG_0__SCAN_IN); 
assign P2_R2099_U72 = ~(P2_R2099_U169 & P2_R2099_U168); 
assign P2_ADD_391_1196_U97 = ~(P2_ADD_391_1196_U385 & P2_ADD_391_1196_U384); 
assign P2_ADD_391_1196_U267 = ~P2_ADD_391_1196_U130; 
assign P2_ADD_391_1196_U269 = ~(P2_ADD_391_1196_U268 & P2_ADD_391_1196_U130); 
assign P2_ADD_391_1196_U377 = ~(P2_ADD_391_1196_U129 & P2_ADD_391_1196_U130); 
assign P2_R2278_U408 = ~(P2_R2278_U305 & P2_R2278_U406); 
assign P2_U2384 = P2_U2368 & P2_U4417; 
assign P2_U2385 = P2_U2368 & P2_U4428; 
assign P2_U3898 = P2_U5687 & P2_U5686; 
assign P2_U3901 = P2_U5695 & P2_U5694; 
assign P2_U3904 = P2_U5703 & P2_U5702; 
assign P2_U3907 = P2_U5711 & P2_U5710; 
assign P2_U3910 = P2_U5719 & P2_U5718; 
assign P2_U3913 = P2_U5727 & P2_U5726; 
assign P2_U3916 = P2_U5735 & P2_U5734; 
assign P2_U3919 = P2_U5743 & P2_U5742; 
assign P2_U3922 = P2_U5751 & P2_U5750; 
assign P2_U3925 = P2_U5759 & P2_U5758; 
assign P2_U3928 = P2_U5767 & P2_U5766; 
assign P2_U3931 = P2_U5775 & P2_U5774; 
assign P2_U3934 = P2_U5783 & P2_U5782; 
assign P2_U3937 = P2_U5791 & P2_U5790; 
assign P2_U3940 = P2_U5799 & P2_U5798; 
assign P2_U3943 = P2_U5807 & P2_U5806; 
assign P2_U3946 = P2_U5815 & P2_U5814; 
assign P2_U3949 = P2_U5823 & P2_U5822; 
assign P2_U3952 = P2_U5831 & P2_U5830; 
assign P2_U3955 = P2_U5839 & P2_U5838; 
assign P2_U3958 = P2_U5847 & P2_U5846; 
assign P2_U3961 = P2_U5855 & P2_U5854; 
assign P2_U3964 = P2_U5863 & P2_U5862; 
assign P2_U3967 = P2_U5871 & P2_U5870; 
assign P2_U3970 = P2_U5879 & P2_U5878; 
assign P2_U3973 = P2_U5887 & P2_U5886; 
assign P2_U3976 = P2_U5895 & P2_U5894; 
assign P2_U3979 = P2_U5903 & P2_U5902; 
assign P2_U3982 = P2_U5911 & P2_U5910; 
assign P2_U3984 = P2_U5919 & P2_U5918; 
assign P2_U3986 = P2_U5927 & P2_U5926; 
assign P2_U3988 = P2_U5935 & P2_U5934; 
assign P2_U4046 = P2_U6107 & P2_U6106 & P2_U6108; 
assign P2_U4048 = P2_U6113 & P2_U6112 & P2_U6114; 
assign P2_U4050 = P2_U6119 & P2_U6118 & P2_U6120; 
assign P2_U4054 = P2_U6131 & P2_U6130 & P2_U6132; 
assign P2_U4619 = ~(P2_U8057 & P2_U8056 & P2_U3715); 
assign P2_U5680 = ~(P2_U2390 & P2_R2096_U68); 
assign P2_U5681 = ~(P2_U2389 & P2_R2099_U94); 
assign P2_U5682 = ~(P2_R2027_U5 & P2_U2388); 
assign P2_U5683 = ~(P2_ADD_394_U4 & P2_U2386); 
assign P2_U5688 = ~(P2_U2390 & P2_R2096_U51); 
assign P2_U5689 = ~(P2_U2389 & P2_R2099_U5); 
assign P2_U5690 = ~(P2_R2027_U85 & P2_U2388); 
assign P2_U5691 = ~(P2_ADD_394_U85 & P2_U2386); 
assign P2_U5696 = ~(P2_U2390 & P2_R2096_U77); 
assign P2_U5697 = ~(P2_U2389 & P2_R2099_U96); 
assign P2_U5698 = ~(P2_R2027_U74 & P2_U2388); 
assign P2_U5699 = ~(P2_ADD_394_U5 & P2_U2386); 
assign P2_U5704 = ~(P2_U2390 & P2_R2096_U75); 
assign P2_U5705 = ~(P2_U2389 & P2_R2099_U95); 
assign P2_U5706 = ~(P2_R2027_U71 & P2_U2388); 
assign P2_U5707 = ~(P2_ADD_394_U95 & P2_U2386); 
assign P2_U5712 = ~(P2_R2096_U74 & P2_U2390); 
assign P2_U5713 = ~(P2_R2099_U98 & P2_U2389); 
assign P2_U5714 = ~(P2_R2027_U70 & P2_U2388); 
assign P2_U5715 = ~(P2_ADD_394_U76 & P2_U2386); 
assign P2_U5720 = ~(P2_R2096_U73 & P2_U2390); 
assign P2_U5721 = ~(P2_R2099_U71 & P2_U2389); 
assign P2_U5722 = ~(P2_R2027_U69 & P2_U2388); 
assign P2_U5723 = ~(P2_ADD_394_U79 & P2_U2386); 
assign P2_U5728 = ~(P2_R2096_U72 & P2_U2390); 
assign P2_U5729 = ~(P2_R2099_U70 & P2_U2389); 
assign P2_U5730 = ~(P2_R2027_U68 & P2_U2388); 
assign P2_U5731 = ~(P2_ADD_394_U63 & P2_U2386); 
assign P2_U5736 = ~(P2_R2096_U71 & P2_U2390); 
assign P2_U5737 = ~(P2_R2099_U69 & P2_U2389); 
assign P2_U5738 = ~(P2_R2027_U67 & P2_U2388); 
assign P2_U5739 = ~(P2_ADD_394_U89 & P2_U2386); 
assign P2_U5744 = ~(P2_R2096_U70 & P2_U2390); 
assign P2_U5745 = ~(P2_R2099_U68 & P2_U2389); 
assign P2_U5746 = ~(P2_R2027_U66 & P2_U2388); 
assign P2_U5747 = ~(P2_ADD_394_U80 & P2_U2386); 
assign P2_U5752 = ~(P2_R2096_U69 & P2_U2390); 
assign P2_U5753 = ~(P2_R2099_U67 & P2_U2389); 
assign P2_U5754 = ~(P2_R2027_U65 & P2_U2388); 
assign P2_U5755 = ~(P2_ADD_394_U70 & P2_U2386); 
assign P2_U5760 = ~(P2_R2096_U97 & P2_U2390); 
assign P2_U5761 = ~(P2_R2099_U93 & P2_U2389); 
assign P2_U5762 = ~(P2_R2027_U95 & P2_U2388); 
assign P2_U5763 = ~(P2_ADD_394_U83 & P2_U2386); 
assign P2_U5768 = ~(P2_R2096_U96 & P2_U2390); 
assign P2_U5769 = ~(P2_R2099_U92 & P2_U2389); 
assign P2_U5770 = ~(P2_R2027_U94 & P2_U2388); 
assign P2_U5771 = ~(P2_ADD_394_U73 & P2_U2386); 
assign P2_U5776 = ~(P2_R2096_U95 & P2_U2390); 
assign P2_U5777 = ~(P2_R2099_U91 & P2_U2389); 
assign P2_U5778 = ~(P2_R2027_U93 & P2_U2388); 
assign P2_U5779 = ~(P2_ADD_394_U88 & P2_U2386); 
assign P2_U5784 = ~(P2_R2096_U94 & P2_U2390); 
assign P2_U5785 = ~(P2_R2099_U90 & P2_U2389); 
assign P2_U5786 = ~(P2_R2027_U92 & P2_U2388); 
assign P2_U5787 = ~(P2_ADD_394_U69 & P2_U2386); 
assign P2_U5792 = ~(P2_R2096_U93 & P2_U2390); 
assign P2_U5793 = ~(P2_R2099_U89 & P2_U2389); 
assign P2_U5794 = ~(P2_R2027_U91 & P2_U2388); 
assign P2_U5795 = ~(P2_ADD_394_U78 & P2_U2386); 
assign P2_U5800 = ~(P2_R2096_U92 & P2_U2390); 
assign P2_U5801 = ~(P2_R2099_U88 & P2_U2389); 
assign P2_U5802 = ~(P2_R2027_U90 & P2_U2388); 
assign P2_U5803 = ~(P2_ADD_394_U75 & P2_U2386); 
assign P2_U5808 = ~(P2_R2096_U91 & P2_U2390); 
assign P2_U5809 = ~(P2_R2099_U87 & P2_U2389); 
assign P2_U5810 = ~(P2_R2027_U89 & P2_U2388); 
assign P2_U5811 = ~(P2_ADD_394_U91 & P2_U2386); 
assign P2_U5816 = ~(P2_R2096_U90 & P2_U2390); 
assign P2_U5817 = ~(P2_R2099_U86 & P2_U2389); 
assign P2_U5818 = ~(P2_R2027_U88 & P2_U2388); 
assign P2_U5819 = ~(P2_ADD_394_U67 & P2_U2386); 
assign P2_U5824 = ~(P2_R2096_U89 & P2_U2390); 
assign P2_U5825 = ~(P2_R2099_U85 & P2_U2389); 
assign P2_U5826 = ~(P2_R2027_U87 & P2_U2388); 
assign P2_U5827 = ~(P2_ADD_394_U72 & P2_U2386); 
assign P2_U5832 = ~(P2_R2096_U88 & P2_U2390); 
assign P2_U5833 = ~(P2_R2099_U84 & P2_U2389); 
assign P2_U5834 = ~(P2_R2027_U86 & P2_U2388); 
assign P2_U5835 = ~(P2_ADD_394_U82 & P2_U2386); 
assign P2_U5840 = ~(P2_R2096_U87 & P2_U2390); 
assign P2_U5841 = ~(P2_R2099_U83 & P2_U2389); 
assign P2_U5842 = ~(P2_R2027_U84 & P2_U2388); 
assign P2_U5843 = ~(P2_ADD_394_U68 & P2_U2386); 
assign P2_U5848 = ~(P2_R2096_U86 & P2_U2390); 
assign P2_U5849 = ~(P2_R2099_U82 & P2_U2389); 
assign P2_U5850 = ~(P2_R2027_U83 & P2_U2388); 
assign P2_U5851 = ~(P2_ADD_394_U87 & P2_U2386); 
assign P2_U5856 = ~(P2_R2096_U85 & P2_U2390); 
assign P2_U5857 = ~(P2_R2099_U81 & P2_U2389); 
assign P2_U5858 = ~(P2_R2027_U82 & P2_U2388); 
assign P2_U5859 = ~(P2_ADD_394_U71 & P2_U2386); 
assign P2_U5864 = ~(P2_R2096_U84 & P2_U2390); 
assign P2_U5865 = ~(P2_R2099_U80 & P2_U2389); 
assign P2_U5866 = ~(P2_R2027_U81 & P2_U2388); 
assign P2_U5867 = ~(P2_ADD_394_U81 & P2_U2386); 
assign P2_U5872 = ~(P2_R2096_U83 & P2_U2390); 
assign P2_U5873 = ~(P2_R2099_U79 & P2_U2389); 
assign P2_U5874 = ~(P2_R2027_U80 & P2_U2388); 
assign P2_U5875 = ~(P2_ADD_394_U66 & P2_U2386); 
assign P2_U5880 = ~(P2_R2096_U82 & P2_U2390); 
assign P2_U5881 = ~(P2_R2099_U78 & P2_U2389); 
assign P2_U5882 = ~(P2_R2027_U79 & P2_U2388); 
assign P2_U5883 = ~(P2_ADD_394_U90 & P2_U2386); 
assign P2_U5888 = ~(P2_R2096_U81 & P2_U2390); 
assign P2_U5889 = ~(P2_R2099_U77 & P2_U2389); 
assign P2_U5890 = ~(P2_R2027_U78 & P2_U2388); 
assign P2_U5891 = ~(P2_ADD_394_U74 & P2_U2386); 
assign P2_U5896 = ~(P2_R2096_U80 & P2_U2390); 
assign P2_U5897 = ~(P2_R2099_U76 & P2_U2389); 
assign P2_U5898 = ~(P2_R2027_U77 & P2_U2388); 
assign P2_U5899 = ~(P2_ADD_394_U77 & P2_U2386); 
assign P2_U5904 = ~(P2_R2096_U79 & P2_U2390); 
assign P2_U5905 = ~(P2_R2099_U75 & P2_U2389); 
assign P2_U5906 = ~(P2_R2027_U76 & P2_U2388); 
assign P2_U5907 = ~(P2_ADD_394_U86 & P2_U2386); 
assign P2_U5912 = ~(P2_R2096_U78 & P2_U2390); 
assign P2_U5913 = ~(P2_R2099_U74 & P2_U2389); 
assign P2_U5914 = ~(P2_R2027_U75 & P2_U2388); 
assign P2_U5915 = ~(P2_ADD_394_U65 & P2_U2386); 
assign P2_U5920 = ~(P2_R2096_U76 & P2_U2390); 
assign P2_U5921 = ~(P2_R2099_U73 & P2_U2389); 
assign P2_U5922 = ~(P2_R2027_U73 & P2_U2388); 
assign P2_U5923 = ~(P2_ADD_394_U64 & P2_U2386); 
assign P2_U5928 = ~(P2_R2096_U50 & P2_U2390); 
assign P2_U5929 = ~(P2_R2099_U72 & P2_U2389); 
assign P2_U5930 = ~(P2_R2027_U72 & P2_U2388); 
assign P2_U5931 = ~(P2_ADD_394_U84 & P2_U2386); 
assign P2_U6129 = ~(P2_U2372 & P2_R2099_U72); 
assign P2_U6438 = ~(P2_ADD_391_1196_U97 & P2_U2397); 
assign P2_U6564 = ~(P2_U2379 & P2_R2099_U72); 
assign P2_U6830 = ~(P2_U2392 & P2_R2099_U72); 
assign P2_ADD_391_1196_U128 = ~(P2_ADD_391_1196_U270 & P2_ADD_391_1196_U269); 
assign P2_ADD_391_1196_U378 = ~(P2_ADD_391_1196_U267 & P2_ADD_391_1196_U376); 
assign P2_R2278_U91 = ~(P2_R2278_U408 & P2_R2278_U407); 
assign P2_U2824 = ~(P2_U6827 & P2_U6829 & P2_U4168 & P2_U6830 & P2_U6828); 
assign P2_U2856 = ~(P2_U6565 & P2_U6564); 
assign P2_U2894 = ~(P2_U6437 & P2_U6436 & P2_U6440 & P2_U6439 & P2_U6438); 
assign P2_U2985 = ~(P2_U4050 & P2_U4049); 
assign P2_U2986 = ~(P2_U4048 & P2_U4047); 
assign P2_U2987 = ~(P2_U4046 & P2_U4045); 
assign P2_U3299 = ~(P2_U4619 & P2_STATE2_REG_0__SCAN_IN); 
assign P2_U3896 = P2_U5681 & P2_U5680; 
assign P2_U3897 = P2_U5683 & P2_U5682; 
assign P2_U3899 = P2_U5689 & P2_U5688; 
assign P2_U3900 = P2_U5691 & P2_U5690; 
assign P2_U3902 = P2_U5697 & P2_U5696; 
assign P2_U3903 = P2_U5699 & P2_U5698; 
assign P2_U3905 = P2_U5705 & P2_U5704; 
assign P2_U3906 = P2_U5707 & P2_U5706; 
assign P2_U3908 = P2_U5713 & P2_U5712; 
assign P2_U3909 = P2_U5715 & P2_U5714; 
assign P2_U3911 = P2_U5721 & P2_U5720; 
assign P2_U3912 = P2_U5723 & P2_U5722; 
assign P2_U3914 = P2_U5729 & P2_U5728; 
assign P2_U3915 = P2_U5731 & P2_U5730; 
assign P2_U3917 = P2_U5737 & P2_U5736; 
assign P2_U3918 = P2_U5739 & P2_U5738; 
assign P2_U3920 = P2_U5745 & P2_U5744; 
assign P2_U3921 = P2_U5747 & P2_U5746; 
assign P2_U3923 = P2_U5753 & P2_U5752; 
assign P2_U3924 = P2_U5755 & P2_U5754; 
assign P2_U3926 = P2_U5761 & P2_U5760; 
assign P2_U3927 = P2_U5763 & P2_U5762; 
assign P2_U3929 = P2_U5769 & P2_U5768; 
assign P2_U3930 = P2_U5771 & P2_U5770; 
assign P2_U3932 = P2_U5777 & P2_U5776; 
assign P2_U3933 = P2_U5779 & P2_U5778; 
assign P2_U3935 = P2_U5785 & P2_U5784; 
assign P2_U3936 = P2_U5787 & P2_U5786; 
assign P2_U3938 = P2_U5793 & P2_U5792; 
assign P2_U3939 = P2_U5795 & P2_U5794; 
assign P2_U3941 = P2_U5801 & P2_U5800; 
assign P2_U3942 = P2_U5803 & P2_U5802; 
assign P2_U3944 = P2_U5809 & P2_U5808; 
assign P2_U3945 = P2_U5811 & P2_U5810; 
assign P2_U3947 = P2_U5817 & P2_U5816; 
assign P2_U3948 = P2_U5819 & P2_U5818; 
assign P2_U3950 = P2_U5825 & P2_U5824; 
assign P2_U3951 = P2_U5827 & P2_U5826; 
assign P2_U3953 = P2_U5833 & P2_U5832; 
assign P2_U3954 = P2_U5835 & P2_U5834; 
assign P2_U3956 = P2_U5841 & P2_U5840; 
assign P2_U3957 = P2_U5843 & P2_U5842; 
assign P2_U3959 = P2_U5849 & P2_U5848; 
assign P2_U3960 = P2_U5851 & P2_U5850; 
assign P2_U3962 = P2_U5857 & P2_U5856; 
assign P2_U3963 = P2_U5859 & P2_U5858; 
assign P2_U3965 = P2_U5865 & P2_U5864; 
assign P2_U3966 = P2_U5867 & P2_U5866; 
assign P2_U3968 = P2_U5873 & P2_U5872; 
assign P2_U3969 = P2_U5875 & P2_U5874; 
assign P2_U3971 = P2_U5881 & P2_U5880; 
assign P2_U3972 = P2_U5883 & P2_U5882; 
assign P2_U3974 = P2_U5889 & P2_U5888; 
assign P2_U3975 = P2_U5891 & P2_U5890; 
assign P2_U3977 = P2_U5897 & P2_U5896; 
assign P2_U3978 = P2_U5899 & P2_U5898; 
assign P2_U3980 = P2_U5905 & P2_U5904; 
assign P2_U3981 = P2_U5907 & P2_U5906; 
assign P2_U3983 = P2_U5915 & P2_U5914 & P2_U5913 & P2_U5912; 
assign P2_U3985 = P2_U5923 & P2_U5922 & P2_U5921; 
assign P2_U3987 = P2_U5931 & P2_U5930 & P2_U5929; 
assign P2_U4053 = P2_U6128 & P2_U6127 & P2_U6129; 
assign P2_U4626 = ~(P2_U4619 & P2_U4465); 
assign P2_U4629 = ~(P2_U2374 & P2_U4619); 
assign P2_U4631 = ~(P2_U4619 & P2_U4464); 
assign P2_U5684 = ~(P2_R2278_U83 & P2_U2385); 
assign P2_U5685 = ~(P2_ADD_371_1212_U68 & P2_U2384); 
assign P2_U5692 = ~(P2_R2278_U6 & P2_U2385); 
assign P2_U5693 = ~(P2_ADD_371_1212_U25 & P2_U2384); 
assign P2_U5700 = ~(P2_R2278_U92 & P2_U2385); 
assign P2_U5701 = ~(P2_ADD_371_1212_U79 & P2_U2384); 
assign P2_U5708 = ~(P2_R2278_U90 & P2_U2385); 
assign P2_U5709 = ~(P2_ADD_371_1212_U84 & P2_U2384); 
assign P2_U5716 = ~(P2_R2278_U89 & P2_U2385); 
assign P2_U5717 = ~(P2_ADD_371_1212_U80 & P2_U2384); 
assign P2_U5724 = ~(P2_R2278_U88 & P2_U2385); 
assign P2_U5725 = ~(P2_ADD_371_1212_U81 & P2_U2384); 
assign P2_U5732 = ~(P2_R2278_U87 & P2_U2385); 
assign P2_U5733 = ~(P2_ADD_371_1212_U78 & P2_U2384); 
assign P2_U5740 = ~(P2_R2278_U86 & P2_U2385); 
assign P2_U5741 = ~(P2_ADD_371_1212_U85 & P2_U2384); 
assign P2_U5748 = ~(P2_R2278_U85 & P2_U2385); 
assign P2_U5749 = ~(P2_ADD_371_1212_U82 & P2_U2384); 
assign P2_U5756 = ~(P2_R2278_U84 & P2_U2385); 
assign P2_U5757 = ~(P2_ADD_371_1212_U118 & P2_U2384); 
assign P2_U5764 = ~(P2_R2278_U112 & P2_U2385); 
assign P2_U5765 = ~(P2_ADD_371_1212_U13 & P2_U2384); 
assign P2_U5772 = ~(P2_R2278_U111 & P2_U2385); 
assign P2_U5773 = ~(P2_ADD_371_1212_U14 & P2_U2384); 
assign P2_U5780 = ~(P2_R2278_U110 & P2_U2385); 
assign P2_U5781 = ~(P2_ADD_371_1212_U76 & P2_U2384); 
assign P2_U5788 = ~(P2_R2278_U109 & P2_U2385); 
assign P2_U5789 = ~(P2_ADD_371_1212_U15 & P2_U2384); 
assign P2_U5796 = ~(P2_R2278_U108 & P2_U2385); 
assign P2_U5797 = ~(P2_ADD_371_1212_U16 & P2_U2384); 
assign P2_U5804 = ~(P2_R2278_U107 & P2_U2385); 
assign P2_U5805 = ~(P2_ADD_371_1212_U73 & P2_U2384); 
assign P2_U5812 = ~(P2_R2278_U106 & P2_U2385); 
assign P2_U5813 = ~(P2_ADD_371_1212_U17 & P2_U2384); 
assign P2_U5820 = ~(P2_R2278_U105 & P2_U2385); 
assign P2_U5821 = ~(P2_ADD_371_1212_U71 & P2_U2384); 
assign P2_U5828 = ~(P2_R2278_U104 & P2_U2385); 
assign P2_U5829 = ~(P2_ADD_371_1212_U72 & P2_U2384); 
assign P2_U5836 = ~(P2_R2278_U103 & P2_U2385); 
assign P2_U5837 = ~(P2_ADD_371_1212_U18 & P2_U2384); 
assign P2_U5844 = ~(P2_R2278_U102 & P2_U2385); 
assign P2_U5845 = ~(P2_ADD_371_1212_U19 & P2_U2384); 
assign P2_U5852 = ~(P2_R2278_U101 & P2_U2385); 
assign P2_U5853 = ~(P2_ADD_371_1212_U75 & P2_U2384); 
assign P2_U5860 = ~(P2_R2278_U100 & P2_U2385); 
assign P2_U5861 = ~(P2_ADD_371_1212_U20 & P2_U2384); 
assign P2_U5868 = ~(P2_R2278_U99 & P2_U2385); 
assign P2_U5869 = ~(P2_ADD_371_1212_U21 & P2_U2384); 
assign P2_U5876 = ~(P2_R2278_U98 & P2_U2385); 
assign P2_U5877 = ~(P2_ADD_371_1212_U70 & P2_U2384); 
assign P2_U5884 = ~(P2_R2278_U97 & P2_U2385); 
assign P2_U5885 = ~(P2_ADD_371_1212_U77 & P2_U2384); 
assign P2_U5892 = ~(P2_R2278_U96 & P2_U2385); 
assign P2_U5893 = ~(P2_ADD_371_1212_U22 & P2_U2384); 
assign P2_U5900 = ~(P2_R2278_U95 & P2_U2385); 
assign P2_U5901 = ~(P2_ADD_371_1212_U74 & P2_U2384); 
assign P2_U5908 = ~(P2_R2278_U94 & P2_U2385); 
assign P2_U5909 = ~(P2_ADD_371_1212_U23 & P2_U2384); 
assign P2_U5916 = ~(P2_R2278_U93 & P2_U2385); 
assign P2_U5917 = ~(P2_ADD_371_1212_U24 & P2_U2384); 
assign P2_U5924 = ~(P2_R2278_U91 & P2_U2385); 
assign P2_U5925 = ~(P2_ADD_371_1212_U69 & P2_U2384); 
assign P2_U5932 = ~(P2_R2278_U5 & P2_U2385); 
assign P2_U5933 = ~(P2_ADD_371_1212_U83 & P2_U2384); 
assign P2_U6125 = ~(P2_U2370 & P2_R2278_U91); 
assign P2_U8061 = ~(P2_U4630 & P2_U4619 & P2_U3284); 
assign P2_ADD_391_1196_U96 = ~(P2_ADD_391_1196_U378 & P2_ADD_391_1196_U377); 
assign P2_ADD_391_1196_U271 = ~P2_ADD_391_1196_U128; 
assign P2_ADD_391_1196_U273 = ~(P2_ADD_391_1196_U272 & P2_ADD_391_1196_U128); 
assign P2_ADD_391_1196_U370 = ~(P2_ADD_391_1196_U127 & P2_ADD_391_1196_U128); 
assign P2_U2983 = ~(P2_U4054 & P2_U4053); 
assign P2_U3015 = ~(P2_U5933 & P2_U5932 & P2_U3988 & P2_U3987 & P2_U5928); 
assign P2_U3016 = ~(P2_U5925 & P2_U5924 & P2_U3986 & P2_U3985 & P2_U5920); 
assign P2_U3017 = ~(P2_U5917 & P2_U5916 & P2_U3984 & P2_U3983); 
assign P2_U3018 = ~(P2_U5909 & P2_U5908 & P2_U3982 & P2_U3981 & P2_U3980); 
assign P2_U3019 = ~(P2_U5901 & P2_U5900 & P2_U3979 & P2_U3978 & P2_U3977); 
assign P2_U3020 = ~(P2_U5893 & P2_U5892 & P2_U3976 & P2_U3975 & P2_U3974); 
assign P2_U3021 = ~(P2_U5885 & P2_U5884 & P2_U3973 & P2_U3972 & P2_U3971); 
assign P2_U3022 = ~(P2_U5877 & P2_U5876 & P2_U3970 & P2_U3969 & P2_U3968); 
assign P2_U3023 = ~(P2_U5869 & P2_U5868 & P2_U3967 & P2_U3966 & P2_U3965); 
assign P2_U3024 = ~(P2_U5861 & P2_U5860 & P2_U3964 & P2_U3963 & P2_U3962); 
assign P2_U3025 = ~(P2_U5853 & P2_U5852 & P2_U3961 & P2_U3960 & P2_U3959); 
assign P2_U3026 = ~(P2_U5845 & P2_U5844 & P2_U3958 & P2_U3957 & P2_U3956); 
assign P2_U3027 = ~(P2_U5837 & P2_U5836 & P2_U3955 & P2_U3954 & P2_U3953); 
assign P2_U3028 = ~(P2_U5829 & P2_U5828 & P2_U3952 & P2_U3951 & P2_U3950); 
assign P2_U3029 = ~(P2_U5821 & P2_U5820 & P2_U3949 & P2_U3948 & P2_U3947); 
assign P2_U3030 = ~(P2_U5813 & P2_U5812 & P2_U3946 & P2_U3945 & P2_U3944); 
assign P2_U3031 = ~(P2_U5805 & P2_U5804 & P2_U3943 & P2_U3942 & P2_U3941); 
assign P2_U3032 = ~(P2_U5797 & P2_U5796 & P2_U3940 & P2_U3939 & P2_U3938); 
assign P2_U3033 = ~(P2_U5789 & P2_U5788 & P2_U3937 & P2_U3936 & P2_U3935); 
assign P2_U3034 = ~(P2_U5781 & P2_U5780 & P2_U3934 & P2_U3933 & P2_U3932); 
assign P2_U3035 = ~(P2_U5773 & P2_U5772 & P2_U3931 & P2_U3930 & P2_U3929); 
assign P2_U3036 = ~(P2_U5765 & P2_U5764 & P2_U3928 & P2_U3927 & P2_U3926); 
assign P2_U3037 = ~(P2_U5757 & P2_U5756 & P2_U3925 & P2_U3924 & P2_U3923); 
assign P2_U3038 = ~(P2_U5749 & P2_U5748 & P2_U3922 & P2_U3921 & P2_U3920); 
assign P2_U3039 = ~(P2_U5741 & P2_U5740 & P2_U3919 & P2_U3918 & P2_U3917); 
assign P2_U3040 = ~(P2_U5733 & P2_U5732 & P2_U3916 & P2_U3915 & P2_U3914); 
assign P2_U3041 = ~(P2_U5725 & P2_U5724 & P2_U3913 & P2_U3912 & P2_U3911); 
assign P2_U3042 = ~(P2_U5717 & P2_U5716 & P2_U3910 & P2_U3909 & P2_U3908); 
assign P2_U3043 = ~(P2_U5709 & P2_U5708 & P2_U3907 & P2_U3906 & P2_U3905); 
assign P2_U3044 = ~(P2_U5701 & P2_U5700 & P2_U3904 & P2_U3903 & P2_U3902); 
assign P2_U3045 = ~(P2_U5693 & P2_U5692 & P2_U3901 & P2_U3900 & P2_U3899); 
assign P2_U3046 = ~(P2_U5685 & P2_U5684 & P2_U3898 & P2_U3897 & P2_U3896); 
assign P2_U4052 = P2_U6126 & P2_U6124 & P2_U6125; 
assign P2_U4620 = ~P2_U3299; 
assign P2_U4625 = ~(P2_U3299 & P2_STATE2_REG_2__SCAN_IN); 
assign P2_U4628 = ~(P2_U4626 & P2_STATE2_REG_1__SCAN_IN); 
assign P2_U6443 = ~(P2_ADD_391_1196_U96 & P2_U2397); 
assign P2_U8058 = ~(P2_U3299 & P2_STATE2_REG_3__SCAN_IN); 
assign P2_U8060 = ~(P2_U4631 & P2_STATE2_REG_0__SCAN_IN); 
assign P2_ADD_391_1196_U126 = ~(P2_ADD_391_1196_U274 & P2_ADD_391_1196_U273); 
assign P2_ADD_391_1196_U371 = ~(P2_ADD_391_1196_U271 & P2_ADD_391_1196_U369); 
assign P2_U2893 = ~(P2_U6442 & P2_U6441 & P2_U6445 & P2_U6444 & P2_U6443); 
assign P2_U2984 = ~(P2_U4052 & P2_U4051); 
assign P2_U3176 = ~(P2_U8061 & P2_U8060 & P2_U3721); 
assign P2_U3178 = ~(P2_U3716 & P2_U4625); 
assign P2_U4627 = ~(P2_U3717 & P2_U4620); 
assign P2_U8059 = ~(P2_U2448 & P2_U4620); 
assign P2_ADD_391_1196_U95 = ~(P2_ADD_391_1196_U371 & P2_ADD_391_1196_U370); 
assign P2_ADD_391_1196_U275 = ~P2_ADD_391_1196_U126; 
assign P2_ADD_391_1196_U277 = ~(P2_ADD_391_1196_U276 & P2_ADD_391_1196_U126); 
assign P2_ADD_391_1196_U363 = ~(P2_ADD_391_1196_U125 & P2_ADD_391_1196_U126); 
assign P2_U3177 = ~(P2_U4629 & P2_U4628 & P2_U4627 & P2_U4454); 
assign P2_U3593 = ~(P2_U8059 & P2_U8058); 
assign P2_U6448 = ~(P2_ADD_391_1196_U95 & P2_U2397); 
assign P2_ADD_391_1196_U82 = ~(P2_ADD_391_1196_U278 & P2_ADD_391_1196_U277); 
assign P2_ADD_391_1196_U364 = ~(P2_ADD_391_1196_U275 & P2_ADD_391_1196_U362); 
assign P2_U2892 = ~(P2_U6447 & P2_U6446 & P2_U6450 & P2_U6449 & P2_U6448); 
assign P2_ADD_391_1196_U94 = ~(P2_ADD_391_1196_U364 & P2_ADD_391_1196_U363); 
assign P2_ADD_391_1196_U279 = ~P2_ADD_391_1196_U82; 
assign P2_ADD_391_1196_U281 = ~(P2_ADD_391_1196_U280 & P2_ADD_391_1196_U82); 
assign P2_ADD_391_1196_U356 = ~(P2_ADD_391_1196_U124 & P2_ADD_391_1196_U82); 
assign P2_U6453 = ~(P2_ADD_391_1196_U94 & P2_U2397); 
assign P2_ADD_391_1196_U283 = ~(P2_ADD_391_1196_U282 & P2_ADD_391_1196_U281 & P2_ADD_391_1196_U121); 
assign P2_ADD_391_1196_U285 = ~(P2_ADD_391_1196_U279 & P2_ADD_391_1196_U284); 
assign P2_ADD_391_1196_U357 = ~(P2_ADD_391_1196_U355 & P2_ADD_391_1196_U279); 
assign P2_U2891 = ~(P2_U6452 & P2_U6451 & P2_U6455 & P2_U6454 & P2_U6453); 
assign P2_ADD_391_1196_U93 = ~(P2_ADD_391_1196_U357 & P2_ADD_391_1196_U356); 
assign P2_ADD_391_1196_U287 = ~(P2_ADD_391_1196_U286 & P2_ADD_391_1196_U285 & P2_ADD_391_1196_U343); 
assign P2_U6458 = ~(P2_ADD_391_1196_U93 & P2_U2397); 
assign P2_ADD_391_1196_U8 = P2_ADD_391_1196_U287 & P2_ADD_391_1196_U283; 
assign P2_U2890 = ~(P2_U6457 & P2_U6456 & P2_U6460 & P2_U6459 & P2_U6458); 
assign P2_U6463 = ~(P2_ADD_391_1196_U8 & P2_U2397); 
assign P2_U2889 = ~(P2_U6462 & P2_U6461 & P2_U6465 & P2_U6464 & P2_U6463); 
endmodule 
