module b09_C( D_IN_REG_0__SCAN_IN, X, D_OUT_REG_7__SCAN_IN, D_OUT_REG_6__SCAN_IN, D_OUT_REG_5__SCAN_IN, D_OUT_REG_4__SCAN_IN, D_OUT_REG_3__SCAN_IN, D_OUT_REG_2__SCAN_IN, D_OUT_REG_1__SCAN_IN, D_OUT_REG_0__SCAN_IN, OLD_REG_7__SCAN_IN, OLD_REG_6__SCAN_IN, OLD_REG_5__SCAN_IN, OLD_REG_4__SCAN_IN, OLD_REG_3__SCAN_IN, OLD_REG_2__SCAN_IN, OLD_REG_1__SCAN_IN, OLD_REG_0__SCAN_IN, Y_REG_SCAN_IN, STATO_REG_1__SCAN_IN, STATO_REG_0__SCAN_IN, D_IN_REG_8__SCAN_IN, D_IN_REG_7__SCAN_IN, D_IN_REG_6__SCAN_IN, D_IN_REG_5__SCAN_IN, D_IN_REG_4__SCAN_IN, D_IN_REG_3__SCAN_IN, D_IN_REG_2__SCAN_IN, D_IN_REG_1__SCAN_IN, U91, U92, U93, U94, U95, U96, U97, U98, U99, U100, U101, U102, U103, U104, U105, U106, U107, U108, U109, U110, U111, U112, U113, U114, U115, U116, U117, U118); 
input D_IN_REG_0__SCAN_IN, X, D_OUT_REG_7__SCAN_IN, D_OUT_REG_6__SCAN_IN, D_OUT_REG_5__SCAN_IN, D_OUT_REG_4__SCAN_IN, D_OUT_REG_3__SCAN_IN, D_OUT_REG_2__SCAN_IN, D_OUT_REG_1__SCAN_IN, D_OUT_REG_0__SCAN_IN, OLD_REG_7__SCAN_IN, OLD_REG_6__SCAN_IN, OLD_REG_5__SCAN_IN, OLD_REG_4__SCAN_IN, OLD_REG_3__SCAN_IN, OLD_REG_2__SCAN_IN, OLD_REG_1__SCAN_IN, OLD_REG_0__SCAN_IN, Y_REG_SCAN_IN, STATO_REG_1__SCAN_IN, STATO_REG_0__SCAN_IN, D_IN_REG_8__SCAN_IN, D_IN_REG_7__SCAN_IN, D_IN_REG_6__SCAN_IN, D_IN_REG_5__SCAN_IN, D_IN_REG_4__SCAN_IN, D_IN_REG_3__SCAN_IN, D_IN_REG_2__SCAN_IN, D_IN_REG_1__SCAN_IN; 
output U91, U92, U93, U94, U95, U96, U97, U98, U99, U100, U101, U102, U103, U104, U105, U106, U107, U108, U109, U110, U111, U112, U113, U114, U115, U116, U117, U118; 
wire U87, U88, U89, U90, U119, U120, U121, U122, U123, U124, U125, U126, U127, U128, U129, U130, U131, U132, U133, U134, U135, U136, U137, U138, U139, U140, U141, U142, U143, U144, U145, U146, U147, U148, U149, U150, U151, U152, U153, U154, U155, U156, U157, U158, U159, U160, U161, U162, U163, U164, U165, U166, U167, U168, U169, U170, U171, U172, U173, U174, U175, U176, U177, U178, U179, U180, U181, U182, U183, U184, U185, U186, U187, U188, U189, U190, U191, U192, U193, U194, U195, U196, U197, U198, U199, U200, U201, U202, U203, U204, U205, U206, U207, U208, U209, U210, U211, U212, U213, U214, U215, U216, U217, U218, U219, U220, U221, U222, U223, U224, U225, U226; 
assign U87 = STATO_REG_1__SCAN_IN & STATO_REG_0__SCAN_IN; 
assign U119 = ~STATO_REG_0__SCAN_IN; 
assign U120 = ~D_IN_REG_0__SCAN_IN; 
assign U121 = ~D_IN_REG_1__SCAN_IN; 
assign U122 = ~OLD_REG_0__SCAN_IN; 
assign U123 = ~D_IN_REG_2__SCAN_IN; 
assign U124 = ~OLD_REG_1__SCAN_IN; 
assign U125 = ~D_IN_REG_3__SCAN_IN; 
assign U126 = ~OLD_REG_2__SCAN_IN; 
assign U127 = ~D_IN_REG_4__SCAN_IN; 
assign U128 = ~OLD_REG_3__SCAN_IN; 
assign U129 = ~D_IN_REG_5__SCAN_IN; 
assign U130 = ~OLD_REG_4__SCAN_IN; 
assign U131 = ~D_IN_REG_6__SCAN_IN; 
assign U132 = ~OLD_REG_5__SCAN_IN; 
assign U133 = ~D_IN_REG_8__SCAN_IN; 
assign U134 = ~OLD_REG_7__SCAN_IN; 
assign U135 = ~D_IN_REG_7__SCAN_IN; 
assign U136 = ~OLD_REG_6__SCAN_IN; 
assign U137 = ~STATO_REG_1__SCAN_IN; 
assign U139 = ~(STATO_REG_0__SCAN_IN & D_IN_REG_0__SCAN_IN); 
assign U196 = Y_REG_SCAN_IN | D_IN_REG_0__SCAN_IN; 
assign U226 = STATO_REG_0__SCAN_IN | D_IN_REG_0__SCAN_IN; 
assign U92 = ~(U137 & U139); 
assign U141 = ~(U119 & STATO_REG_1__SCAN_IN); 
assign U142 = ~(U137 & STATO_REG_0__SCAN_IN); 
assign U151 = ~U139; 
assign U152 = ~(U120 & STATO_REG_1__SCAN_IN); 
assign U178 = ~(U120 & STATO_REG_0__SCAN_IN); 
assign U201 = ~(U87 & U120); 
assign U207 = ~(U122 & D_IN_REG_1__SCAN_IN); 
assign U208 = ~(U121 & OLD_REG_0__SCAN_IN); 
assign U209 = ~(U124 & D_IN_REG_2__SCAN_IN); 
assign U210 = ~(U123 & OLD_REG_1__SCAN_IN); 
assign U211 = ~(U126 & D_IN_REG_3__SCAN_IN); 
assign U212 = ~(U125 & OLD_REG_2__SCAN_IN); 
assign U213 = ~(U128 & D_IN_REG_4__SCAN_IN); 
assign U214 = ~(U127 & OLD_REG_3__SCAN_IN); 
assign U215 = ~(U130 & D_IN_REG_5__SCAN_IN); 
assign U216 = ~(U129 & OLD_REG_4__SCAN_IN); 
assign U217 = ~(U132 & D_IN_REG_6__SCAN_IN); 
assign U218 = ~(U131 & OLD_REG_5__SCAN_IN); 
assign U219 = ~(U134 & D_IN_REG_8__SCAN_IN); 
assign U220 = ~(U133 & OLD_REG_7__SCAN_IN); 
assign U221 = ~(U136 & D_IN_REG_7__SCAN_IN); 
assign U222 = ~(U135 & OLD_REG_6__SCAN_IN); 
assign U223 = ~(U120 & STATO_REG_0__SCAN_IN); 
assign U225 = ~(U137 & D_IN_REG_0__SCAN_IN); 
assign U90 = U141 & U201; 
assign U143 = U210 & U209 & U208 & U207; 
assign U144 = U214 & U213 & U212 & U211; 
assign U145 = U218 & U217 & U216 & U215; 
assign U146 = U222 & U221 & U220 & U219; 
assign U148 = ~U142; 
assign U149 = ~U141; 
assign U179 = ~(U141 & U178); 
assign U180 = ~(U151 & D_IN_REG_8__SCAN_IN); 
assign U182 = ~(U151 & D_IN_REG_7__SCAN_IN); 
assign U184 = ~(U151 & D_IN_REG_6__SCAN_IN); 
assign U186 = ~(U151 & D_IN_REG_5__SCAN_IN); 
assign U188 = ~(U151 & D_IN_REG_4__SCAN_IN); 
assign U190 = ~(U151 & D_IN_REG_3__SCAN_IN); 
assign U192 = ~(U151 & D_IN_REG_2__SCAN_IN); 
assign U194 = ~(U151 & D_IN_REG_1__SCAN_IN); 
assign U224 = ~(U152 & U119); 
assign U138 = ~(U146 & U145 & U144 & U143); 
assign U181 = ~(U179 & OLD_REG_7__SCAN_IN); 
assign U183 = ~(U179 & OLD_REG_6__SCAN_IN); 
assign U185 = ~(U179 & OLD_REG_5__SCAN_IN); 
assign U187 = ~(U179 & OLD_REG_4__SCAN_IN); 
assign U189 = ~(U179 & OLD_REG_3__SCAN_IN); 
assign U191 = ~(U179 & OLD_REG_2__SCAN_IN); 
assign U193 = ~(U179 & OLD_REG_1__SCAN_IN); 
assign U195 = ~(U179 & OLD_REG_0__SCAN_IN); 
assign U197 = ~(U120 & U149 & D_OUT_REG_0__SCAN_IN); 
assign U198 = ~(U148 & U196); 
assign U202 = ~(U90 & U142); 
assign U205 = ~(U148 & U120); 
assign U103 = ~(U195 & U194); 
assign U104 = ~(U193 & U192); 
assign U105 = ~(U191 & U190); 
assign U106 = ~(U189 & U188); 
assign U107 = ~(U187 & U186); 
assign U108 = ~(U185 & U184); 
assign U109 = ~(U183 & U182); 
assign U110 = ~(U181 & U180); 
assign U147 = ~U138; 
assign U150 = ~(U151 & U138); 
assign U199 = ~(U87 & U138); 
assign U203 = ~(X & U202); 
assign U206 = ~(U90 & U205); 
assign U93 = U206 & D_IN_REG_1__SCAN_IN; 
assign U94 = U206 & D_IN_REG_2__SCAN_IN; 
assign U95 = U206 & D_IN_REG_3__SCAN_IN; 
assign U96 = U206 & D_IN_REG_4__SCAN_IN; 
assign U97 = U206 & D_IN_REG_5__SCAN_IN; 
assign U98 = U206 & D_IN_REG_6__SCAN_IN; 
assign U99 = U206 & D_IN_REG_7__SCAN_IN; 
assign U100 = U206 & D_IN_REG_8__SCAN_IN; 
assign U102 = ~(U197 & U198 & U150); 
assign U140 = ~(U226 & U225 & U150); 
assign U153 = ~(U147 & U87); 
assign U200 = ~(U142 & U199); 
assign U88 = U140 & STATO_REG_0__SCAN_IN; 
assign U89 = U149 & U140; 
assign U91 = ~(U224 & U223 & U153); 
assign U154 = ~U140; 
assign U204 = ~(U200 & D_IN_REG_0__SCAN_IN); 
assign U101 = ~(U204 & U203); 
assign U155 = ~(U88 & D_IN_REG_8__SCAN_IN); 
assign U156 = ~(U154 & D_OUT_REG_7__SCAN_IN); 
assign U157 = ~(U89 & D_OUT_REG_7__SCAN_IN); 
assign U158 = ~(U88 & D_IN_REG_7__SCAN_IN); 
assign U159 = ~(U154 & D_OUT_REG_6__SCAN_IN); 
assign U160 = ~(U89 & D_OUT_REG_6__SCAN_IN); 
assign U161 = ~(U88 & D_IN_REG_6__SCAN_IN); 
assign U162 = ~(U154 & D_OUT_REG_5__SCAN_IN); 
assign U163 = ~(U89 & D_OUT_REG_5__SCAN_IN); 
assign U164 = ~(U88 & D_IN_REG_5__SCAN_IN); 
assign U165 = ~(U154 & D_OUT_REG_4__SCAN_IN); 
assign U166 = ~(U89 & D_OUT_REG_4__SCAN_IN); 
assign U167 = ~(U88 & D_IN_REG_4__SCAN_IN); 
assign U168 = ~(U154 & D_OUT_REG_3__SCAN_IN); 
assign U169 = ~(U89 & D_OUT_REG_3__SCAN_IN); 
assign U170 = ~(U88 & D_IN_REG_3__SCAN_IN); 
assign U171 = ~(U154 & D_OUT_REG_2__SCAN_IN); 
assign U172 = ~(U89 & D_OUT_REG_2__SCAN_IN); 
assign U173 = ~(U88 & D_IN_REG_2__SCAN_IN); 
assign U174 = ~(U154 & D_OUT_REG_1__SCAN_IN); 
assign U175 = ~(U89 & D_OUT_REG_1__SCAN_IN); 
assign U176 = ~(U88 & D_IN_REG_1__SCAN_IN); 
assign U177 = ~(U154 & D_OUT_REG_0__SCAN_IN); 
assign U111 = ~(U176 & U175 & U177); 
assign U112 = ~(U173 & U172 & U174); 
assign U113 = ~(U170 & U169 & U171); 
assign U114 = ~(U167 & U166 & U168); 
assign U115 = ~(U164 & U163 & U165); 
assign U116 = ~(U161 & U160 & U162); 
assign U117 = ~(U158 & U157 & U159); 
assign U118 = ~(U156 & U155); 
endmodule 
