module b07_C( START, STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, PUNTI_RETTA_REG_7__SCAN_IN, PUNTI_RETTA_REG_6__SCAN_IN, PUNTI_RETTA_REG_5__SCAN_IN, PUNTI_RETTA_REG_4__SCAN_IN, PUNTI_RETTA_REG_3__SCAN_IN, PUNTI_RETTA_REG_2__SCAN_IN, PUNTI_RETTA_REG_1__SCAN_IN, PUNTI_RETTA_REG_0__SCAN_IN, CONT_REG_7__SCAN_IN, CONT_REG_6__SCAN_IN, CONT_REG_5__SCAN_IN, CONT_REG_4__SCAN_IN, CONT_REG_3__SCAN_IN, CONT_REG_2__SCAN_IN, CONT_REG_1__SCAN_IN, CONT_REG_0__SCAN_IN, MAR_REG_7__SCAN_IN, MAR_REG_6__SCAN_IN, MAR_REG_5__SCAN_IN, MAR_REG_4__SCAN_IN, MAR_REG_3__SCAN_IN, MAR_REG_2__SCAN_IN, MAR_REG_1__SCAN_IN, MAR_REG_0__SCAN_IN, X_REG_7__SCAN_IN, X_REG_6__SCAN_IN, X_REG_5__SCAN_IN, X_REG_4__SCAN_IN, X_REG_3__SCAN_IN, X_REG_2__SCAN_IN, X_REG_1__SCAN_IN, X_REG_0__SCAN_IN, Y_REG_3__SCAN_IN, Y_REG_1__SCAN_IN, Y_REG_5__SCAN_IN, T_REG_3__SCAN_IN, T_REG_5__SCAN_IN, T_REG_1__SCAN_IN, T_REG_0__SCAN_IN, T_REG_4__SCAN_IN, T_REG_6__SCAN_IN, T_REG_2__SCAN_IN, Y_REG_4__SCAN_IN, Y_REG_0__SCAN_IN, Y_REG_2__SCAN_IN, Y_REG_6__SCAN_IN, STATO_REG_2__SCAN_IN, U324, U325, U326, U327, U328, U329, U330, U331, U332, U333, U334, U335, U336, U337, U338, U339, U340, U341, U342, U343, U344, U345, U346, U347, U348, U349, U350, U351, U352, U353, U354, U355, U356, U357, U358, U388, U389, U390, U391, U394, U395, U396, U397, U398, U399, U400, U401, U402, U403); 
input START, STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, PUNTI_RETTA_REG_7__SCAN_IN, PUNTI_RETTA_REG_6__SCAN_IN, PUNTI_RETTA_REG_5__SCAN_IN, PUNTI_RETTA_REG_4__SCAN_IN, PUNTI_RETTA_REG_3__SCAN_IN, PUNTI_RETTA_REG_2__SCAN_IN, PUNTI_RETTA_REG_1__SCAN_IN, PUNTI_RETTA_REG_0__SCAN_IN, CONT_REG_7__SCAN_IN, CONT_REG_6__SCAN_IN, CONT_REG_5__SCAN_IN, CONT_REG_4__SCAN_IN, CONT_REG_3__SCAN_IN, CONT_REG_2__SCAN_IN, CONT_REG_1__SCAN_IN, CONT_REG_0__SCAN_IN, MAR_REG_7__SCAN_IN, MAR_REG_6__SCAN_IN, MAR_REG_5__SCAN_IN, MAR_REG_4__SCAN_IN, MAR_REG_3__SCAN_IN, MAR_REG_2__SCAN_IN, MAR_REG_1__SCAN_IN, MAR_REG_0__SCAN_IN, X_REG_7__SCAN_IN, X_REG_6__SCAN_IN, X_REG_5__SCAN_IN, X_REG_4__SCAN_IN, X_REG_3__SCAN_IN, X_REG_2__SCAN_IN, X_REG_1__SCAN_IN, X_REG_0__SCAN_IN, Y_REG_3__SCAN_IN, Y_REG_1__SCAN_IN, Y_REG_5__SCAN_IN, T_REG_3__SCAN_IN, T_REG_5__SCAN_IN, T_REG_1__SCAN_IN, T_REG_0__SCAN_IN, T_REG_4__SCAN_IN, T_REG_6__SCAN_IN, T_REG_2__SCAN_IN, Y_REG_4__SCAN_IN, Y_REG_0__SCAN_IN, Y_REG_2__SCAN_IN, Y_REG_6__SCAN_IN, STATO_REG_2__SCAN_IN; 
output U324, U325, U326, U327, U328, U329, U330, U331, U332, U333, U334, U335, U336, U337, U338, U339, U340, U341, U342, U343, U344, U345, U346, U347, U348, U349, U350, U351, U352, U353, U354, U355, U356, U357, U358, U388, U389, U390, U391, U394, U395, U396, U397, U398, U399, U400, U401, U402, U403; 
wire U300, U301, U302, U303, U304, U305, U306, U307, U308, U309, U310, U311, U312, U313, U314, U315, U316, U317, U318, U319, U320, U321, U322, U323, U359, U360, U361, U362, U363, U364, U365, U366, U367, U368, U369, U370, U371, U372, U373, U374, U375, U376, U377, U378, U379, U380, U381, U382, U383, U384, U385, U386, U387, U392, U393, U404, U405, U406, U407, U408, U409, U410, U411, U412, U413, U414, U415, U416, U417, U418, U419, U420, U421, U422, U423, U424, U425, U426, U427, U428, U429, U430, U431, U432, U433, U434, U435, U436, U437, U438, U439, U440, U441, U442, U443, U444, U445, U446, U447, U448, U449, U450, U451, U452, U453, U454, U455, U456, U457, U458, U459, U460, U461, U462, U463, U464, U465, U466, U467, U468, U469, U470, U471, U472, U473, U474, U475, U476, U477, U478, U479, U480, U481, U482, U483, U484, U485, U486, U487, U488, U489, U490, U491, U492, U493, U494, U495, U496, U497, U498, U499, U500, U501, U502, U503, U504, U505, U506, U507, U508, U509, U510, U511, U512, U513, U514, U515, U516, U517, U518, U519, U520, U521, U522, U523, U524, U525, U526, U527, U528, U529, U530, U531, U532, U533, U534, U535, U536, U537, U538, U539, U540, U541, U542, U543, U544, U545, U546, U547, U548, U549, U550, U551, U552, U553, U554, U555, U556, U557, U558, U559, U560, U561, U562, U563, U564, U565, U566, U567, U568, U569, U570, U571, U572, U573, U574, U575, U576, U577, U578, U579, U580, U581, U582, U583, U584, U585, U586, U587, R182_U4, R182_U5, R182_U6, R182_U7, R182_U8, R182_U9, R182_U10, R182_U11, R182_U12, R182_U13, R182_U14, R182_U15, R182_U16, R182_U17, R182_U18, R182_U19, R182_U20, R182_U21, R182_U22, R182_U23, R182_U24, R182_U25, R182_U26, R182_U27, R182_U28, R182_U29, R182_U30, R182_U31, R182_U32, R182_U33, R182_U34, R182_U35, R182_U36, R182_U37, R182_U38, R182_U39, R182_U40, R182_U41, R182_U42, R182_U43, R182_U44, R182_U45, R182_U46, R182_U47, R182_U48, R182_U49, R182_U50, R182_U51, R182_U52, R182_U53, R182_U54, R182_U55, R182_U56, R182_U57, R182_U58, R182_U59, R182_U60, R182_U61, R182_U62, R182_U63, R182_U64, R182_U65, R182_U66, R182_U67, R182_U68, R182_U69, R182_U70, R182_U71, R182_U72, R182_U73, R182_U74, R182_U75, R182_U76, R182_U77, R182_U78, R182_U79, R182_U80, R182_U81, R182_U82, R182_U83, R182_U84, R182_U85, R182_U86, R182_U87, R182_U88, R182_U89, R182_U90, R182_U91, R182_U92, R182_U93, R182_U94, R182_U95, R182_U96, R182_U97, R182_U98; 
assign U307 = START & STATO_REG_0__SCAN_IN; 
assign U359 = ~MAR_REG_1__SCAN_IN; 
assign U360 = ~MAR_REG_0__SCAN_IN; 
assign U361 = ~(MAR_REG_1__SCAN_IN & MAR_REG_0__SCAN_IN); 
assign U362 = ~MAR_REG_2__SCAN_IN; 
assign U364 = ~MAR_REG_3__SCAN_IN; 
assign U366 = ~START; 
assign U367 = ~STATO_REG_1__SCAN_IN; 
assign U368 = ~STATO_REG_2__SCAN_IN; 
assign U369 = ~STATO_REG_0__SCAN_IN; 
assign U370 = ~(STATO_REG_2__SCAN_IN & STATO_REG_1__SCAN_IN); 
assign U371 = STATO_REG_2__SCAN_IN | STATO_REG_1__SCAN_IN; 
assign U377 = ~MAR_REG_7__SCAN_IN; 
assign U378 = ~MAR_REG_6__SCAN_IN; 
assign U379 = ~MAR_REG_5__SCAN_IN; 
assign U380 = ~MAR_REG_4__SCAN_IN; 
assign U381 = ~X_REG_3__SCAN_IN; 
assign U382 = ~X_REG_2__SCAN_IN; 
assign U384 = ~X_REG_0__SCAN_IN; 
assign U385 = STATO_REG_1__SCAN_IN | STATO_REG_0__SCAN_IN; 
assign U387 = ~(STATO_REG_2__SCAN_IN & STATO_REG_0__SCAN_IN); 
assign U405 = ~(X_REG_7__SCAN_IN | X_REG_6__SCAN_IN | X_REG_5__SCAN_IN | X_REG_4__SCAN_IN); 
assign U406 = STATO_REG_2__SCAN_IN | STATO_REG_0__SCAN_IN; 
assign U407 = ~(STATO_REG_1__SCAN_IN & STATO_REG_0__SCAN_IN); 
assign U505 = MAR_REG_3__SCAN_IN | MAR_REG_2__SCAN_IN | MAR_REG_1__SCAN_IN; 
assign U308 = U362 & MAR_REG_3__SCAN_IN; 
assign U373 = ~(U384 & U382 & U381 & U405 & X_REG_1__SCAN_IN); 
assign U404 = U378 & U377 & U379 & U380 & MAR_REG_3__SCAN_IN; 
assign U408 = ~U385; 
assign U409 = ~U387; 
assign U415 = ~U370; 
assign U416 = ~U407; 
assign U417 = ~U361; 
assign U423 = ~U406; 
assign U427 = ~U371; 
assign U476 = ~(U307 & U368); 
assign U480 = ~(U371 & U361); 
assign U482 = ~(U371 & U360); 
assign U499 = ~(U359 & MAR_REG_0__SCAN_IN); 
assign U517 = ~(U368 & X_REG_6__SCAN_IN); 
assign U520 = ~(U368 & X_REG_5__SCAN_IN); 
assign U523 = ~(U368 & X_REG_4__SCAN_IN); 
assign U526 = ~(U368 & X_REG_3__SCAN_IN); 
assign U529 = ~(U368 & X_REG_2__SCAN_IN); 
assign U532 = ~(U368 & X_REG_1__SCAN_IN); 
assign U535 = ~(U368 & X_REG_0__SCAN_IN); 
assign U537 = ~(U385 & U387 & STATO_REG_2__SCAN_IN); 
assign U552 = ~(U307 & U367); 
assign U562 = ~(U367 & STATO_REG_2__SCAN_IN); 
assign U565 = ~(U364 & U362 & U359 & MAR_REG_0__SCAN_IN); 
assign U570 = ~(U407 & T_REG_3__SCAN_IN); 
assign U572 = ~(U407 & T_REG_5__SCAN_IN); 
assign U574 = ~(U407 & T_REG_1__SCAN_IN); 
assign U576 = ~(U407 & T_REG_0__SCAN_IN); 
assign U578 = ~(U407 & T_REG_4__SCAN_IN); 
assign U580 = ~(U407 & T_REG_6__SCAN_IN); 
assign U582 = ~(U407 & T_REG_2__SCAN_IN); 
assign U363 = ~(U417 & MAR_REG_2__SCAN_IN); 
assign U386 = ~(U408 & STATO_REG_2__SCAN_IN); 
assign U430 = ~(U427 & STATO_REG_0__SCAN_IN); 
assign U432 = ~U373; 
assign U457 = ~(U427 & U307); 
assign U494 = ~(U308 & U417); 
assign U515 = ~(U409 & Y_REG_6__SCAN_IN); 
assign U516 = ~(U408 & T_REG_6__SCAN_IN); 
assign U518 = ~(U409 & Y_REG_5__SCAN_IN); 
assign U519 = ~(U408 & T_REG_5__SCAN_IN); 
assign U521 = ~(U409 & Y_REG_4__SCAN_IN); 
assign U522 = ~(U408 & T_REG_4__SCAN_IN); 
assign U524 = ~(U409 & Y_REG_3__SCAN_IN); 
assign U525 = ~(U408 & T_REG_3__SCAN_IN); 
assign U527 = ~(U409 & Y_REG_2__SCAN_IN); 
assign U528 = ~(U408 & T_REG_2__SCAN_IN); 
assign U530 = ~(U409 & Y_REG_1__SCAN_IN); 
assign U531 = ~(U408 & T_REG_1__SCAN_IN); 
assign U533 = ~(U409 & Y_REG_0__SCAN_IN); 
assign U534 = ~(U408 & T_REG_0__SCAN_IN); 
assign U539 = ~(U537 & X_REG_6__SCAN_IN); 
assign U541 = ~(U537 & X_REG_5__SCAN_IN); 
assign U543 = ~(U537 & X_REG_4__SCAN_IN); 
assign U545 = ~(U537 & X_REG_3__SCAN_IN); 
assign U547 = ~(U537 & X_REG_2__SCAN_IN); 
assign U549 = ~(U537 & X_REG_1__SCAN_IN); 
assign U551 = ~(U537 & X_REG_0__SCAN_IN); 
assign U563 = ~(U423 & STATO_REG_1__SCAN_IN); 
assign U566 = ~(U308 & U360 & MAR_REG_1__SCAN_IN); 
assign U317 = ~(U516 & U517 & U515); 
assign U318 = ~(U519 & U520 & U518); 
assign U319 = ~(U522 & U523 & U521); 
assign U320 = ~(U525 & U526 & U524); 
assign U321 = ~(U528 & U529 & U527); 
assign U322 = ~(U531 & U532 & U530); 
assign U323 = ~(U535 & U534 & U533 & U370); 
assign U392 = ~(U566 & U565); 
assign U393 = ~(U563 & U562); 
assign U418 = ~U363; 
assign U478 = ~(U371 & U363); 
assign U510 = ~U386; 
assign U511 = ~(U386 & Y_REG_3__SCAN_IN); 
assign U512 = ~(U386 & Y_REG_5__SCAN_IN); 
assign U513 = ~(U386 & Y_REG_4__SCAN_IN); 
assign U514 = ~(U386 & Y_REG_6__SCAN_IN); 
assign U569 = ~(U386 & Y_REG_1__SCAN_IN); 
assign U585 = ~(U386 & Y_REG_0__SCAN_IN); 
assign U587 = ~(U386 & Y_REG_2__SCAN_IN); 
assign U304 = U393 & U406; 
assign U305 = U393 & U368; 
assign U365 = ~(U404 & U418); 
assign U414 = ~(U510 & U392); 
assign U500 = ~(U418 & MAR_REG_3__SCAN_IN); 
assign U564 = ~U393; 
assign U567 = ~U392; 
assign R182_U5 = ~U323; 
assign R182_U8 = ~U322; 
assign R182_U10 = ~U321; 
assign R182_U12 = ~U320; 
assign R182_U14 = ~U319; 
assign R182_U16 = ~U318; 
assign R182_U18 = ~U317; 
assign U327 = ~(U414 & U514); 
assign U328 = ~(U414 & U513); 
assign U329 = ~(U414 & U512); 
assign U330 = ~(U414 & U511); 
assign U374 = ~(U415 & U365); 
assign U383 = ~(U567 & U494); 
assign U413 = ~(U305 & U392); 
assign U419 = ~U365; 
assign U485 = ~(U564 & X_REG_7__SCAN_IN); 
assign U487 = ~(U564 & X_REG_6__SCAN_IN); 
assign U489 = ~(U564 & X_REG_5__SCAN_IN); 
assign U491 = ~(U564 & X_REG_4__SCAN_IN); 
assign U493 = ~(U564 & X_REG_3__SCAN_IN); 
assign U498 = ~(U564 & X_REG_2__SCAN_IN); 
assign U501 = ~(U567 & U499 & U500); 
assign U504 = ~(U564 & X_REG_1__SCAN_IN); 
assign U509 = ~(U564 & X_REG_0__SCAN_IN); 
assign U376 = ~(U407 & U476 & U374); 
assign U410 = ~U374; 
assign U411 = ~(U415 & U419); 
assign U420 = ~(START & U419); 
assign U424 = ~(U419 & U366); 
assign U495 = ~U383; 
assign U496 = ~(U305 & U383); 
assign U502 = ~(U305 & U501); 
assign U568 = ~(U510 & U501); 
assign U586 = ~(U510 & U383); 
assign U306 = U376 & U371; 
assign U394 = ~(U569 & U568); 
assign U403 = ~(U587 & U586); 
assign U421 = ~(U420 & STATO_REG_1__SCAN_IN); 
assign U425 = ~(U424 & U369); 
assign U428 = ~(U411 & U371); 
assign U431 = ~(U411 & U430); 
assign U458 = ~(U410 & U432); 
assign U477 = ~U376; 
assign U479 = ~(U376 & U478); 
assign U481 = ~(U376 & U480); 
assign U483 = ~(U376 & U482); 
assign U506 = ~(U495 & U505); 
assign U536 = ~(U374 & U411); 
assign U309 = U536 & CONT_REG_7__SCAN_IN; 
assign U339 = U477 & MAR_REG_4__SCAN_IN; 
assign U340 = U477 & MAR_REG_5__SCAN_IN; 
assign U341 = U477 & MAR_REG_6__SCAN_IN; 
assign U342 = U477 & MAR_REG_7__SCAN_IN; 
assign U372 = ~(U431 & U366); 
assign U375 = ~(U458 & U457); 
assign U422 = ~(U421 & STATO_REG_2__SCAN_IN); 
assign U426 = ~(U406 & U425); 
assign U429 = ~(U428 & U366); 
assign U507 = ~(U305 & U506); 
assign U538 = ~(U536 & CONT_REG_6__SCAN_IN); 
assign U540 = ~(U536 & CONT_REG_5__SCAN_IN); 
assign U542 = ~(U536 & CONT_REG_4__SCAN_IN); 
assign U544 = ~(U536 & CONT_REG_3__SCAN_IN); 
assign U546 = ~(U536 & CONT_REG_2__SCAN_IN); 
assign U548 = ~(U536 & CONT_REG_1__SCAN_IN); 
assign U550 = ~(U536 & CONT_REG_0__SCAN_IN); 
assign U554 = ~(U479 & MAR_REG_3__SCAN_IN); 
assign U555 = ~(U306 & U418 & U364); 
assign U556 = ~(U481 & MAR_REG_2__SCAN_IN); 
assign U557 = ~(U306 & U417 & U362); 
assign U558 = ~(U483 & MAR_REG_1__SCAN_IN); 
assign U559 = ~(U306 & U359 & MAR_REG_0__SCAN_IN); 
assign U560 = ~(U306 & U360); 
assign U561 = ~(U477 & MAR_REG_0__SCAN_IN); 
assign U584 = ~(U510 & U506); 
assign U301 = U375 & STATO_REG_2__SCAN_IN; 
assign U310 = ~(U539 & U538); 
assign U311 = ~(U541 & U540); 
assign U312 = ~(U543 & U542); 
assign U313 = ~(U545 & U544); 
assign U314 = ~(U547 & U546); 
assign U315 = ~(U549 & U548); 
assign U316 = ~(U551 & U550); 
assign U324 = ~(U407 & U422); 
assign U326 = ~(U406 & U385 & U429); 
assign U388 = ~(U555 & U554); 
assign U389 = ~(U557 & U556); 
assign U390 = ~(U559 & U558); 
assign U391 = ~(U561 & U560); 
assign U402 = ~(U585 & U584); 
assign U412 = ~U372; 
assign U435 = ~(U372 & PUNTI_RETTA_REG_7__SCAN_IN); 
assign U438 = ~(U372 & PUNTI_RETTA_REG_6__SCAN_IN); 
assign U441 = ~(U372 & PUNTI_RETTA_REG_5__SCAN_IN); 
assign U444 = ~(U372 & PUNTI_RETTA_REG_4__SCAN_IN); 
assign U447 = ~(U372 & PUNTI_RETTA_REG_3__SCAN_IN); 
assign U450 = ~(U372 & PUNTI_RETTA_REG_2__SCAN_IN); 
assign U453 = ~(U372 & PUNTI_RETTA_REG_1__SCAN_IN); 
assign U456 = ~(U372 & PUNTI_RETTA_REG_0__SCAN_IN); 
assign U459 = ~U375; 
assign U553 = ~(U426 & STATO_REG_1__SCAN_IN); 
assign R182_U28 = ~U309; 
assign U300 = U412 & STATO_REG_2__SCAN_IN; 
assign U325 = ~(U553 & U552 & U387); 
assign U461 = ~(U459 & CONT_REG_7__SCAN_IN); 
assign U463 = ~(U459 & CONT_REG_6__SCAN_IN); 
assign U465 = ~(U459 & CONT_REG_5__SCAN_IN); 
assign U467 = ~(U459 & CONT_REG_4__SCAN_IN); 
assign U469 = ~(U459 & CONT_REG_3__SCAN_IN); 
assign U471 = ~(U459 & CONT_REG_2__SCAN_IN); 
assign U473 = ~(U459 & CONT_REG_1__SCAN_IN); 
assign U475 = ~(U459 & CONT_REG_0__SCAN_IN); 
assign R182_U4 = ~U316; 
assign R182_U6 = ~(U323 & U316); 
assign R182_U7 = ~U315; 
assign R182_U9 = ~U314; 
assign R182_U11 = ~U313; 
assign R182_U13 = ~U312; 
assign R182_U15 = ~U311; 
assign R182_U19 = ~U310; 
assign R182_U41 = U315 | U322; 
assign R182_U43 = ~(U322 & U315); 
assign R182_U45 = U314 | U321; 
assign R182_U47 = ~(U321 & U314); 
assign R182_U49 = U313 | U320; 
assign R182_U51 = ~(U320 & U313); 
assign R182_U53 = U312 | U319; 
assign R182_U55 = ~(U319 & U312); 
assign R182_U57 = U311 | U318; 
assign R182_U59 = ~(U318 & U311); 
assign R182_U68 = ~(U310 & R182_U18); 
assign R182_U73 = ~(U311 & R182_U16); 
assign R182_U78 = ~(U312 & R182_U14); 
assign R182_U83 = ~(U313 & R182_U12); 
assign R182_U88 = ~(U314 & R182_U10); 
assign R182_U92 = ~(U315 & R182_U8); 
assign R182_U98 = ~(U316 & R182_U5); 
assign U302 = U300 & U373; 
assign U303 = U300 & U432; 
assign R182_U40 = ~R182_U6; 
assign R182_U67 = ~(U317 & R182_U19); 
assign R182_U72 = ~(U318 & R182_U15); 
assign R182_U77 = ~(U319 & R182_U13); 
assign R182_U82 = ~(U320 & R182_U11); 
assign R182_U87 = ~(U321 & R182_U9); 
assign R182_U93 = ~(U322 & R182_U7); 
assign R182_U97 = ~(U323 & R182_U4); 
assign U434 = ~(U302 & CONT_REG_7__SCAN_IN); 
assign U437 = ~(U302 & CONT_REG_6__SCAN_IN); 
assign U440 = ~(U302 & CONT_REG_5__SCAN_IN); 
assign U443 = ~(U302 & CONT_REG_4__SCAN_IN); 
assign U446 = ~(U302 & CONT_REG_3__SCAN_IN); 
assign U449 = ~(U302 & CONT_REG_2__SCAN_IN); 
assign U452 = ~(U302 & CONT_REG_1__SCAN_IN); 
assign U455 = ~(U302 & CONT_REG_0__SCAN_IN); 
assign R182_U21 = ~(R182_U98 & R182_U97); 
assign R182_U22 = ~(R182_U68 & R182_U67); 
assign R182_U23 = ~(R182_U73 & R182_U72); 
assign R182_U24 = ~(R182_U78 & R182_U77); 
assign R182_U25 = ~(R182_U83 & R182_U82); 
assign R182_U26 = ~(R182_U88 & R182_U87); 
assign R182_U27 = ~(R182_U93 & R182_U92); 
assign R182_U42 = ~(R182_U40 & R182_U41); 
assign U454 = ~(R182_U21 & U303); 
assign U474 = ~(U301 & R182_U21); 
assign U508 = ~(U304 & R182_U21); 
assign U577 = ~(U416 & R182_U21); 
assign R182_U38 = ~(R182_U43 & R182_U42); 
assign R182_U69 = ~R182_U22; 
assign R182_U74 = ~R182_U23; 
assign R182_U79 = ~R182_U24; 
assign R182_U84 = ~R182_U25; 
assign R182_U89 = ~R182_U26; 
assign R182_U94 = ~R182_U27; 
assign R182_U96 = ~(R182_U27 & R182_U6); 
assign U331 = ~(U509 & U507 & U508); 
assign U343 = ~(U475 & U474); 
assign U351 = ~(U455 & U454 & U456); 
assign U398 = ~(U577 & U576); 
assign R182_U44 = ~R182_U38; 
assign R182_U46 = ~(R182_U45 & R182_U38); 
assign R182_U91 = ~(R182_U26 & R182_U38); 
assign R182_U95 = ~(R182_U94 & R182_U40); 
assign R182_U20 = ~(R182_U96 & R182_U95); 
assign R182_U36 = ~(R182_U47 & R182_U46); 
assign R182_U90 = ~(R182_U44 & R182_U89); 
assign U451 = ~(R182_U20 & U303); 
assign U472 = ~(U301 & R182_U20); 
assign U503 = ~(U304 & R182_U20); 
assign U575 = ~(U416 & R182_U20); 
assign R182_U39 = R182_U91 & R182_U90; 
assign R182_U48 = ~R182_U36; 
assign R182_U50 = ~(R182_U49 & R182_U36); 
assign R182_U86 = ~(R182_U25 & R182_U36); 
assign U332 = ~(U504 & U502 & U503); 
assign U344 = ~(U473 & U472); 
assign U352 = ~(U452 & U453 & U451); 
assign U397 = ~(U575 & U574); 
assign U448 = ~(R182_U39 & U303); 
assign U470 = ~(U301 & R182_U39); 
assign U497 = ~(U304 & R182_U39); 
assign U583 = ~(U416 & R182_U39); 
assign R182_U34 = ~(R182_U51 & R182_U50); 
assign R182_U85 = ~(R182_U48 & R182_U84); 
assign U333 = ~(U498 & U496 & U497); 
assign U345 = ~(U471 & U470); 
assign U353 = ~(U449 & U450 & U448); 
assign U401 = ~(U583 & U582); 
assign R182_U37 = R182_U86 & R182_U85; 
assign R182_U52 = ~R182_U34; 
assign R182_U54 = ~(R182_U53 & R182_U34); 
assign R182_U81 = ~(R182_U24 & R182_U34); 
assign U445 = ~(R182_U37 & U303); 
assign U468 = ~(U301 & R182_U37); 
assign U492 = ~(U304 & R182_U37); 
assign U571 = ~(U416 & R182_U37); 
assign R182_U32 = ~(R182_U55 & R182_U54); 
assign R182_U80 = ~(R182_U52 & R182_U79); 
assign U334 = ~(U493 & U413 & U492); 
assign U346 = ~(U469 & U468); 
assign U354 = ~(U446 & U447 & U445); 
assign U395 = ~(U571 & U570); 
assign R182_U35 = R182_U81 & R182_U80; 
assign R182_U56 = ~R182_U32; 
assign R182_U58 = ~(R182_U57 & R182_U32); 
assign R182_U76 = ~(R182_U23 & R182_U32); 
assign U442 = ~(R182_U35 & U303); 
assign U466 = ~(U301 & R182_U35); 
assign U490 = ~(U304 & R182_U35); 
assign U579 = ~(U416 & R182_U35); 
assign R182_U17 = ~(R182_U59 & R182_U58); 
assign R182_U75 = ~(R182_U56 & R182_U74); 
assign U335 = ~(U491 & U413 & U490); 
assign U347 = ~(U467 & U466); 
assign U355 = ~(U443 & U444 & U442); 
assign U399 = ~(U579 & U578); 
assign R182_U33 = R182_U76 & R182_U75; 
assign R182_U60 = ~R182_U17; 
assign R182_U63 = ~(U310 & R182_U17); 
assign R182_U71 = ~(R182_U22 & R182_U17); 
assign U439 = ~(R182_U33 & U303); 
assign U464 = ~(U301 & R182_U33); 
assign U488 = ~(U304 & R182_U33); 
assign U573 = ~(U416 & R182_U33); 
assign R182_U61 = ~(R182_U60 & R182_U19); 
assign R182_U70 = ~(R182_U69 & R182_U60); 
assign U336 = ~(U489 & U413 & U488); 
assign U348 = ~(U465 & U464); 
assign U356 = ~(U440 & U441 & U439); 
assign U396 = ~(U573 & U572); 
assign R182_U31 = R182_U71 & R182_U70; 
assign R182_U62 = ~(U317 & R182_U61); 
assign U436 = ~(R182_U31 & U303); 
assign U462 = ~(U301 & R182_U31); 
assign U486 = ~(U304 & R182_U31); 
assign U581 = ~(U416 & R182_U31); 
assign R182_U29 = ~(R182_U63 & R182_U62); 
assign U337 = ~(U487 & U413 & U486); 
assign U349 = ~(U463 & U462); 
assign U357 = ~(U437 & U438 & U436); 
assign U400 = ~(U581 & U580); 
assign R182_U64 = ~R182_U29; 
assign R182_U65 = ~(U309 & R182_U29); 
assign R182_U66 = ~(R182_U64 & R182_U28); 
assign R182_U30 = R182_U66 & R182_U65; 
assign U433 = ~(R182_U30 & U303); 
assign U460 = ~(U301 & R182_U30); 
assign U484 = ~(U304 & R182_U30); 
assign U338 = ~(U485 & U413 & U484); 
assign U350 = ~(U461 & U460); 
assign U358 = ~(U434 & U435 & U433); 
endmodule 
