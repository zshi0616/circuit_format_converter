module b15_C( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U2788, U2789, U2790, U2791, U2792, U2793, U2794, U2795, U2796, U2797, U2798, U2799, U2800, U2801, U2802, U2803, U2804, U2805, U2806, U2807, U2808, U2809, U2810, U2811, U2812, U2813, U2814, U2815, U2816, U2817, U2818, U2819, U2820, U2821, U2822, U2823, U2824, U2825, U2826, U2827, U2828, U2829, U2830, U2831, U2832, U2833, U2834, U2835, U2836, U2837, U2838, U2839, U2840, U2841, U2842, U2843, U2844, U2845, U2846, U2847, U2848, U2849, U2850, U2851, U2852, U2853, U2854, U2855, U2856, U2857, U2858, U2859, U2860, U2861, U2862, U2863, U2864, U2865, U2866, U2867, U2868, U2869, U2870, U2871, U2872, U2873, U2874, U2875, U2876, U2877, U2878, U2879, U2880, U2881, U2882, U2883, U2884, U2885, U2886, U2887, U2888, U2889, U2890, U2891, U2892, U2893, U2894, U2895, U2896, U2897, U2898, U2899, U2900, U2901, U2902, U2903, U2904, U2905, U2906, U2907, U2908, U2909, U2910, U2911, U2912, U2913, U2914, U2915, U2916, U2917, U2918, U2919, U2920, U2921, U2922, U2923, U2924, U2925, U2926, U2927, U2928, U2929, U2930, U2931, U2932, U2933, U2934, U2935, U2936, U2937, U2938, U2939, U2940, U2941, U2942, U2943, U2944, U2945, U2946, U2947, U2948, U2949, U2950, U2951, U2952, U2953, U2954, U2955, U2956, U2957, U2958, U2959, U2960, U2961, U2962, U2963, U2964, U2965, U2966, U2967, U2968, U2969, U2970, U2971, U2972, U2973, U2974, U2975, U2976, U2977, U2978, U2979, U2980, U2981, U2982, U2983, U2984, U2985, U2986, U2987, U2988, U2989, U2990, U2991, U2992, U2993, U2994, U2995, U2996, U2997, U2998, U2999, U3000, U3001, U3002, U3003, U3004, U3005, U3006, U3007, U3008, U3009, U3010, U3011, U3012, U3013, U3014, U3015, U3016, U3017, U3018, U3019, U3020, U3021, U3022, U3023, U3024, U3025, U3026, U3027, U3028, U3029, U3030, U3031, U3032, U3033, U3034, U3035, U3036, U3037, U3038, U3039, U3040, U3041, U3042, U3043, U3044, U3045, U3046, U3047, U3048, U3049, U3050, U3051, U3052, U3053, U3054, U3055, U3056, U3057, U3058, U3059, U3060, U3061, U3062, U3063, U3064, U3065, U3066, U3067, U3068, U3069, U3070, U3071, U3072, U3073, U3074, U3075, U3076, U3077, U3078, U3079, U3080, U3081, U3082, U3083, U3084, U3085, U3086, U3087, U3088, U3089, U3090, U3091, U3092, U3093, U3094, U3095, U3096, U3097, U3098, U3099, U3100, U3101, U3102, U3103, U3104, U3105, U3106, U3107, U3108, U3109, U3110, U3111, U3112, U3113, U3114, U3115, U3116, U3117, U3118, U3119, U3120, U3121, U3122, U3123, U3124, U3125, U3126, U3127, U3128, U3129, U3130, U3131, U3132, U3133, U3134, U3135, U3136, U3137, U3138, U3139, U3140, U3141, U3142, U3143, U3144, U3145, U3146, U3147, U3148, U3149, U3150, U3151, U3152, U3153, U3154, U3155, U3156, U3157, U3158, U3159, U3160, U3161, U3162, U3163, U3164, U3165, U3166, U3167, U3168, U3169, U3170, U3171, U3172, U3173, U3174, U3175, U3176, U3177, U3178, U3179, U3180, U3181, U3182, U3183, U3184, U3185, U3186, U3187, U3188, U3189, U3190, U3191, U3192, U3193, U3194, U3195, U3196, U3197, U3198, U3199, U3200, U3201, U3202, U3203, U3204, U3205, U3206, U3207, U3208, U3209, U3210, U3211, U3212, U3213, U3445, U3446, U3447, U3448, U3451, U3452, U3453, U3455, U3456, U3459, U3460, U3461, U3462, U3463, U3464, U3465, U3468, U3469, U3470, U3471, U3472, U3473, U3474); 
input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN; 
output U2788, U2789, U2790, U2791, U2792, U2793, U2794, U2795, U2796, U2797, U2798, U2799, U2800, U2801, U2802, U2803, U2804, U2805, U2806, U2807, U2808, U2809, U2810, U2811, U2812, U2813, U2814, U2815, U2816, U2817, U2818, U2819, U2820, U2821, U2822, U2823, U2824, U2825, U2826, U2827, U2828, U2829, U2830, U2831, U2832, U2833, U2834, U2835, U2836, U2837, U2838, U2839, U2840, U2841, U2842, U2843, U2844, U2845, U2846, U2847, U2848, U2849, U2850, U2851, U2852, U2853, U2854, U2855, U2856, U2857, U2858, U2859, U2860, U2861, U2862, U2863, U2864, U2865, U2866, U2867, U2868, U2869, U2870, U2871, U2872, U2873, U2874, U2875, U2876, U2877, U2878, U2879, U2880, U2881, U2882, U2883, U2884, U2885, U2886, U2887, U2888, U2889, U2890, U2891, U2892, U2893, U2894, U2895, U2896, U2897, U2898, U2899, U2900, U2901, U2902, U2903, U2904, U2905, U2906, U2907, U2908, U2909, U2910, U2911, U2912, U2913, U2914, U2915, U2916, U2917, U2918, U2919, U2920, U2921, U2922, U2923, U2924, U2925, U2926, U2927, U2928, U2929, U2930, U2931, U2932, U2933, U2934, U2935, U2936, U2937, U2938, U2939, U2940, U2941, U2942, U2943, U2944, U2945, U2946, U2947, U2948, U2949, U2950, U2951, U2952, U2953, U2954, U2955, U2956, U2957, U2958, U2959, U2960, U2961, U2962, U2963, U2964, U2965, U2966, U2967, U2968, U2969, U2970, U2971, U2972, U2973, U2974, U2975, U2976, U2977, U2978, U2979, U2980, U2981, U2982, U2983, U2984, U2985, U2986, U2987, U2988, U2989, U2990, U2991, U2992, U2993, U2994, U2995, U2996, U2997, U2998, U2999, U3000, U3001, U3002, U3003, U3004, U3005, U3006, U3007, U3008, U3009, U3010, U3011, U3012, U3013, U3014, U3015, U3016, U3017, U3018, U3019, U3020, U3021, U3022, U3023, U3024, U3025, U3026, U3027, U3028, U3029, U3030, U3031, U3032, U3033, U3034, U3035, U3036, U3037, U3038, U3039, U3040, U3041, U3042, U3043, U3044, U3045, U3046, U3047, U3048, U3049, U3050, U3051, U3052, U3053, U3054, U3055, U3056, U3057, U3058, U3059, U3060, U3061, U3062, U3063, U3064, U3065, U3066, U3067, U3068, U3069, U3070, U3071, U3072, U3073, U3074, U3075, U3076, U3077, U3078, U3079, U3080, U3081, U3082, U3083, U3084, U3085, U3086, U3087, U3088, U3089, U3090, U3091, U3092, U3093, U3094, U3095, U3096, U3097, U3098, U3099, U3100, U3101, U3102, U3103, U3104, U3105, U3106, U3107, U3108, U3109, U3110, U3111, U3112, U3113, U3114, U3115, U3116, U3117, U3118, U3119, U3120, U3121, U3122, U3123, U3124, U3125, U3126, U3127, U3128, U3129, U3130, U3131, U3132, U3133, U3134, U3135, U3136, U3137, U3138, U3139, U3140, U3141, U3142, U3143, U3144, U3145, U3146, U3147, U3148, U3149, U3150, U3151, U3152, U3153, U3154, U3155, U3156, U3157, U3158, U3159, U3160, U3161, U3162, U3163, U3164, U3165, U3166, U3167, U3168, U3169, U3170, U3171, U3172, U3173, U3174, U3175, U3176, U3177, U3178, U3179, U3180, U3181, U3182, U3183, U3184, U3185, U3186, U3187, U3188, U3189, U3190, U3191, U3192, U3193, U3194, U3195, U3196, U3197, U3198, U3199, U3200, U3201, U3202, U3203, U3204, U3205, U3206, U3207, U3208, U3209, U3210, U3211, U3212, U3213, U3445, U3446, U3447, U3448, U3451, U3452, U3453, U3455, U3456, U3459, U3460, U3461, U3462, U3463, U3464, U3465, U3468, U3469, U3470, U3471, U3472, U3473, U3474; 
wire U2352, U2353, U2354, U2355, U2356, U2357, U2358, U2359, U2360, U2361, U2362, U2363, U2364, U2365, U2366, U2367, U2368, U2369, U2370, U2371, U2372, U2373, U2374, U2375, U2376, U2377, U2378, U2379, U2380, U2381, U2382, U2383, U2384, U2385, U2386, U2387, U2388, U2389, U2390, U2391, U2392, U2393, U2394, U2395, U2396, U2397, U2398, U2399, U2400, U2401, U2402, U2403, U2404, U2405, U2406, U2407, U2408, U2409, U2410, U2411, U2412, U2413, U2414, U2415, U2416, U2417, U2418, U2419, U2420, U2421, U2422, U2423, U2424, U2425, U2426, U2427, U2428, U2429, U2430, U2431, U2432, U2433, U2434, U2435, U2436, U2437, U2438, U2439, U2440, U2441, U2442, U2443, U2444, U2445, U2446, U2447, U2448, U2449, U2450, U2451, U2452, U2453, U2454, U2455, U2456, U2457, U2458, U2459, U2460, U2461, U2462, U2463, U2464, U2465, U2466, U2467, U2468, U2469, U2470, U2471, U2472, U2473, U2474, U2475, U2476, U2477, U2478, U2479, U2480, U2481, U2482, U2483, U2484, U2485, U2486, U2487, U2488, U2489, U2490, U2491, U2492, U2493, U2494, U2495, U2496, U2497, U2498, U2499, U2500, U2501, U2502, U2503, U2504, U2505, U2506, U2507, U2508, U2509, U2510, U2511, U2512, U2513, U2514, U2515, U2516, U2517, U2518, U2519, U2520, U2521, U2522, U2523, U2524, U2525, U2526, U2527, U2528, U2529, U2530, U2531, U2532, U2533, U2534, U2535, U2536, U2537, U2538, U2539, U2540, U2541, U2542, U2543, U2544, U2545, U2546, U2547, U2548, U2549, U2550, U2551, U2552, U2553, U2554, U2555, U2556, U2557, U2558, U2559, U2560, U2561, U2562, U2563, U2564, U2565, U2566, U2567, U2568, U2569, U2570, U2571, U2572, U2573, U2574, U2575, U2576, U2577, U2578, U2579, U2580, U2581, U2582, U2583, U2584, U2585, U2586, U2587, U2588, U2589, U2590, U2591, U2592, U2593, U2594, U2595, U2596, U2597, U2598, U2599, U2600, U2601, U2602, U2603, U2604, U2605, U2606, U2607, U2608, U2609, U2610, U2611, U2612, U2613, U2614, U2615, U2616, U2617, U2618, U2620, U2621, U2622, U2623, U2624, U2625, U2626, U2627, U2628, U2629, U2630, U2631, U2632, U2633, U2634, U2635, U2636, U2637, U2638, U2639, U2640, U2641, U2642, U2643, U2644, U2645, U2646, U2647, U2648, U2649, U2650, U2651, U2652, U2653, U2654, U2655, U2656, U2657, U2658, U2659, U2660, U2661, U2662, U2663, U2664, U2665, U2666, U2667, U2668, U2669, U2670, U2671, U2672, U2673, U2674, U2675, U2676, U2677, U2678, U2679, U2680, U2681, U2682, U2683, U2684, U2685, U2686, U2687, U2688, U2689, U2690, U2691, U2692, U2693, U2694, U2695, U2696, U2697, U2698, U2699, U2700, U2701, U2702, U2703, U2704, U2705, U2706, U2707, U2708, U2709, U2710, U2711, U2712, U2713, U2714, U2715, U2716, U2717, U2718, U2719, U2720, U2721, U2722, U2723, U2724, U2725, U2726, U2727, U2728, U2729, U2730, U2731, U2732, U2733, U2734, U2735, U2736, U2737, U2738, U2739, U2740, U2741, U2742, U2743, U2744, U2745, U2746, U2747, U2748, U2749, U2750, U2751, U2752, U2753, U2754, U2755, U2756, U2757, U2758, U2759, U2760, U2761, U2762, U2763, U2764, U2765, U2766, U2767, U2768, U2769, U2770, U2771, U2772, U2773, U2774, U2775, U2776, U2777, U2778, U2779, U2780, U2781, U2782, U2783, U2784, U2785, U2786, U2787, U3214, U3215, U3216, U3217, U3218, U3219, U3220, U3221, U3222, U3223, U3224, U3225, U3226, U3227, U3228, U3229, U3230, U3231, U3232, U3233, U3234, U3235, U3236, U3237, U3238, U3239, U3240, U3241, U3242, U3243, U3244, U3245, U3246, U3247, U3248, U3249, U3250, U3251, U3252, U3253, U3254, U3255, U3256, U3257, U3258, U3259, U3260, U3261, U3262, U3263, U3264, U3265, U3266, U3267, U3268, U3269, U3270, U3271, U3272, U3273, U3274, U3275, U3276, U3277, U3278, U3279, U3280, U3281, U3282, U3283, U3284, U3285, U3286, U3287, U3288, U3289, U3290, U3291, U3292, U3293, U3294, U3295, U3296, U3297, U3298, U3299, U3300, U3301, U3302, U3303, U3304, U3305, U3306, U3307, U3308, U3309, U3310, U3311, U3312, U3313, U3314, U3315, U3316, U3317, U3318, U3319, U3320, U3321, U3322, U3323, U3324, U3325, U3326, U3327, U3328, U3329, U3330, U3331, U3332, U3333, U3334, U3335, U3336, U3337, U3338, U3339, U3340, U3341, U3342, U3343, U3344, U3345, U3346, U3347, U3348, U3349, U3350, U3351, U3352, U3353, U3354, U3355, U3356, U3357, U3358, U3359, U3360, U3361, U3362, U3363, U3364, U3365, U3366, U3367, U3368, U3369, U3370, U3371, U3372, U3373, U3374, U3375, U3376, U3377, U3378, U3379, U3380, U3381, U3382, U3383, U3384, U3385, U3386, U3387, U3388, U3389, U3390, U3391, U3392, U3393, U3394, U3395, U3396, U3397, U3398, U3399, U3400, U3401, U3402, U3403, U3404, U3405, U3406, U3407, U3408, U3409, U3410, U3411, U3412, U3413, U3414, U3415, U3416, U3417, U3418, U3419, U3420, U3421, U3422, U3423, U3424, U3425, U3426, U3427, U3428, U3429, U3430, U3431, U3432, U3433, U3434, U3435, U3436, U3437, U3438, U3439, U3440, U3441, U3442, U3443, U3444, U3449, U3450, U3454, U3457, U3458, U3466, U3467, U3475, U3476, U3477, U3478, U3479, U3480, U3481, U3482, U3483, U3484, U3485, U3486, U3487, U3488, U3489, U3490, U3491, U3492, U3493, U3494, U3495, U3496, U3497, U3498, U3499, U3500, U3501, U3502, U3503, U3504, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3582, U3583, U3584, U3585, U3586, U3587, U3588, U3589, U3590, U3591, U3592, U3593, U3594, U3595, U3596, U3597, U3598, U3599, U3600, U3601, U3602, U3603, U3604, U3605, U3606, U3607, U3608, U3609, U3610, U3611, U3612, U3613, U3614, U3615, U3616, U3617, U3618, U3619, U3620, U3621, U3622, U3623, U3624, U3625, U3626, U3627, U3628, U3629, U3630, U3631, U3632, U3633, U3634, U3635, U3636, U3637, U3638, U3639, U3640, U3641, U3642, U3643, U3644, U3645, U3646, U3647, U3648, U3649, U3650, U3651, U3652, U3653, U3654, U3655, U3656, U3657, U3658, U3659, U3660, U3661, U3662, U3663, U3664, U3665, U3666, U3667, U3668, U3669, U3670, U3671, U3672, U3673, U3674, U3675, U3676, U3677, U3678, U3679, U3680, U3681, U3682, U3683, U3684, U3685, U3686, U3687, U3688, U3689, U3690, U3691, U3692, U3693, U3694, U3695, U3696, U3697, U3698, U3699, U3700, U3701, U3702, U3703, U3704, U3705, U3706, U3707, U3708, U3709, U3710, U3711, U3712, U3713, U3714, U3715, U3716, U3717, U3718, U3719, U3720, U3721, U3722, U3723, U3724, U3725, U3726, U3727, U3728, U3729, U3730, U3731, U3732, U3733, U3734, U3735, U3736, U3737, U3738, U3739, U3740, U3741, U3742, U3743, U3744, U3745, U3746, U3747, U3748, U3749, U3750, U3751, U3752, U3753, U3754, U3755, U3756, U3757, U3758, U3759, U3760, U3761, U3762, U3763, U3764, U3765, U3766, U3767, U3768, U3769, U3770, U3771, U3772, U3773, U3774, U3775, U3776, U3777, U3778, U3779, U3780, U3781, U3782, U3783, U3784, U3785, U3786, U3787, U3788, U3789, U3790, U3791, U3792, U3793, U3794, U3795, U3796, U3797, U3798, U3799, U3800, U3801, U3802, U3803, U3804, U3805, U3806, U3807, U3808, U3809, U3810, U3811, U3812, U3813, U3814, U3815, U3816, U3817, U3818, U3819, U3820, U3821, U3822, U3823, U3824, U3825, U3826, U3827, U3828, U3829, U3830, U3831, U3832, U3833, U3834, U3835, U3836, U3837, U3838, U3839, U3840, U3841, U3842, U3843, U3844, U3845, U3846, U3847, U3848, U3849, U3850, U3851, U3852, U3853, U3854, U3855, U3856, U3857, U3858, U3859, U3860, U3861, U3862, U3863, U3864, U3865, U3866, U3867, U3868, U3869, U3870, U3871, U3872, U3873, U3874, U3875, U3876, U3877, U3878, U3879, U3880, U3881, U3882, U3883, U3884, U3885, U3886, U3887, U3888, U3889, U3890, U3891, U3892, U3893, U3894, U3895, U3896, U3897, U3898, U3899, U3900, U3901, U3902, U3903, U3904, U3905, U3906, U3907, U3908, U3909, U3910, U3911, U3912, U3913, U3914, U3915, U3916, U3917, U3918, U3919, U3920, U3921, U3922, U3923, U3924, U3925, U3926, U3927, U3928, U3929, U3930, U3931, U3932, U3933, U3934, U3935, U3936, U3937, U3938, U3939, U3940, U3941, U3942, U3943, U3944, U3945, U3946, U3947, U3948, U3949, U3950, U3951, U3952, U3953, U3954, U3955, U3956, U3957, U3958, U3959, U3960, U3961, U3962, U3963, U3964, U3965, U3966, U3967, U3968, U3969, U3970, U3971, U3972, U3973, U3974, U3975, U3976, U3977, U3978, U3979, U3980, U3981, U3982, U3983, U3984, U3985, U3986, U3987, U3988, U3989, U3990, U3991, U3992, U3993, U3994, U3995, U3996, U3997, U3998, U3999, U4000, U4001, U4002, U4003, U4004, U4005, U4006, U4007, U4008, U4009, U4010, U4011, U4012, U4013, U4014, U4015, U4016, U4017, U4018, U4019, U4020, U4021, U4022, U4023, U4024, U4025, U4026, U4027, U4028, U4029, U4030, U4031, U4032, U4033, U4034, U4035, U4036, U4037, U4038, U4039, U4040, U4041, U4042, U4043, U4044, U4045, U4046, U4047, U4048, U4049, U4050, U4051, U4052, U4053, U4054, U4055, U4056, U4057, U4058, U4059, U4060, U4061, U4062, U4063, U4064, U4065, U4066, U4067, U4068, U4069, U4070, U4071, U4072, U4073, U4074, U4075, U4076, U4077, U4078, U4079, U4080, U4081, U4082, U4083, U4084, U4085, U4086, U4087, U4088, U4089, U4090, U4091, U4092, U4093, U4094, U4095, U4096, U4097, U4098, U4099, U4100, U4101, U4102, U4103, U4104, U4105, U4106, U4107, U4108, U4109, U4110, U4111, U4112, U4113, U4114, U4115, U4116, U4117, U4118, U4119, U4120, U4121, U4122, U4123, U4124, U4125, U4126, U4127, U4128, U4129, U4130, U4131, U4132, U4133, U4134, U4135, U4136, U4137, U4138, U4139, U4140, U4141, U4142, U4143, U4144, U4145, U4146, U4147, U4148, U4149, U4150, U4151, U4152, U4153, U4154, U4155, U4156, U4157, U4158, U4159, U4160, U4161, U4162, U4163, U4164, U4165, U4166, U4167, U4168, U4169, U4170, U4171, U4172, U4173, U4174, U4175, U4176, U4177, U4178, U4179, U4180, U4181, U4182, U4183, U4184, U4185, U4186, U4187, U4188, U4189, U4190, U4191, U4192, U4193, U4194, U4195, U4196, U4197, U4198, U4199, U4200, U4201, U4202, U4203, U4204, U4205, U4206, U4207, U4208, U4209, U4210, U4211, U4212, U4213, U4214, U4215, U4216, U4217, U4218, U4219, U4220, U4221, U4222, U4223, U4224, U4225, U4226, U4227, U4228, U4229, U4230, U4231, U4232, U4233, U4234, U4235, U4236, U4237, U4238, U4239, U4240, U4241, U4242, U4243, U4244, U4245, U4246, U4247, U4248, U4249, U4250, U4251, U4252, U4253, U4254, U4255, U4256, U4257, U4258, U4259, U4260, U4261, U4262, U4263, U4264, U4265, U4266, U4267, U4268, U4269, U4270, U4271, U4272, U4273, U4274, U4275, U4276, U4277, U4278, U4279, U4280, U4281, U4282, U4283, U4284, U4285, U4286, U4287, U4288, U4289, U4290, U4291, U4292, U4293, U4294, U4295, U4296, U4297, U4298, U4299, U4300, U4301, U4302, U4303, U4304, U4305, U4306, U4307, U4308, U4309, U4310, U4311, U4312, U4313, U4314, U4315, U4316, U4317, U4318, U4319, U4320, U4321, U4322, U4323, U4324, U4325, U4326, U4327, U4328, U4329, U4330, U4331, U4332, U4333, U4334, U4335, U4336, U4337, U4338, U4339, U4340, U4341, U4342, U4343, U4344, U4345, U4346, U4347, U4348, U4349, U4350, U4351, U4352, U4353, U4354, U4355, U4356, U4357, U4358, U4359, U4360, U4361, U4362, U4363, U4364, U4365, U4366, U4367, U4368, U4369, U4370, U4371, U4372, U4373, U4374, U4375, U4376, U4377, U4378, U4379, U4380, U4381, U4382, U4383, U4384, U4385, U4386, U4387, U4388, U4389, U4390, U4391, U4392, U4393, U4394, U4395, U4396, U4397, U4398, U4399, U4400, U4401, U4402, U4403, U4404, U4405, U4406, U4407, U4408, U4409, U4410, U4411, U4412, U4413, U4414, U4415, U4416, U4417, U4418, U4419, U4420, U4421, U4422, U4423, U4424, U4425, U4426, U4427, U4428, U4429, U4430, U4431, U4432, U4433, U4434, U4435, U4436, U4437, U4438, U4439, U4440, U4441, U4442, U4443, U4444, U4445, U4446, U4447, U4448, U4449, U4450, U4451, U4452, U4453, U4454, U4455, U4456, U4457, U4458, U4459, U4460, U4461, U4462, U4463, U4464, U4465, U4466, U4467, U4468, U4469, U4470, U4471, U4472, U4473, U4474, U4475, U4476, U4477, U4478, U4479, U4480, U4481, U4482, U4483, U4484, U4485, U4486, U4487, U4488, U4489, U4490, U4491, U4492, U4493, U4494, U4495, U4496, U4497, U4498, U4499, U4500, U4501, U4502, U4503, U4504, U4505, U4506, U4507, U4508, U4509, U4510, U4511, U4512, U4513, U4514, U4515, U4516, U4517, U4518, U4519, U4520, U4521, U4522, U4523, U4524, U4525, U4526, U4527, U4528, U4529, U4530, U4531, U4532, U4533, U4534, U4535, U4536, U4537, U4538, U4539, U4540, U4541, U4542, U4543, U4544, U4545, U4546, U4547, U4548, U4549, U4550, U4551, U4552, U4553, U4554, U4555, U4556, U4557, U4558, U4559, U4560, U4561, U4562, U4563, U4564, U4565, U4566, U4567, U4568, U4569, U4570, U4571, U4572, U4573, U4574, U4575, U4576, U4577, U4578, U4579, U4580, U4581, U4582, U4583, U4584, U4585, U4586, U4587, U4588, U4589, U4590, U4591, U4592, U4593, U4594, U4595, U4596, U4597, U4598, U4599, U4600, U4601, U4602, U4603, U4604, U4605, U4606, U4607, U4608, U4609, U4610, U4611, U4612, U4613, U4614, U4615, U4616, U4617, U4618, U4619, U4620, U4621, U4622, U4623, U4624, U4625, U4626, U4627, U4628, U4629, U4630, U4631, U4632, U4633, U4634, U4635, U4636, U4637, U4638, U4639, U4640, U4641, U4642, U4643, U4644, U4645, U4646, U4647, U4648, U4649, U4650, U4651, U4652, U4653, U4654, U4655, U4656, U4657, U4658, U4659, U4660, U4661, U4662, U4663, U4664, U4665, U4666, U4667, U4668, U4669, U4670, U4671, U4672, U4673, U4674, U4675, U4676, U4677, U4678, U4679, U4680, U4681, U4682, U4683, U4684, U4685, U4686, U4687, U4688, U4689, U4690, U4691, U4692, U4693, U4694, U4695, U4696, U4697, U4698, U4699, U4700, U4701, U4702, U4703, U4704, U4705, U4706, U4707, U4708, U4709, U4710, U4711, U4712, U4713, U4714, U4715, U4716, U4717, U4718, U4719, U4720, U4721, U4722, U4723, U4724, U4725, U4726, U4727, U4728, U4729, U4730, U4731, U4732, U4733, U4734, U4735, U4736, U4737, U4738, U4739, U4740, U4741, U4742, U4743, U4744, U4745, U4746, U4747, U4748, U4749, U4750, U4751, U4752, U4753, U4754, U4755, U4756, U4757, U4758, U4759, U4760, U4761, U4762, U4763, U4764, U4765, U4766, U4767, U4768, U4769, U4770, U4771, U4772, U4773, U4774, U4775, U4776, U4777, U4778, U4779, U4780, U4781, U4782, U4783, U4784, U4785, U4786, U4787, U4788, U4789, U4790, U4791, U4792, U4793, U4794, U4795, U4796, U4797, U4798, U4799, U4800, U4801, U4802, U4803, U4804, U4805, U4806, U4807, U4808, U4809, U4810, U4811, U4812, U4813, U4814, U4815, U4816, U4817, U4818, U4819, U4820, U4821, U4822, U4823, U4824, U4825, U4826, U4827, U4828, U4829, U4830, U4831, U4832, U4833, U4834, U4835, U4836, U4837, U4838, U4839, U4840, U4841, U4842, U4843, U4844, U4845, U4846, U4847, U4848, U4849, U4850, U4851, U4852, U4853, U4854, U4855, U4856, U4857, U4858, U4859, U4860, U4861, U4862, U4863, U4864, U4865, U4866, U4867, U4868, U4869, U4870, U4871, U4872, U4873, U4874, U4875, U4876, U4877, U4878, U4879, U4880, U4881, U4882, U4883, U4884, U4885, U4886, U4887, U4888, U4889, U4890, U4891, U4892, U4893, U4894, U4895, U4896, U4897, U4898, U4899, U4900, U4901, U4902, U4903, U4904, U4905, U4906, U4907, U4908, U4909, U4910, U4911, U4912, U4913, U4914, U4915, U4916, U4917, U4918, U4919, U4920, U4921, U4922, U4923, U4924, U4925, U4926, U4927, U4928, U4929, U4930, U4931, U4932, U4933, U4934, U4935, U4936, U4937, U4938, U4939, U4940, U4941, U4942, U4943, U4944, U4945, U4946, U4947, U4948, U4949, U4950, U4951, U4952, U4953, U4954, U4955, U4956, U4957, U4958, U4959, U4960, U4961, U4962, U4963, U4964, U4965, U4966, U4967, U4968, U4969, U4970, U4971, U4972, U4973, U4974, U4975, U4976, U4977, U4978, U4979, U4980, U4981, U4982, U4983, U4984, U4985, U4986, U4987, U4988, U4989, U4990, U4991, U4992, U4993, U4994, U4995, U4996, U4997, U4998, U4999, U5000, U5001, U5002, U5003, U5004, U5005, U5006, U5007, U5008, U5009, U5010, U5011, U5012, U5013, U5014, U5015, U5016, U5017, U5018, U5019, U5020, U5021, U5022, U5023, U5024, U5025, U5026, U5027, U5028, U5029, U5030, U5031, U5032, U5033, U5034, U5035, U5036, U5037, U5038, U5039, U5040, U5041, U5042, U5043, U5044, U5045, U5046, U5047, U5048, U5049, U5050, U5051, U5052, U5053, U5054, U5055, U5056, U5057, U5058, U5059, U5060, U5061, U5062, U5063, U5064, U5065, U5066, U5067, U5068, U5069, U5070, U5071, U5072, U5073, U5074, U5075, U5076, U5077, U5078, U5079, U5080, U5081, U5082, U5083, U5084, U5085, U5086, U5087, U5088, U5089, U5090, U5091, U5092, U5093, U5094, U5095, U5096, U5097, U5098, U5099, U5100, U5101, U5102, U5103, U5104, U5105, U5106, U5107, U5108, U5109, U5110, U5111, U5112, U5113, U5114, U5115, U5116, U5117, U5118, U5119, U5120, U5121, U5122, U5123, U5124, U5125, U5126, U5127, U5128, U5129, U5130, U5131, U5132, U5133, U5134, U5135, U5136, U5137, U5138, U5139, U5140, U5141, U5142, U5143, U5144, U5145, U5146, U5147, U5148, U5149, U5150, U5151, U5152, U5153, U5154, U5155, U5156, U5157, U5158, U5159, U5160, U5161, U5162, U5163, U5164, U5165, U5166, U5167, U5168, U5169, U5170, U5171, U5172, U5173, U5174, U5175, U5176, U5177, U5178, U5179, U5180, U5181, U5182, U5183, U5184, U5185, U5186, U5187, U5188, U5189, U5190, U5191, U5192, U5193, U5194, U5195, U5196, U5197, U5198, U5199, U5200, U5201, U5202, U5203, U5204, U5205, U5206, U5207, U5208, U5209, U5210, U5211, U5212, U5213, U5214, U5215, U5216, U5217, U5218, U5219, U5220, U5221, U5222, U5223, U5224, U5225, U5226, U5227, U5228, U5229, U5230, U5231, U5232, U5233, U5234, U5235, U5236, U5237, U5238, U5239, U5240, U5241, U5242, U5243, U5244, U5245, U5246, U5247, U5248, U5249, U5250, U5251, U5252, U5253, U5254, U5255, U5256, U5257, U5258, U5259, U5260, U5261, U5262, U5263, U5264, U5265, U5266, U5267, U5268, U5269, U5270, U5271, U5272, U5273, U5274, U5275, U5276, U5277, U5278, U5279, U5280, U5281, U5282, U5283, U5284, U5285, U5286, U5287, U5288, U5289, U5290, U5291, U5292, U5293, U5294, U5295, U5296, U5297, U5298, U5299, U5300, U5301, U5302, U5303, U5304, U5305, U5306, U5307, U5308, U5309, U5310, U5311, U5312, U5313, U5314, U5315, U5316, U5317, U5318, U5319, U5320, U5321, U5322, U5323, U5324, U5325, U5326, U5327, U5328, U5329, U5330, U5331, U5332, U5333, U5334, U5335, U5336, U5337, U5338, U5339, U5340, U5341, U5342, U5343, U5344, U5345, U5346, U5347, U5348, U5349, U5350, U5351, U5352, U5353, U5354, U5355, U5356, U5357, U5358, U5359, U5360, U5361, U5362, U5363, U5364, U5365, U5366, U5367, U5368, U5369, U5370, U5371, U5372, U5373, U5374, U5375, U5376, U5377, U5378, U5379, U5380, U5381, U5382, U5383, U5384, U5385, U5386, U5387, U5388, U5389, U5390, U5391, U5392, U5393, U5394, U5395, U5396, U5397, U5398, U5399, U5400, U5401, U5402, U5403, U5404, U5405, U5406, U5407, U5408, U5409, U5410, U5411, U5412, U5413, U5414, U5415, U5416, U5417, U5418, U5419, U5420, U5421, U5422, U5423, U5424, U5425, U5426, U5427, U5428, U5429, U5430, U5431, U5432, U5433, U5434, U5435, U5436, U5437, U5438, U5439, U5440, U5441, U5442, U5443, U5444, U5445, U5446, U5447, U5448, U5449, U5450, U5451, U5452, U5453, U5454, U5455, U5456, U5457, U5458, U5459, U5460, U5461, U5462, U5463, U5464, U5465, U5466, U5467, U5468, U5469, U5470, U5471, U5472, U5473, U5474, U5475, U5476, U5477, U5478, U5479, U5480, U5481, U5482, U5483, U5484, U5485, U5486, U5487, U5488, U5489, U5490, U5491, U5492, U5493, U5494, U5495, U5496, U5497, U5498, U5499, U5500, U5501, U5502, U5503, U5504, U5505, U5506, U5507, U5508, U5509, U5510, U5511, U5512, U5513, U5514, U5515, U5516, U5517, U5518, U5519, U5520, U5521, U5522, U5523, U5524, U5525, U5526, U5527, U5528, U5529, U5530, U5531, U5532, U5533, U5534, U5535, U5536, U5537, U5538, U5539, U5540, U5541, U5542, U5543, U5544, U5545, U5546, U5547, U5548, U5549, U5550, U5551, U5552, U5553, U5554, U5555, U5556, U5557, U5558, U5559, U5560, U5561, U5562, U5563, U5564, U5565, U5566, U5567, U5568, U5569, U5570, U5571, U5572, U5573, U5574, U5575, U5576, U5577, U5578, U5579, U5580, U5581, U5582, U5583, U5584, U5585, U5586, U5587, U5588, U5589, U5590, U5591, U5592, U5593, U5594, U5595, U5596, U5597, U5598, U5599, U5600, U5601, U5602, U5603, U5604, U5605, U5606, U5607, U5608, U5609, U5610, U5611, U5612, U5613, U5614, U5615, U5616, U5617, U5618, U5619, U5620, U5621, U5622, U5623, U5624, U5625, U5626, U5627, U5628, U5629, U5630, U5631, U5632, U5633, U5634, U5635, U5636, U5637, U5638, U5639, U5640, U5641, U5642, U5643, U5644, U5645, U5646, U5647, U5648, U5649, U5650, U5651, U5652, U5653, U5654, U5655, U5656, U5657, U5658, U5659, U5660, U5661, U5662, U5663, U5664, U5665, U5666, U5667, U5668, U5669, U5670, U5671, U5672, U5673, U5674, U5675, U5676, U5677, U5678, U5679, U5680, U5681, U5682, U5683, U5684, U5685, U5686, U5687, U5688, U5689, U5690, U5691, U5692, U5693, U5694, U5695, U5696, U5697, U5698, U5699, U5700, U5701, U5702, U5703, U5704, U5705, U5706, U5707, U5708, U5709, U5710, U5711, U5712, U5713, U5714, U5715, U5716, U5717, U5718, U5719, U5720, U5721, U5722, U5723, U5724, U5725, U5726, U5727, U5728, U5729, U5730, U5731, U5732, U5733, U5734, U5735, U5736, U5737, U5738, U5739, U5740, U5741, U5742, U5743, U5744, U5745, U5746, U5747, U5748, U5749, U5750, U5751, U5752, U5753, U5754, U5755, U5756, U5757, U5758, U5759, U5760, U5761, U5762, U5763, U5764, U5765, U5766, U5767, U5768, U5769, U5770, U5771, U5772, U5773, U5774, U5775, U5776, U5777, U5778, U5779, U5780, U5781, U5782, U5783, U5784, U5785, U5786, U5787, U5788, U5789, U5790, U5791, U5792, U5793, U5794, U5795, U5796, U5797, U5798, U5799, U5800, U5801, U5802, U5803, U5804, U5805, U5806, U5807, U5808, U5809, U5810, U5811, U5812, U5813, U5814, U5815, U5816, U5817, U5818, U5819, U5820, U5821, U5822, U5823, U5824, U5825, U5826, U5827, U5828, U5829, U5830, U5831, U5832, U5833, U5834, U5835, U5836, U5837, U5838, U5839, U5840, U5841, U5842, U5843, U5844, U5845, U5846, U5847, U5848, U5849, U5850, U5851, U5852, U5853, U5854, U5855, U5856, U5857, U5858, U5859, U5860, U5861, U5862, U5863, U5864, U5865, U5866, U5867, U5868, U5869, U5870, U5871, U5872, U5873, U5874, U5875, U5876, U5877, U5878, U5879, U5880, U5881, U5882, U5883, U5884, U5885, U5886, U5887, U5888, U5889, U5890, U5891, U5892, U5893, U5894, U5895, U5896, U5897, U5898, U5899, U5900, U5901, U5902, U5903, U5904, U5905, U5906, U5907, U5908, U5909, U5910, U5911, U5912, U5913, U5914, U5915, U5916, U5917, U5918, U5919, U5920, U5921, U5922, U5923, U5924, U5925, U5926, U5927, U5928, U5929, U5930, U5931, U5932, U5933, U5934, U5935, U5936, U5937, U5938, U5939, U5940, U5941, U5942, U5943, U5944, U5945, U5946, U5947, U5948, U5949, U5950, U5951, U5952, U5953, U5954, U5955, U5956, U5957, U5958, U5959, U5960, U5961, U5962, U5963, U5964, U5965, U5966, U5967, U5968, U5969, U5970, U5971, U5972, U5973, U5974, U5975, U5976, U5977, U5978, U5979, U5980, U5981, U5982, U5983, U5984, U5985, U5986, U5987, U5988, U5989, U5990, U5991, U5992, U5993, U5994, U5995, U5996, U5997, U5998, U5999, U6000, U6001, U6002, U6003, U6004, U6005, U6006, U6007, U6008, U6009, U6010, U6011, U6012, U6013, U6014, U6015, U6016, U6017, U6018, U6019, U6020, U6021, U6022, U6023, U6024, U6025, U6026, U6027, U6028, U6029, U6030, U6031, U6032, U6033, U6034, U6035, U6036, U6037, U6038, U6039, U6040, U6041, U6042, U6043, U6044, U6045, U6046, U6047, U6048, U6049, U6050, U6051, U6052, U6053, U6054, U6055, U6056, U6057, U6058, U6059, U6060, U6061, U6062, U6063, U6064, U6065, U6066, U6067, U6068, U6069, U6070, U6071, U6072, U6073, U6074, U6075, U6076, U6077, U6078, U6079, U6080, U6081, U6082, U6083, U6084, U6085, U6086, U6087, U6088, U6089, U6090, U6091, U6092, U6093, U6094, U6095, U6096, U6097, U6098, U6099, U6100, U6101, U6102, U6103, U6104, U6105, U6106, U6107, U6108, U6109, U6110, U6111, U6112, U6113, U6114, U6115, U6116, U6117, U6118, U6119, U6120, U6121, U6122, U6123, U6124, U6125, U6126, U6127, U6128, U6129, U6130, U6131, U6132, U6133, U6134, U6135, U6136, U6137, U6138, U6139, U6140, U6141, U6142, U6143, U6144, U6145, U6146, U6147, U6148, U6149, U6150, U6151, U6152, U6153, U6154, U6155, U6156, U6157, U6158, U6159, U6160, U6161, U6162, U6163, U6164, U6165, U6166, U6167, U6168, U6169, U6170, U6171, U6172, U6173, U6174, U6175, U6176, U6177, U6178, U6179, U6180, U6181, U6182, U6183, U6184, U6185, U6186, U6187, U6188, U6189, U6190, U6191, U6192, U6193, U6194, U6195, U6196, U6197, U6198, U6199, U6200, U6201, U6202, U6203, U6204, U6205, U6206, U6207, U6208, U6209, U6210, U6211, U6212, U6213, U6214, U6215, U6216, U6217, U6218, U6219, U6220, U6221, U6222, U6223, U6224, U6225, U6226, U6227, U6228, U6229, U6230, U6231, U6232, U6233, U6234, U6235, U6236, U6237, U6238, U6239, U6240, U6241, U6242, U6243, U6244, U6245, U6246, U6247, U6248, U6249, U6250, U6251, U6252, U6253, U6254, U6255, U6256, U6257, U6258, U6259, U6260, U6261, U6262, U6263, U6264, U6265, U6266, U6267, U6268, U6269, U6270, U6271, U6272, U6273, U6274, U6275, U6276, U6277, U6278, U6279, U6280, U6281, U6282, U6283, U6284, U6285, U6286, U6287, U6288, U6289, U6290, U6291, U6292, U6293, U6294, U6295, U6296, U6297, U6298, U6299, U6300, U6301, U6302, U6303, U6304, U6305, U6306, U6307, U6308, U6309, U6310, U6311, U6312, U6313, U6314, U6315, U6316, U6317, U6318, U6319, U6320, U6321, U6322, U6323, U6324, U6325, U6326, U6327, U6328, U6329, U6330, U6331, U6332, U6333, U6334, U6335, U6336, U6337, U6338, U6339, U6340, U6341, U6342, U6343, U6344, U6345, U6346, U6347, U6348, U6349, U6350, U6351, U6352, U6353, U6354, U6355, U6356, U6357, U6358, U6359, U6360, U6361, U6362, U6363, U6364, U6365, U6366, U6367, U6368, U6369, U6370, U6371, U6372, U6373, U6374, U6375, U6376, U6377, U6378, U6379, U6380, U6381, U6382, U6383, U6384, U6385, U6386, U6387, U6388, U6389, U6390, U6391, U6392, U6393, U6394, U6395, U6396, U6397, U6398, U6399, U6400, U6401, U6402, U6403, U6404, U6405, U6406, U6407, U6408, U6409, U6410, U6411, U6412, U6413, U6414, U6415, U6416, U6417, U6418, U6419, U6420, U6421, U6422, U6423, U6424, U6425, U6426, U6427, U6428, U6429, U6430, U6431, U6432, U6433, U6434, U6435, U6436, U6437, U6438, U6439, U6440, U6441, U6442, U6443, U6444, U6445, U6446, U6447, U6448, U6449, U6450, U6451, U6452, U6453, U6454, U6455, U6456, U6457, U6458, U6459, U6460, U6461, U6462, U6463, U6464, U6465, U6466, U6467, U6468, U6469, U6470, U6471, U6472, U6473, U6474, U6475, U6476, U6477, U6478, U6479, U6480, U6481, U6482, U6483, U6484, U6485, U6486, U6487, U6488, U6489, U6490, U6491, U6492, U6493, U6494, U6495, U6496, U6497, U6498, U6499, U6500, U6501, U6502, U6503, U6504, U6505, U6506, U6507, U6508, U6509, U6510, U6511, U6512, U6513, U6514, U6515, U6516, U6517, U6518, U6519, U6520, U6521, U6522, U6523, U6524, U6525, U6526, U6527, U6528, U6529, U6530, U6531, U6532, U6533, U6534, U6535, U6536, U6537, U6538, U6539, U6540, U6541, U6542, U6543, U6544, U6545, U6546, U6547, U6548, U6549, U6550, U6551, U6552, U6553, U6554, U6555, U6556, U6557, U6558, U6559, U6560, U6561, U6562, U6563, U6564, U6565, U6566, U6567, U6568, U6569, U6570, U6571, U6572, U6573, U6574, U6575, U6576, U6577, U6578, U6579, U6580, U6581, U6582, U6583, U6584, U6585, U6586, U6587, U6588, U6589, U6590, U6591, U6592, U6593, U6594, U6595, U6596, U6597, U6598, U6599, U6600, U6601, U6602, U6603, U6604, U6605, U6606, U6607, U6608, U6609, U6610, U6611, U6612, U6613, U6614, U6615, U6616, U6617, U6618, U6619, U6620, U6621, U6622, U6623, U6624, U6625, U6626, U6627, U6628, U6629, U6630, U6631, U6632, U6633, U6634, U6635, U6636, U6637, U6638, U6639, U6640, U6641, U6642, U6643, U6644, U6645, U6646, U6647, U6648, U6649, U6650, U6651, U6652, U6653, U6654, U6655, U6656, U6657, U6658, U6659, U6660, U6661, U6662, U6663, U6664, U6665, U6666, U6667, U6668, U6669, U6670, U6671, U6672, U6673, U6674, U6675, U6676, U6677, U6678, U6679, U6680, U6681, U6682, U6683, U6684, U6685, U6686, U6687, U6688, U6689, U6690, U6691, U6692, U6693, U6694, U6695, U6696, U6697, U6698, U6699, U6700, U6701, U6702, U6703, U6704, U6705, U6706, U6707, U6708, U6709, U6710, U6711, U6712, U6713, U6714, U6715, U6716, U6717, U6718, U6719, U6720, U6721, U6722, U6723, U6724, U6725, U6726, U6727, U6728, U6729, U6730, U6731, U6732, U6733, U6734, U6735, U6736, U6737, U6738, U6739, U6740, U6741, U6742, U6743, U6744, U6745, U6746, U6747, U6748, U6749, U6750, U6751, U6752, U6753, U6754, U6755, U6756, U6757, U6758, U6759, U6760, U6761, U6762, U6763, U6764, U6765, U6766, U6767, U6768, U6769, U6770, U6771, U6772, U6773, U6774, U6775, U6776, U6777, U6778, U6779, U6780, U6781, U6782, U6783, U6784, U6785, U6786, U6787, U6788, U6789, U6790, U6791, U6792, U6793, U6794, U6795, U6796, U6797, U6798, U6799, U6800, U6801, U6802, U6803, U6804, U6805, U6806, U6807, U6808, U6809, U6810, U6811, U6812, U6813, U6814, U6815, U6816, U6817, U6818, U6819, U6820, U6821, U6822, U6823, U6824, U6825, U6826, U6827, U6828, U6829, U6830, U6831, U6832, U6833, U6834, U6835, U6836, U6837, U6838, U6839, U6840, U6841, U6842, U6843, U6844, U6845, U6846, U6847, U6848, U6849, U6850, U6851, U6852, U6853, U6854, U6855, U6856, U6857, U6858, U6859, U6860, U6861, U6862, U6863, U6864, U6865, U6866, U6867, U6868, U6869, U6870, U6871, U6872, U6873, U6874, U6875, U6876, U6877, U6878, U6879, U6880, U6881, U6882, U6883, U6884, U6885, U6886, U6887, U6888, U6889, U6890, U6891, U6892, U6893, U6894, U6895, U6896, U6897, U6898, U6899, U6900, U6901, U6902, U6903, U6904, U6905, U6906, U6907, U6908, U6909, U6910, U6911, U6912, U6913, U6914, U6915, U6916, U6917, U6918, U6919, U6920, U6921, U6922, U6923, U6924, U6925, U6926, U6927, U6928, U6929, U6930, U6931, U6932, U6933, U6934, U6935, U6936, U6937, U6938, U6939, U6940, U6941, U6942, U6943, U6944, U6945, U6946, U6947, U6948, U6949, U6950, U6951, U6952, U6953, U6954, U6955, U6956, U6957, U6958, U6959, U6960, U6961, U6962, U6963, U6964, U6965, U6966, U6967, U6968, U6969, U6970, U6971, U6972, U6973, U6974, U6975, U6976, U6977, U6978, U6979, U6980, U6981, U6982, U6983, U6984, U6985, U6986, U6987, U6988, U6989, U6990, U6991, U6992, U6993, U6994, U6995, U6996, U6997, U6998, U6999, U7000, U7001, U7002, U7003, U7004, U7005, U7006, U7007, U7008, U7009, U7010, U7011, U7012, U7013, U7014, U7015, U7016, U7017, U7018, U7019, U7020, U7021, U7022, U7023, U7024, U7025, U7026, U7027, U7028, U7029, U7030, U7031, U7032, U7033, U7034, U7035, U7036, U7037, U7038, U7039, U7040, U7041, U7042, U7043, U7044, U7045, U7046, U7047, U7048, U7049, U7050, U7051, U7052, U7053, U7054, U7055, U7056, U7057, U7058, U7059, U7060, U7061, U7062, U7063, U7064, U7065, U7066, U7067, U7068, U7069, U7070, U7071, U7072, U7073, U7074, U7075, U7076, U7077, U7078, U7079, U7080, U7081, U7082, U7083, U7084, U7085, U7086, U7087, U7088, U7089, U7090, U7091, U7092, U7093, U7094, U7095, U7096, U7097, U7098, U7099, U7100, U7101, U7102, U7103, U7104, U7105, U7106, U7107, U7108, U7109, U7110, U7111, U7112, U7113, U7114, U7115, U7116, U7117, U7118, U7119, U7120, U7121, U7122, U7123, U7124, U7125, U7126, U7127, U7128, U7129, U7130, U7131, U7132, U7133, U7134, U7135, U7136, U7137, U7138, U7139, U7140, U7141, U7142, U7143, U7144, U7145, U7146, U7147, U7148, U7149, U7150, U7151, U7152, U7153, U7154, U7155, U7156, U7157, U7158, U7159, U7160, U7161, U7162, U7163, U7164, U7165, U7166, U7167, U7168, U7169, U7170, U7171, U7172, U7173, U7174, U7175, U7176, U7177, U7178, U7179, U7180, U7181, U7182, U7183, U7184, U7185, U7186, U7187, U7188, U7189, U7190, U7191, U7192, U7193, U7194, U7195, U7196, U7197, U7198, U7199, U7200, U7201, U7202, U7203, U7204, U7205, U7206, U7207, U7208, U7209, U7210, U7211, U7212, U7213, U7214, U7215, U7216, U7217, U7218, U7219, U7220, U7221, U7222, U7223, U7224, U7225, U7226, U7227, U7228, U7229, U7230, U7231, U7232, U7233, U7234, U7235, U7236, U7237, U7238, U7239, U7240, U7241, U7242, U7243, U7244, U7245, U7246, U7247, U7248, U7249, U7250, U7251, U7252, U7253, U7254, U7255, U7256, U7257, U7258, U7259, U7260, U7261, U7262, U7263, U7264, U7265, U7266, U7267, U7268, U7269, U7270, U7271, U7272, U7273, U7274, U7275, U7276, U7277, U7278, U7279, U7280, U7281, U7282, U7283, U7284, U7285, U7286, U7287, U7288, U7289, U7290, U7291, U7292, U7293, U7294, U7295, U7296, U7297, U7298, U7299, U7300, U7301, U7302, U7303, U7304, U7305, U7306, U7307, U7308, U7309, U7310, U7311, U7312, U7313, U7314, U7315, U7316, U7317, U7318, U7319, U7320, U7321, U7322, U7323, U7324, U7325, U7326, U7327, U7328, U7329, U7330, U7331, U7332, U7333, U7334, U7335, U7336, U7337, U7338, U7339, U7340, U7341, U7342, U7343, U7344, U7345, U7346, U7347, U7348, U7349, U7350, U7351, U7352, U7353, U7354, U7355, U7356, U7357, U7358, U7359, U7360, U7361, U7362, U7363, U7364, U7365, U7366, U7367, U7368, U7369, U7370, U7371, U7372, U7373, U7374, U7375, U7376, U7377, U7378, U7379, U7380, U7381, U7382, U7383, U7384, U7385, U7386, U7387, U7388, U7389, U7390, U7391, U7392, U7393, U7394, U7395, U7396, U7397, U7398, U7399, U7400, U7401, U7402, U7403, U7404, U7405, U7406, U7407, U7408, U7409, U7410, U7411, U7412, U7413, U7414, U7415, U7416, U7417, U7418, U7419, U7420, U7421, U7422, U7423, U7424, U7425, U7426, U7427, U7428, U7429, U7430, U7431, U7432, U7433, U7434, U7435, U7436, U7437, U7438, U7439, U7440, U7441, U7442, U7443, U7444, U7445, U7446, U7447, U7448, U7449, U7450, U7451, U7452, U7453, U7454, U7455, U7456, U7457, U7458, U7459, U7460, U7461, U7462, U7463, U7464, U7465, U7466, U7467, U7468, U7469, U7470, U7471, U7472, U7473, U7474, U7475, U7476, U7477, U7478, U7479, U7480, U7481, U7482, U7483, U7484, U7485, U7486, U7487, U7488, U7489, U7490, U7491, U7492, U7493, U7494, U7495, U7496, U7497, U7498, U7499, U7500, U7501, U7502, U7503, U7504, U7505, U7506, U7507, U7508, U7509, U7510, U7511, U7512, U7513, U7514, U7515, U7516, U7517, U7518, U7519, U7520, U7521, U7522, U7523, U7524, U7525, U7526, U7527, U7528, U7529, U7530, U7531, U7532, U7533, U7534, U7535, U7536, U7537, U7538, U7539, U7540, U7541, U7542, U7543, U7544, U7545, U7546, U7547, U7548, U7549, U7550, U7551, U7552, U7553, U7554, U7555, U7556, U7557, U7558, U7559, U7560, U7561, U7562, U7563, U7564, U7565, U7566, U7567, U7568, U7569, U7570, U7571, U7572, U7573, U7574, U7575, U7576, U7577, U7578, U7579, U7580, U7581, U7582, U7583, U7584, U7585, U7586, U7587, U7588, U7589, U7590, U7591, U7592, U7593, U7594, U7595, U7596, U7597, U7598, U7599, U7600, U7601, U7602, U7603, U7604, U7605, U7606, U7607, U7608, U7609, U7610, U7611, U7612, U7613, U7614, U7615, U7616, U7617, U7618, U7619, U7620, U7621, U7622, U7623, U7624, U7625, U7626, U7627, U7628, U7629, U7630, U7631, U7632, U7633, U7634, U7635, U7636, U7637, U7638, U7639, U7640, U7641, U7642, U7643, U7644, U7645, U7646, U7647, U7648, U7649, U7650, U7651, U7652, U7653, U7654, U7655, U7656, U7657, U7658, U7659, U7660, U7661, U7662, U7663, U7664, U7665, U7666, U7667, U7668, U7669, U7670, U7671, U7672, U7673, U7674, U7675, U7676, U7677, U7678, U7679, U7680, U7681, U7682, U7683, U7684, U7685, U7686, U7687, U7688, U7689, U7690, U7691, U7692, U7693, U7694, U7695, U7696, U7697, U7698, U7699, U7700, U7701, U7702, U7703, U7704, U7705, U7706, U7707, U7708, U7709, U7710, U7711, U7712, U7713, U7714, U7715, U7716, U7717, U7718, U7719, U7720, U7721, U7722, U7723, U7724, U7725, U7726, U7727, U7728, U7729, U7730, U7731, U7732, U7733, U7734, U7735, U7736, U7737, U7738, U7739, U7740, U7741, U7742, U7743, U7744, U7745, U7746, U7747, U7748, U7749, U7750, U7751, U7752, U7753, U7754, U7755, U7756, U7757, U7758, U7759, U7760, U7761, U7762, U7763, U7764, U7765, U7766, U7767, U7768, U7769, U7770, U7771, U7772, U7773, U7774, U7775, U7776, U7777, U7778, U7779, U7780, U7781, U7782, R2027_U5, R2027_U6, R2027_U7, R2027_U8, R2027_U9, R2027_U10, R2027_U11, R2027_U12, R2027_U13, R2027_U14, R2027_U15, R2027_U16, R2027_U17, R2027_U18, R2027_U19, R2027_U20, R2027_U21, R2027_U22, R2027_U23, R2027_U24, R2027_U25, R2027_U26, R2027_U27, R2027_U28, R2027_U29, R2027_U30, R2027_U31, R2027_U32, R2027_U33, R2027_U34, R2027_U35, R2027_U36, R2027_U37, R2027_U38, R2027_U39, R2027_U40, R2027_U41, R2027_U42, R2027_U43, R2027_U44, R2027_U45, R2027_U46, R2027_U47, R2027_U48, R2027_U49, R2027_U50, R2027_U51, R2027_U52, R2027_U53, R2027_U54, R2027_U55, R2027_U56, R2027_U57, R2027_U58, R2027_U59, R2027_U60, R2027_U61, R2027_U62, R2027_U63, R2027_U64, R2027_U65, R2027_U66, R2027_U67, R2027_U68, R2027_U69, R2027_U70, R2027_U71, R2027_U72, R2027_U73, R2027_U74, R2027_U75, R2027_U76, R2027_U77, R2027_U78, R2027_U79, R2027_U80, R2027_U81, R2027_U82, R2027_U83, R2027_U84, R2027_U85, R2027_U86, R2027_U87, R2027_U88, R2027_U89, R2027_U90, R2027_U91, R2027_U92, R2027_U93, R2027_U94, R2027_U95, R2027_U96, R2027_U97, R2027_U98, R2027_U99, R2027_U100, R2027_U101, R2027_U102, R2027_U103, R2027_U104, R2027_U105, R2027_U106, R2027_U107, R2027_U108, R2027_U109, R2027_U110, R2027_U111, R2027_U112, R2027_U113, R2027_U114, R2027_U115, R2027_U116, R2027_U117, R2027_U118, R2027_U119, R2027_U120, R2027_U121, R2027_U122, R2027_U123, R2027_U124, R2027_U125, R2027_U126, R2027_U127, R2027_U128, R2027_U129, R2027_U130, R2027_U131, R2027_U132, R2027_U133, R2027_U134, R2027_U135, R2027_U136, R2027_U137, R2027_U138, R2027_U139, R2027_U140, R2027_U141, R2027_U142, R2027_U143, R2027_U144, R2027_U145, R2027_U146, R2027_U147, R2027_U148, R2027_U149, R2027_U150, R2027_U151, R2027_U152, R2027_U153, R2027_U154, R2027_U155, R2027_U156, R2027_U157, R2027_U158, R2027_U159, R2027_U160, R2027_U161, R2027_U162, R2027_U163, R2027_U164, R2027_U165, R2027_U166, R2027_U167, R2027_U168, R2027_U169, R2027_U170, R2027_U171, R2027_U172, R2027_U173, R2027_U174, R2027_U175, R2027_U176, R2027_U177, R2027_U178, R2027_U179, R2027_U180, R2027_U181, R2027_U182, R2027_U183, R2027_U184, R2027_U185, R2027_U186, R2027_U187, R2027_U188, R2027_U189, R2027_U190, R2027_U191, R2027_U192, R2027_U193, R2027_U194, R2027_U195, R2027_U196, R2027_U197, R2027_U198, R2027_U199, R2027_U200, R2027_U201, R2027_U202, R2278_U5, R2278_U6, R2278_U7, R2278_U8, R2278_U9, R2278_U10, R2278_U11, R2278_U12, R2278_U13, R2278_U14, R2278_U15, R2278_U16, R2278_U17, R2278_U18, R2278_U19, R2278_U20, R2278_U21, R2278_U22, R2278_U23, R2278_U24, R2278_U25, R2278_U26, R2278_U27, R2278_U28, R2278_U29, R2278_U30, R2278_U31, R2278_U32, R2278_U33, R2278_U34, R2278_U35, R2278_U36, R2278_U37, R2278_U38, R2278_U39, R2278_U40, R2278_U41, R2278_U42, R2278_U43, R2278_U44, R2278_U45, R2278_U46, R2278_U47, R2278_U48, R2278_U49, R2278_U50, R2278_U51, R2278_U52, R2278_U53, R2278_U54, R2278_U55, R2278_U56, R2278_U57, R2278_U58, R2278_U59, R2278_U60, R2278_U61, R2278_U62, R2278_U63, R2278_U64, R2278_U65, R2278_U66, R2278_U67, R2278_U68, R2278_U69, R2278_U70, R2278_U71, R2278_U72, R2278_U73, R2278_U74, R2278_U75, R2278_U76, R2278_U77, R2278_U78, R2278_U79, R2278_U80, R2278_U81, R2278_U82, R2278_U83, R2278_U84, R2278_U85, R2278_U86, R2278_U87, R2278_U88, R2278_U89, R2278_U90, R2278_U91, R2278_U92, R2278_U93, R2278_U94, R2278_U95, R2278_U96, R2278_U97, R2278_U98, R2278_U99, R2278_U100, R2278_U101, R2278_U102, R2278_U103, R2278_U104, R2278_U105, R2278_U106, R2278_U107, R2278_U108, R2278_U109, R2278_U110, R2278_U111, R2278_U112, R2278_U113, R2278_U114, R2278_U115, R2278_U116, R2278_U117, R2278_U118, R2278_U119, R2278_U120, R2278_U121, R2278_U122, R2278_U123, R2278_U124, R2278_U125, R2278_U126, R2278_U127, R2278_U128, R2278_U129, R2278_U130, R2278_U131, R2278_U132, R2278_U133, R2278_U134, R2278_U135, R2278_U136, R2278_U137, R2278_U138, R2278_U139, R2278_U140, R2278_U141, R2278_U142, R2278_U143, R2278_U144, R2278_U145, R2278_U146, R2278_U147, R2278_U148, R2278_U149, R2278_U150, R2278_U151, R2278_U152, R2278_U153, R2278_U154, R2278_U155, R2278_U156, R2278_U157, R2278_U158, R2278_U159, R2278_U160, R2278_U161, R2278_U162, R2278_U163, R2278_U164, R2278_U165, R2278_U166, R2278_U167, R2278_U168, R2278_U169, R2278_U170, R2278_U171, R2278_U172, R2278_U173, R2278_U174, R2278_U175, R2278_U176, R2278_U177, R2278_U178, R2278_U179, R2278_U180, R2278_U181, R2278_U182, R2278_U183, R2278_U184, R2278_U185, R2278_U186, R2278_U187, R2278_U188, R2278_U189, R2278_U190, R2278_U191, R2278_U192, R2278_U193, R2278_U194, R2278_U195, R2278_U196, R2278_U197, R2278_U198, R2278_U199, R2278_U200, R2278_U201, R2278_U202, R2278_U203, R2278_U204, R2278_U205, R2278_U206, R2278_U207, R2278_U208, R2278_U209, R2278_U210, R2278_U211, R2278_U212, R2278_U213, R2278_U214, R2278_U215, R2278_U216, R2278_U217, R2278_U218, R2278_U219, R2278_U220, R2278_U221, R2278_U222, R2278_U223, R2278_U224, R2278_U225, R2278_U226, R2278_U227, R2278_U228, R2278_U229, R2278_U230, R2278_U231, R2278_U232, R2278_U233, R2278_U234, R2278_U235, R2278_U236, R2278_U237, R2278_U238, R2278_U239, R2278_U240, R2278_U241, R2278_U242, R2278_U243, R2278_U244, R2278_U245, R2278_U246, R2278_U247, R2278_U248, R2278_U249, R2278_U250, R2278_U251, R2278_U252, R2278_U253, R2278_U254, R2278_U255, R2278_U256, R2278_U257, R2278_U258, R2278_U259, R2278_U260, R2278_U261, R2278_U262, R2278_U263, R2278_U264, R2278_U265, R2278_U266, R2278_U267, R2278_U268, R2278_U269, R2278_U270, R2278_U271, R2278_U272, R2278_U273, R2278_U274, R2278_U275, R2278_U276, R2278_U277, R2278_U278, R2278_U279, R2278_U280, R2278_U281, R2278_U282, R2278_U283, R2278_U284, R2278_U285, R2278_U286, R2278_U287, R2278_U288, R2278_U289, R2278_U290, R2278_U291, R2278_U292, R2278_U293, R2278_U294, R2278_U295, R2278_U296, R2278_U297, R2278_U298, R2278_U299, R2278_U300, R2278_U301, R2278_U302, R2278_U303, R2278_U304, R2278_U305, R2278_U306, R2278_U307, R2278_U308, R2278_U309, R2278_U310, R2278_U311, R2278_U312, R2278_U313, R2278_U314, R2278_U315, R2278_U316, R2278_U317, R2278_U318, R2278_U319, R2278_U320, R2278_U321, R2278_U322, R2278_U323, R2278_U324, R2278_U325, R2278_U326, R2278_U327, R2278_U328, R2278_U329, R2278_U330, R2278_U331, R2278_U332, R2278_U333, R2278_U334, R2278_U335, R2278_U336, R2278_U337, R2278_U338, R2278_U339, R2278_U340, R2278_U341, R2278_U342, R2278_U343, R2278_U344, R2278_U345, R2278_U346, R2278_U347, R2278_U348, R2278_U349, R2278_U350, R2278_U351, R2278_U352, R2278_U353, R2278_U354, R2278_U355, R2278_U356, R2278_U357, R2278_U358, R2278_U359, R2278_U360, R2278_U361, R2278_U362, R2278_U363, R2278_U364, R2278_U365, R2278_U366, R2278_U367, R2278_U368, R2278_U369, R2278_U370, R2278_U371, R2278_U372, R2278_U373, R2278_U374, R2278_U375, R2278_U376, R2278_U377, R2278_U378, R2278_U379, R2278_U380, R2278_U381, R2278_U382, R2278_U383, R2278_U384, R2278_U385, R2278_U386, R2278_U387, R2278_U388, R2278_U389, R2278_U390, R2278_U391, R2278_U392, R2278_U393, R2278_U394, R2278_U395, R2278_U396, R2278_U397, R2278_U398, R2278_U399, R2278_U400, R2278_U401, R2278_U402, R2278_U403, R2278_U404, R2278_U405, R2278_U406, R2278_U407, R2278_U408, R2278_U409, R2278_U410, R2278_U411, R2278_U412, R2278_U413, R2278_U414, R2278_U415, R2278_U416, R2278_U417, R2278_U418, R2278_U419, R2278_U420, R2278_U421, R2278_U422, R2358_U5, R2358_U6, R2358_U7, R2358_U8, R2358_U9, R2358_U10, R2358_U11, R2358_U12, R2358_U13, R2358_U14, R2358_U15, R2358_U16, R2358_U17, R2358_U18, R2358_U19, R2358_U20, R2358_U21, R2358_U22, R2358_U23, R2358_U24, R2358_U25, R2358_U26, R2358_U27, R2358_U28, R2358_U29, R2358_U30, R2358_U31, R2358_U32, R2358_U33, R2358_U34, R2358_U35, R2358_U36, R2358_U37, R2358_U38, R2358_U39, R2358_U40, R2358_U41, R2358_U42, R2358_U43, R2358_U44, R2358_U45, R2358_U46, R2358_U47, R2358_U48, R2358_U49, R2358_U50, R2358_U51, R2358_U52, R2358_U53, R2358_U54, R2358_U55, R2358_U56, R2358_U57, R2358_U58, R2358_U59, R2358_U60, R2358_U61, R2358_U62, R2358_U63, R2358_U64, R2358_U65, R2358_U66, R2358_U67, R2358_U68, R2358_U69, R2358_U70, R2358_U71, R2358_U72, R2358_U73, R2358_U74, R2358_U75, R2358_U76, R2358_U77, R2358_U78, R2358_U79, R2358_U80, R2358_U81, R2358_U82, R2358_U83, R2358_U84, R2358_U85, R2358_U86, R2358_U87, R2358_U88, R2358_U89, R2358_U90, R2358_U91, R2358_U92, R2358_U93, R2358_U94, R2358_U95, R2358_U96, R2358_U97, R2358_U98, R2358_U99, R2358_U100, R2358_U101, R2358_U102, R2358_U103, R2358_U104, R2358_U105, R2358_U106, R2358_U107, R2358_U108, R2358_U109, R2358_U110, R2358_U111, R2358_U112, R2358_U113, R2358_U114, R2358_U115, R2358_U116, R2358_U117, R2358_U118, R2358_U119, R2358_U120, R2358_U121, R2358_U122, R2358_U123, R2358_U124, R2358_U125, R2358_U126, R2358_U127, R2358_U128, R2358_U129, R2358_U130, R2358_U131, R2358_U132, R2358_U133, R2358_U134, R2358_U135, R2358_U136, R2358_U137, R2358_U138, R2358_U139, R2358_U140, R2358_U141, R2358_U142, R2358_U143, R2358_U144, R2358_U145, R2358_U146, R2358_U147, R2358_U148, R2358_U149, R2358_U150, R2358_U151, R2358_U152, R2358_U153, R2358_U154, R2358_U155, R2358_U156, R2358_U157, R2358_U158, R2358_U159, R2358_U160, R2358_U161, R2358_U162, R2358_U163, R2358_U164, R2358_U165, R2358_U166, R2358_U167, R2358_U168, R2358_U169, R2358_U170, R2358_U171, R2358_U172, R2358_U173, R2358_U174, R2358_U175, R2358_U176, R2358_U177, R2358_U178, R2358_U179, R2358_U180, R2358_U181, R2358_U182, R2358_U183, R2358_U184, R2358_U185, R2358_U186, R2358_U187, R2358_U188, R2358_U189, R2358_U190, R2358_U191, R2358_U192, R2358_U193, R2358_U194, R2358_U195, R2358_U196, R2358_U197, R2358_U198, R2358_U199, R2358_U200, R2358_U201, R2358_U202, R2358_U203, R2358_U204, R2358_U205, R2358_U206, R2358_U207, R2358_U208, R2358_U209, R2358_U210, R2358_U211, R2358_U212, R2358_U213, R2358_U214, R2358_U215, R2358_U216, R2358_U217, R2358_U218, R2358_U219, R2358_U220, R2358_U221, R2358_U222, R2358_U223, R2358_U224, R2358_U225, R2358_U226, R2358_U227, R2358_U228, R2358_U229, R2358_U230, R2358_U231, R2358_U232, R2358_U233, R2358_U234, R2358_U235, R2358_U236, R2358_U237, R2358_U238, R2358_U239, R2358_U240, R2358_U241, R2358_U242, R2358_U243, R2358_U244, R2358_U245, R2358_U246, R2358_U247, R2358_U248, R2358_U249, R2358_U250, R2358_U251, R2358_U252, R2358_U253, R2358_U254, R2358_U255, R2358_U256, R2358_U257, R2358_U258, R2358_U259, R2358_U260, R2358_U261, R2358_U262, R2358_U263, R2358_U264, R2358_U265, R2358_U266, R2358_U267, R2358_U268, R2358_U269, R2358_U270, R2358_U271, R2358_U272, R2358_U273, R2358_U274, R2358_U275, R2358_U276, R2358_U277, R2358_U278, R2358_U279, R2358_U280, R2358_U281, R2358_U282, R2358_U283, R2358_U284, R2358_U285, R2358_U286, R2358_U287, R2358_U288, R2358_U289, R2358_U290, R2358_U291, R2358_U292, R2358_U293, R2358_U294, R2358_U295, R2358_U296, R2358_U297, R2358_U298, R2358_U299, R2358_U300, R2358_U301, R2358_U302, R2358_U303, R2358_U304, R2358_U305, R2358_U306, R2358_U307, R2358_U308, R2358_U309, R2358_U310, R2358_U311, R2358_U312, R2358_U313, R2358_U314, R2358_U315, R2358_U316, R2358_U317, R2358_U318, R2358_U319, R2358_U320, R2358_U321, R2358_U322, R2358_U323, R2358_U324, R2358_U325, R2358_U326, R2358_U327, R2358_U328, R2358_U329, R2358_U330, R2358_U331, R2358_U332, R2358_U333, R2358_U334, R2358_U335, R2358_U336, R2358_U337, R2358_U338, R2358_U339, R2358_U340, R2358_U341, R2358_U342, R2358_U343, R2358_U344, R2358_U345, R2358_U346, R2358_U347, R2358_U348, R2358_U349, R2358_U350, R2358_U351, R2358_U352, R2358_U353, R2358_U354, R2358_U355, R2358_U356, R2358_U357, R2358_U358, R2358_U359, R2358_U360, R2358_U361, R2358_U362, R2358_U363, R2358_U364, R2358_U365, R2358_U366, R2358_U367, R2358_U368, R2358_U369, R2358_U370, R2358_U371, R2358_U372, R2358_U373, R2358_U374, R2358_U375, R2358_U376, R2358_U377, R2358_U378, R2358_U379, R2358_U380, R2358_U381, R2358_U382, R2358_U383, R2358_U384, R2358_U385, R2358_U386, R2358_U387, R2358_U388, R2358_U389, R2358_U390, R2358_U391, R2358_U392, R2358_U393, R2358_U394, R2358_U395, R2358_U396, R2358_U397, R2358_U398, R2358_U399, R2358_U400, R2358_U401, R2358_U402, R2358_U403, R2358_U404, R2358_U405, R2358_U406, R2358_U407, R2358_U408, R2358_U409, R2358_U410, R2358_U411, R2358_U412, R2358_U413, R2358_U414, R2358_U415, R2358_U416, R2358_U417, R2358_U418, R2358_U419, R2358_U420, R2358_U421, R2358_U422, R2358_U423, R2358_U424, R2358_U425, R2358_U426, R2358_U427, R2358_U428, R2358_U429, R2358_U430, R2358_U431, R2358_U432, R2358_U433, R2358_U434, R2358_U435, R2358_U436, R2358_U437, R2358_U438, R2358_U439, R2358_U440, R2358_U441, R2358_U442, R2358_U443, R2358_U444, R2358_U445, R2358_U446, R2358_U447, R2358_U448, R2358_U449, R2358_U450, R2358_U451, R2358_U452, R2358_U453, R2358_U454, R2358_U455, R2358_U456, R2358_U457, R2358_U458, R2358_U459, R2358_U460, R2358_U461, R2358_U462, R2358_U463, R2358_U464, R2358_U465, R2358_U466, R2358_U467, R2358_U468, R2358_U469, R2358_U470, R2358_U471, R2358_U472, R2358_U473, R2358_U474, R2358_U475, R2358_U476, R2358_U477, R2358_U478, R2358_U479, R2358_U480, R2358_U481, R2358_U482, R2358_U483, R2358_U484, R2358_U485, R2358_U486, R2358_U487, R2358_U488, R2358_U489, R2358_U490, R2358_U491, R2358_U492, R2358_U493, R2358_U494, R2358_U495, R2358_U496, R2358_U497, R2358_U498, R2358_U499, R2358_U500, R2358_U501, R2358_U502, R2358_U503, R2358_U504, R2358_U505, R2358_U506, R2358_U507, R2358_U508, R2358_U509, R2358_U510, R2358_U511, R2358_U512, R2358_U513, R2358_U514, R2358_U515, R2358_U516, R2358_U517, R2358_U518, R2358_U519, R2358_U520, R2358_U521, R2358_U522, R2358_U523, R2358_U524, R2358_U525, R2358_U526, R2358_U527, R2358_U528, R2358_U529, R2358_U530, R2358_U531, R2358_U532, R2358_U533, R2358_U534, R2358_U535, R2358_U536, R2358_U537, R2358_U538, R2358_U539, R2358_U540, R2358_U541, R2358_U542, R2358_U543, R2358_U544, R2358_U545, R2358_U546, R2358_U547, R2358_U548, R2358_U549, R2358_U550, R2358_U551, R2358_U552, R2358_U553, R2358_U554, R2358_U555, R2358_U556, R2358_U557, R2358_U558, R2358_U559, R2358_U560, R2358_U561, R2358_U562, R2358_U563, R2358_U564, R2358_U565, R2358_U566, R2358_U567, R2358_U568, R2358_U569, R2358_U570, R2358_U571, R2358_U572, R2358_U573, R2358_U574, R2358_U575, R2358_U576, R2358_U577, R2358_U578, R2358_U579, R2358_U580, R2358_U581, R2358_U582, R2358_U583, R2358_U584, R2358_U585, R2358_U586, R2358_U587, R2358_U588, R2358_U589, R2358_U590, R2358_U591, R2358_U592, R2358_U593, R2358_U594, R2358_U595, R2358_U596, R2358_U597, R2358_U598, R2358_U599, R2358_U600, R2358_U601, R2358_U602, R2358_U603, R2358_U604, R2358_U605, R2358_U606, R2358_U607, R2358_U608, R2358_U609, R2358_U610, R2358_U611, R2358_U612, R2358_U613, R2358_U614, R2358_U615, R2358_U616, R2358_U617, R2358_U618, R2358_U619, R2358_U620, R2358_U621, R2358_U622, R2358_U623, R2358_U624, R2358_U625, R2358_U626, R2358_U627, R2358_U628, R2358_U629, R2358_U630, R2358_U631, R2358_U632, R2358_U633, R2358_U634, R2358_U635, R2358_U636, R2358_U637, R2358_U638, R2358_U639, R2358_U640, R2358_U641, R2358_U642, R2358_U643, R2358_U644, R2358_U645, R2358_U646, R2358_U647, R2358_U648, R2358_U649, R2358_U650, R2358_U651, R2358_U652, R2358_U653, R2358_U654, R2337_U5, R2337_U6, R2337_U7, R2337_U8, R2337_U9, R2337_U10, R2337_U11, R2337_U12, R2337_U13, R2337_U14, R2337_U15, R2337_U16, R2337_U17, R2337_U18, R2337_U19, R2337_U20, R2337_U21, R2337_U22, R2337_U23, R2337_U24, R2337_U25, R2337_U26, R2337_U27, R2337_U28, R2337_U29, R2337_U30, R2337_U31, R2337_U32, R2337_U33, R2337_U34, R2337_U35, R2337_U36, R2337_U37, R2337_U38, R2337_U39, R2337_U40, R2337_U41, R2337_U42, R2337_U43, R2337_U44, R2337_U45, R2337_U46, R2337_U47, R2337_U48, R2337_U49, R2337_U50, R2337_U51, R2337_U52, R2337_U53, R2337_U54, R2337_U55, R2337_U56, R2337_U57, R2337_U58, R2337_U59, R2337_U60, R2337_U61, R2337_U62, R2337_U63, R2337_U64, R2337_U65, R2337_U66, R2337_U67, R2337_U68, R2337_U69, R2337_U70, R2337_U71, R2337_U72, R2337_U73, R2337_U74, R2337_U75, R2337_U76, R2337_U77, R2337_U78, R2337_U79, R2337_U80, R2337_U81, R2337_U82, R2337_U83, R2337_U84, R2337_U85, R2337_U86, R2337_U87, R2337_U88, R2337_U89, R2337_U90, R2337_U91, R2337_U92, R2337_U93, R2337_U94, R2337_U95, R2337_U96, R2337_U97, R2337_U98, R2337_U99, R2337_U100, R2337_U101, R2337_U102, R2337_U103, R2337_U104, R2337_U105, R2337_U106, R2337_U107, R2337_U108, R2337_U109, R2337_U110, R2337_U111, R2337_U112, R2337_U113, R2337_U114, R2337_U115, R2337_U116, R2337_U117, R2337_U118, R2337_U119, R2337_U120, R2337_U121, R2337_U122, R2337_U123, R2337_U124, R2337_U125, R2337_U126, R2337_U127, R2337_U128, R2337_U129, R2337_U130, R2337_U131, R2337_U132, R2337_U133, R2337_U134, R2337_U135, R2337_U136, R2337_U137, R2337_U138, R2337_U139, R2337_U140, R2337_U141, R2337_U142, R2337_U143, R2337_U144, R2337_U145, R2337_U146, R2337_U147, R2337_U148, R2337_U149, R2337_U150, R2337_U151, R2337_U152, R2337_U153, R2337_U154, R2337_U155, R2337_U156, R2337_U157, R2337_U158, R2337_U159, R2337_U160, R2337_U161, R2337_U162, R2337_U163, R2337_U164, R2337_U165, R2337_U166, R2337_U167, R2337_U168, R2337_U169, R2337_U170, R2337_U171, R2337_U172, R2337_U173, R2337_U174, R2337_U175, R2337_U176, R2337_U177, R2337_U178, R2337_U179, R2337_U180, R2337_U181, R2337_U182, R2337_U183, R2337_U184, R2337_U185, R2337_U186, R2337_U187, R2337_U188, R2337_U189, R2337_U190, R2337_U191, R2337_U192, R2337_U193, R2182_U5, R2182_U6, R2182_U7, R2182_U8, R2182_U9, R2182_U10, R2182_U11, R2182_U12, R2182_U13, R2182_U14, R2182_U15, R2182_U16, R2182_U17, R2182_U18, R2182_U19, R2182_U20, R2182_U21, R2182_U22, R2182_U23, R2182_U24, R2182_U25, R2182_U26, R2182_U27, R2182_U28, R2182_U29, R2182_U30, R2182_U31, R2182_U32, R2182_U33, R2182_U34, R2182_U35, R2182_U36, R2182_U37, R2182_U38, R2182_U39, R2182_U40, R2182_U41, R2182_U42, R2182_U43, R2182_U44, R2182_U45, R2182_U46, R2182_U47, R2182_U48, R2182_U49, R2182_U50, R2182_U51, R2182_U52, R2182_U53, R2182_U54, R2182_U55, R2182_U56, R2182_U57, R2182_U58, R2182_U59, R2182_U60, R2182_U61, R2182_U62, R2182_U63, R2182_U64, R2182_U65, R2182_U66, R2182_U67, R2182_U68, R2182_U69, R2182_U70, R2182_U71, R2182_U72, R2182_U73, R2182_U74, R2182_U75, R2182_U76, R2182_U77, R2182_U78, R2182_U79, R2182_U80, R2182_U81, R2182_U82, R2182_U83, R2182_U84, R2182_U85, R2182_U86, R2144_U5, R2144_U6, R2144_U7, R2144_U8, R2144_U9, R2144_U10, R2144_U11, R2144_U12, R2144_U13, R2144_U14, R2144_U15, R2144_U16, R2144_U17, R2144_U18, R2144_U19, R2144_U20, R2144_U21, R2144_U22, R2144_U23, R2144_U24, R2144_U25, R2144_U26, R2144_U27, R2144_U28, R2144_U29, R2144_U30, R2144_U31, R2144_U32, R2144_U33, R2144_U34, R2144_U35, R2144_U36, R2144_U37, R2144_U38, R2144_U39, R2144_U40, R2144_U41, R2144_U42, R2144_U43, R2144_U44, R2144_U45, R2144_U46, R2144_U47, R2144_U48, R2144_U49, R2144_U50, R2144_U51, R2144_U52, R2144_U53, R2144_U54, R2144_U55, R2144_U56, R2144_U57, R2144_U58, R2144_U59, R2144_U60, R2144_U61, R2144_U62, R2144_U63, R2144_U64, R2144_U65, R2144_U66, R2144_U67, R2144_U68, R2144_U69, R2144_U70, R2144_U71, R2144_U72, R2144_U73, R2144_U74, R2144_U75, R2144_U76, R2144_U77, R2144_U78, R2144_U79, R2144_U80, R2144_U81, R2144_U82, R2144_U83, R2144_U84, R2144_U85, R2144_U86, R2144_U87, R2144_U88, R2144_U89, R2144_U90, R2144_U91, R2144_U92, R2144_U93, R2144_U94, R2144_U95, R2144_U96, R2144_U97, R2144_U98, R2144_U99, R2144_U100, R2144_U101, R2144_U102, R2144_U103, R2144_U104, R2144_U105, R2144_U106, R2144_U107, R2144_U108, R2144_U109, R2144_U110, R2144_U111, R2144_U112, R2144_U113, R2144_U114, R2144_U115, R2144_U116, R2144_U117, R2144_U118, R2144_U119, R2144_U120, R2144_U121, R2144_U122, R2144_U123, R2144_U124, R2144_U125, R2144_U126, R2144_U127, R2144_U128, R2144_U129, R2144_U130, R2144_U131, R2144_U132, R2144_U133, R2144_U134, R2144_U135, R2144_U136, R2144_U137, R2144_U138, R2144_U139, R2144_U140, R2144_U141, R2144_U142, R2144_U143, R2144_U144, R2144_U145, R2144_U146, R2144_U147, R2144_U148, R2144_U149, R2144_U150, R2144_U151, R2144_U152, R2144_U153, R2144_U154, R2144_U155, R2144_U156, R2144_U157, R2144_U158, R2144_U159, R2144_U160, R2144_U161, R2144_U162, R2144_U163, R2144_U164, R2144_U165, R2144_U166, R2144_U167, R2144_U168, R2144_U169, R2144_U170, R2144_U171, R2144_U172, R2144_U173, R2144_U174, R2144_U175, R2144_U176, R2144_U177, R2144_U178, R2144_U179, R2144_U180, R2144_U181, R2144_U182, R2144_U183, R2144_U184, R2144_U185, R2144_U186, R2144_U187, R2144_U188, R2144_U189, R2144_U190, R2144_U191, R2144_U192, R2144_U193, R2144_U194, R2144_U195, R2144_U196, R2144_U197, R2144_U198, R2144_U199, R2144_U200, R2144_U201, R2144_U202, R2144_U203, R2144_U204, R2144_U205, R2144_U206, R2144_U207, R2144_U208, R2144_U209, R2144_U210, R2144_U211, R2144_U212, R2144_U213, R2144_U214, R2144_U215, R2144_U216, R2144_U217, R2144_U218, R2144_U219, R2144_U220, R2144_U221, R2144_U222, R2144_U223, R2144_U224, R2144_U225, R2144_U226, R2144_U227, R2144_U228, R2144_U229, R2144_U230, R2144_U231, R2144_U232, R2144_U233, R2144_U234, R2144_U235, R2144_U236, R2144_U237, R2144_U238, R2144_U239, R2144_U240, R2144_U241, R2144_U242, R2144_U243, R2144_U244, R2144_U245, R2144_U246, R2144_U247, R2144_U248, R2144_U249, R2144_U250, R2144_U251, R2144_U252, R2144_U253, R2144_U254, R2144_U255, R2144_U256, R2144_U257, R2144_U258, R2144_U259, R2144_U260, LT_589_U6, LT_589_U7, LT_589_U8, R584_U6, R584_U7, R584_U8, R584_U9, R2099_U4, R2099_U5, R2099_U6, R2099_U7, R2099_U8, R2099_U9, R2099_U10, R2099_U11, R2099_U12, R2099_U13, R2099_U14, R2099_U15, R2099_U16, R2099_U17, R2099_U18, R2099_U19, R2099_U20, R2099_U21, R2099_U22, R2099_U23, R2099_U24, R2099_U25, R2099_U26, R2099_U27, R2099_U28, R2099_U29, R2099_U30, R2099_U31, R2099_U32, R2099_U33, R2099_U34, R2099_U35, R2099_U36, R2099_U37, R2099_U38, R2099_U39, R2099_U40, R2099_U41, R2099_U42, R2099_U43, R2099_U44, R2099_U45, R2099_U46, R2099_U47, R2099_U48, R2099_U49, R2099_U50, R2099_U51, R2099_U52, R2099_U53, R2099_U54, R2099_U55, R2099_U56, R2099_U57, R2099_U58, R2099_U59, R2099_U60, R2099_U61, R2099_U62, R2099_U63, R2099_U64, R2099_U65, R2099_U66, R2099_U67, R2099_U68, R2099_U69, R2099_U70, R2099_U71, R2099_U72, R2099_U73, R2099_U74, R2099_U75, R2099_U76, R2099_U77, R2099_U78, R2099_U79, R2099_U80, R2099_U81, R2099_U82, R2099_U83, R2099_U84, R2099_U85, R2099_U86, R2099_U87, R2099_U88, R2099_U89, R2099_U90, R2099_U91, R2099_U92, R2099_U93, R2099_U94, R2099_U95, R2099_U96, R2099_U97, R2099_U98, R2099_U99, R2099_U100, R2099_U101, R2099_U102, R2099_U103, R2099_U104, R2099_U105, R2099_U106, R2099_U107, R2099_U108, R2099_U109, R2099_U110, R2099_U111, R2099_U112, R2099_U113, R2099_U114, R2099_U115, R2099_U116, R2099_U117, R2099_U118, R2099_U119, R2099_U120, R2099_U121, R2099_U122, R2099_U123, R2099_U124, R2099_U125, R2099_U126, R2099_U127, R2099_U128, R2099_U129, R2099_U130, R2099_U131, R2099_U132, R2099_U133, R2099_U134, R2099_U135, R2099_U136, R2099_U137, R2099_U138, R2099_U139, R2099_U140, R2099_U141, R2099_U142, R2099_U143, R2099_U144, R2099_U145, R2099_U146, R2099_U147, R2099_U148, R2099_U149, R2099_U150, R2099_U151, R2099_U152, R2099_U153, R2099_U154, R2099_U155, R2099_U156, R2099_U157, R2099_U158, R2099_U159, R2099_U160, R2099_U161, R2099_U162, R2099_U163, R2099_U164, R2099_U165, R2099_U166, R2099_U167, R2099_U168, R2099_U169, R2099_U170, R2099_U171, R2099_U172, R2099_U173, R2099_U174, R2099_U175, R2099_U176, R2099_U177, R2099_U178, R2099_U179, R2099_U180, R2099_U181, R2099_U182, R2099_U183, R2099_U184, R2099_U185, R2099_U186, R2099_U187, R2099_U188, R2099_U189, R2099_U190, R2099_U191, R2099_U192, R2099_U193, R2099_U194, R2099_U195, R2099_U196, R2099_U197, R2099_U198, R2099_U199, R2099_U200, R2099_U201, R2099_U202, R2099_U203, R2099_U204, R2099_U205, R2099_U206, R2099_U207, R2099_U208, R2099_U209, R2099_U210, R2099_U211, R2099_U212, R2099_U213, R2099_U214, R2099_U215, R2099_U216, R2099_U217, R2099_U218, R2099_U219, R2099_U220, R2099_U221, R2099_U222, R2099_U223, R2099_U224, R2099_U225, R2099_U226, R2099_U227, R2099_U228, R2099_U229, R2099_U230, R2099_U231, R2099_U232, R2099_U233, R2099_U234, R2099_U235, R2099_U236, R2099_U237, R2099_U238, R2099_U239, R2099_U240, R2099_U241, R2099_U242, R2099_U243, R2099_U244, R2099_U245, R2099_U246, R2099_U247, R2099_U248, R2099_U249, R2099_U250, R2099_U251, R2099_U252, R2099_U253, R2099_U254, R2099_U255, R2099_U256, R2099_U257, R2099_U258, R2099_U259, R2099_U260, R2099_U261, R2099_U262, R2099_U263, R2099_U264, R2099_U265, R2099_U266, R2099_U267, R2099_U268, R2099_U269, R2099_U270, R2099_U271, R2099_U272, R2099_U273, R2099_U274, R2099_U275, R2099_U276, R2099_U277, R2099_U278, R2099_U279, R2099_U280, R2099_U281, R2099_U282, R2099_U283, R2099_U284, R2099_U285, R2099_U286, R2099_U287, R2099_U288, R2099_U289, R2099_U290, R2099_U291, R2099_U292, R2099_U293, R2099_U294, R2099_U295, R2099_U296, R2099_U297, R2099_U298, R2099_U299, R2099_U300, R2099_U301, R2099_U302, R2099_U303, R2099_U304, R2099_U305, R2099_U306, R2099_U307, R2099_U308, R2099_U309, R2099_U310, R2099_U311, R2099_U312, R2099_U313, R2099_U314, R2099_U315, R2099_U316, R2099_U317, R2099_U318, R2099_U319, R2099_U320, R2099_U321, R2099_U322, R2099_U323, R2099_U324, R2099_U325, R2099_U326, R2099_U327, R2099_U328, R2099_U329, R2099_U330, R2099_U331, R2099_U332, R2099_U333, R2099_U334, R2099_U335, R2099_U336, R2099_U337, R2099_U338, R2099_U339, R2099_U340, R2099_U341, R2099_U342, R2099_U343, R2099_U344, R2099_U345, R2099_U346, R2099_U347, R2099_U348, R2099_U349, R2167_U6, R2167_U7, R2167_U8, R2167_U9, R2167_U10, R2167_U11, R2167_U12, R2167_U13, R2167_U14, R2167_U15, R2167_U16, R2167_U17, R2167_U18, R2167_U19, R2167_U20, R2167_U21, R2167_U22, R2167_U23, R2167_U24, R2167_U25, R2167_U26, R2167_U27, R2167_U28, R2167_U29, R2167_U30, R2167_U31, R2167_U32, R2167_U33, R2167_U34, R2167_U35, R2167_U36, R2167_U37, R2167_U38, R2167_U39, R2167_U40, R2167_U41, R2167_U42, R2167_U43, R2167_U44, R2167_U45, R2167_U46, R2167_U47, R2167_U48, R2167_U49, R2167_U50, SUB_357_U6, SUB_357_U7, SUB_357_U8, SUB_357_U9, SUB_357_U10, SUB_357_U11, SUB_357_U12, SUB_357_U13, LT_563_1260_U6, LT_563_1260_U7, LT_563_1260_U8, LT_563_1260_U9, SUB_580_U6, SUB_580_U7, SUB_580_U8, SUB_580_U9, SUB_580_U10, R2096_U4, R2096_U5, R2096_U6, R2096_U7, R2096_U8, R2096_U9, R2096_U10, R2096_U11, R2096_U12, R2096_U13, R2096_U14, R2096_U15, R2096_U16, R2096_U17, R2096_U18, R2096_U19, R2096_U20, R2096_U21, R2096_U22, R2096_U23, R2096_U24, R2096_U25, R2096_U26, R2096_U27, R2096_U28, R2096_U29, R2096_U30, R2096_U31, R2096_U32, R2096_U33, R2096_U34, R2096_U35, R2096_U36, R2096_U37, R2096_U38, R2096_U39, R2096_U40, R2096_U41, R2096_U42, R2096_U43, R2096_U44, R2096_U45, R2096_U46, R2096_U47, R2096_U48, R2096_U49, R2096_U50, R2096_U51, R2096_U52, R2096_U53, R2096_U54, R2096_U55, R2096_U56, R2096_U57, R2096_U58, R2096_U59, R2096_U60, R2096_U61, R2096_U62, R2096_U63, R2096_U64, R2096_U65, R2096_U66, R2096_U67, R2096_U68, R2096_U69, R2096_U70, R2096_U71, R2096_U72, R2096_U73, R2096_U74, R2096_U75, R2096_U76, R2096_U77, R2096_U78, R2096_U79, R2096_U80, R2096_U81, R2096_U82, R2096_U83, R2096_U84, R2096_U85, R2096_U86, R2096_U87, R2096_U88, R2096_U89, R2096_U90, R2096_U91, R2096_U92, R2096_U93, R2096_U94, R2096_U95, R2096_U96, R2096_U97, R2096_U98, R2096_U99, R2096_U100, R2096_U101, R2096_U102, R2096_U103, R2096_U104, R2096_U105, R2096_U106, R2096_U107, R2096_U108, R2096_U109, R2096_U110, R2096_U111, R2096_U112, R2096_U113, R2096_U114, R2096_U115, R2096_U116, R2096_U117, R2096_U118, R2096_U119, R2096_U120, R2096_U121, R2096_U122, R2096_U123, R2096_U124, R2096_U125, R2096_U126, R2096_U127, R2096_U128, R2096_U129, R2096_U130, R2096_U131, R2096_U132, R2096_U133, R2096_U134, R2096_U135, R2096_U136, R2096_U137, R2096_U138, R2096_U139, R2096_U140, R2096_U141, R2096_U142, R2096_U143, R2096_U144, R2096_U145, R2096_U146, R2096_U147, R2096_U148, R2096_U149, R2096_U150, R2096_U151, R2096_U152, R2096_U153, R2096_U154, R2096_U155, R2096_U156, R2096_U157, R2096_U158, R2096_U159, R2096_U160, R2096_U161, R2096_U162, R2096_U163, R2096_U164, R2096_U165, R2096_U166, R2096_U167, R2096_U168, R2096_U169, R2096_U170, R2096_U171, R2096_U172, R2096_U173, R2096_U174, R2096_U175, R2096_U176, R2096_U177, R2096_U178, R2096_U179, R2096_U180, R2096_U181, R2096_U182, LT_563_U6, LT_563_U7, LT_563_U8, LT_563_U9, LT_563_U10, LT_563_U11, LT_563_U12, LT_563_U13, LT_563_U14, LT_563_U15, LT_563_U16, LT_563_U17, LT_563_U18, LT_563_U19, LT_563_U20, LT_563_U21, LT_563_U22, LT_563_U23, LT_563_U24, LT_563_U25, LT_563_U26, LT_563_U27, LT_563_U28, R2238_U6, R2238_U7, R2238_U8, R2238_U9, R2238_U10, R2238_U11, R2238_U12, R2238_U13, R2238_U14, R2238_U15, R2238_U16, R2238_U17, R2238_U18, R2238_U19, R2238_U20, R2238_U21, R2238_U22, R2238_U23, R2238_U24, R2238_U25, R2238_U26, R2238_U27, R2238_U28, R2238_U29, R2238_U30, R2238_U31, R2238_U32, R2238_U33, R2238_U34, R2238_U35, R2238_U36, R2238_U37, R2238_U38, R2238_U39, R2238_U40, R2238_U41, R2238_U42, R2238_U43, R2238_U44, R2238_U45, R2238_U46, R2238_U47, R2238_U48, R2238_U49, R2238_U50, R2238_U51, R2238_U52, R2238_U53, R2238_U54, R2238_U55, R2238_U56, R2238_U57, R2238_U58, R2238_U59, R2238_U60, R2238_U61, R2238_U62, R2238_U63, R2238_U64, R2238_U65, R2238_U66, SUB_450_U6, SUB_450_U7, SUB_450_U8, SUB_450_U9, SUB_450_U10, SUB_450_U11, SUB_450_U12, SUB_450_U13, SUB_450_U14, SUB_450_U15, SUB_450_U16, SUB_450_U17, SUB_450_U18, SUB_450_U19, SUB_450_U20, SUB_450_U21, SUB_450_U22, SUB_450_U23, SUB_450_U24, SUB_450_U25, SUB_450_U26, SUB_450_U27, SUB_450_U28, SUB_450_U29, SUB_450_U30, SUB_450_U31, SUB_450_U32, SUB_450_U33, SUB_450_U34, SUB_450_U35, SUB_450_U36, SUB_450_U37, SUB_450_U38, SUB_450_U39, SUB_450_U40, SUB_450_U41, SUB_450_U42, SUB_450_U43, SUB_450_U44, SUB_450_U45, SUB_450_U46, SUB_450_U47, SUB_450_U48, SUB_450_U49, SUB_450_U50, SUB_450_U51, SUB_450_U52, SUB_450_U53, SUB_450_U54, SUB_450_U55, SUB_450_U56, SUB_450_U57, SUB_450_U58, SUB_450_U59, SUB_450_U60, SUB_450_U61, SUB_450_U62, SUB_450_U63, SUB_450_U64, SUB_450_U65, SUB_450_U66, ADD_371_U4, ADD_371_U5, ADD_371_U6, ADD_371_U7, ADD_371_U8, ADD_371_U9, ADD_371_U10, ADD_371_U11, ADD_371_U12, ADD_371_U13, ADD_371_U14, ADD_371_U15, ADD_371_U16, ADD_371_U17, ADD_371_U18, ADD_371_U19, ADD_371_U20, ADD_371_U21, ADD_371_U22, ADD_371_U23, ADD_371_U24, ADD_371_U25, ADD_371_U26, ADD_371_U27, ADD_371_U28, ADD_371_U29, ADD_371_U30, ADD_371_U31, ADD_371_U32, ADD_371_U33, ADD_371_U34, ADD_371_U35, ADD_371_U36, ADD_371_U37, ADD_371_U38, ADD_371_U39, ADD_371_U40, ADD_371_U41, ADD_371_U42, ADD_371_U43, ADD_371_U44, ADD_405_U4, ADD_405_U5, ADD_405_U6, ADD_405_U7, ADD_405_U8, ADD_405_U9, ADD_405_U10, ADD_405_U11, ADD_405_U12, ADD_405_U13, ADD_405_U14, ADD_405_U15, ADD_405_U16, ADD_405_U17, ADD_405_U18, ADD_405_U19, ADD_405_U20, ADD_405_U21, ADD_405_U22, ADD_405_U23, ADD_405_U24, ADD_405_U25, ADD_405_U26, ADD_405_U27, ADD_405_U28, ADD_405_U29, ADD_405_U30, ADD_405_U31, ADD_405_U32, ADD_405_U33, ADD_405_U34, ADD_405_U35, ADD_405_U36, ADD_405_U37, ADD_405_U38, ADD_405_U39, ADD_405_U40, ADD_405_U41, ADD_405_U42, ADD_405_U43, ADD_405_U44, ADD_405_U45, ADD_405_U46, ADD_405_U47, ADD_405_U48, ADD_405_U49, ADD_405_U50, ADD_405_U51, ADD_405_U52, ADD_405_U53, ADD_405_U54, ADD_405_U55, ADD_405_U56, ADD_405_U57, ADD_405_U58, ADD_405_U59, ADD_405_U60, ADD_405_U61, ADD_405_U62, ADD_405_U63, ADD_405_U64, ADD_405_U65, ADD_405_U66, ADD_405_U67, ADD_405_U68, ADD_405_U69, ADD_405_U70, ADD_405_U71, ADD_405_U72, ADD_405_U73, ADD_405_U74, ADD_405_U75, ADD_405_U76, ADD_405_U77, ADD_405_U78, ADD_405_U79, ADD_405_U80, ADD_405_U81, ADD_405_U82, ADD_405_U83, ADD_405_U84, ADD_405_U85, ADD_405_U86, ADD_405_U87, ADD_405_U88, ADD_405_U89, ADD_405_U90, ADD_405_U91, ADD_405_U92, ADD_405_U93, ADD_405_U94, ADD_405_U95, ADD_405_U96, ADD_405_U97, ADD_405_U98, ADD_405_U99, ADD_405_U100, ADD_405_U101, ADD_405_U102, ADD_405_U103, ADD_405_U104, ADD_405_U105, ADD_405_U106, ADD_405_U107, ADD_405_U108, ADD_405_U109, ADD_405_U110, ADD_405_U111, ADD_405_U112, ADD_405_U113, ADD_405_U114, ADD_405_U115, ADD_405_U116, ADD_405_U117, ADD_405_U118, ADD_405_U119, ADD_405_U120, ADD_405_U121, ADD_405_U122, ADD_405_U123, ADD_405_U124, ADD_405_U125, ADD_405_U126, ADD_405_U127, ADD_405_U128, ADD_405_U129, ADD_405_U130, ADD_405_U131, ADD_405_U132, ADD_405_U133, ADD_405_U134, ADD_405_U135, ADD_405_U136, ADD_405_U137, ADD_405_U138, ADD_405_U139, ADD_405_U140, ADD_405_U141, ADD_405_U142, ADD_405_U143, ADD_405_U144, ADD_405_U145, ADD_405_U146, ADD_405_U147, ADD_405_U148, ADD_405_U149, ADD_405_U150, ADD_405_U151, ADD_405_U152, ADD_405_U153, ADD_405_U154, ADD_405_U155, ADD_405_U156, ADD_405_U157, ADD_405_U158, ADD_405_U159, ADD_405_U160, ADD_405_U161, ADD_405_U162, ADD_405_U163, ADD_405_U164, ADD_405_U165, ADD_405_U166, ADD_405_U167, ADD_405_U168, ADD_405_U169, ADD_405_U170, ADD_405_U171, ADD_405_U172, ADD_405_U173, ADD_405_U174, ADD_405_U175, ADD_405_U176, ADD_405_U177, ADD_405_U178, ADD_405_U179, ADD_405_U180, ADD_405_U181, ADD_405_U182, ADD_405_U183, ADD_405_U184, ADD_405_U185, ADD_405_U186, GTE_485_U6, GTE_485_U7, ADD_515_U4, ADD_515_U5, ADD_515_U6, ADD_515_U7, ADD_515_U8, ADD_515_U9, ADD_515_U10, ADD_515_U11, ADD_515_U12, ADD_515_U13, ADD_515_U14, ADD_515_U15, ADD_515_U16, ADD_515_U17, ADD_515_U18, ADD_515_U19, ADD_515_U20, ADD_515_U21, ADD_515_U22, ADD_515_U23, ADD_515_U24, ADD_515_U25, ADD_515_U26, ADD_515_U27, ADD_515_U28, ADD_515_U29, ADD_515_U30, ADD_515_U31, ADD_515_U32, ADD_515_U33, ADD_515_U34, ADD_515_U35, ADD_515_U36, ADD_515_U37, ADD_515_U38, ADD_515_U39, ADD_515_U40, ADD_515_U41, ADD_515_U42, ADD_515_U43, ADD_515_U44, ADD_515_U45, ADD_515_U46, ADD_515_U47, ADD_515_U48, ADD_515_U49, ADD_515_U50, ADD_515_U51, ADD_515_U52, ADD_515_U53, ADD_515_U54, ADD_515_U55, ADD_515_U56, ADD_515_U57, ADD_515_U58, ADD_515_U59, ADD_515_U60, ADD_515_U61, ADD_515_U62, ADD_515_U63, ADD_515_U64, ADD_515_U65, ADD_515_U66, ADD_515_U67, ADD_515_U68, ADD_515_U69, ADD_515_U70, ADD_515_U71, ADD_515_U72, ADD_515_U73, ADD_515_U74, ADD_515_U75, ADD_515_U76, ADD_515_U77, ADD_515_U78, ADD_515_U79, ADD_515_U80, ADD_515_U81, ADD_515_U82, ADD_515_U83, ADD_515_U84, ADD_515_U85, ADD_515_U86, ADD_515_U87, ADD_515_U88, ADD_515_U89, ADD_515_U90, ADD_515_U91, ADD_515_U92, ADD_515_U93, ADD_515_U94, ADD_515_U95, ADD_515_U96, ADD_515_U97, ADD_515_U98, ADD_515_U99, ADD_515_U100, ADD_515_U101, ADD_515_U102, ADD_515_U103, ADD_515_U104, ADD_515_U105, ADD_515_U106, ADD_515_U107, ADD_515_U108, ADD_515_U109, ADD_515_U110, ADD_515_U111, ADD_515_U112, ADD_515_U113, ADD_515_U114, ADD_515_U115, ADD_515_U116, ADD_515_U117, ADD_515_U118, ADD_515_U119, ADD_515_U120, ADD_515_U121, ADD_515_U122, ADD_515_U123, ADD_515_U124, ADD_515_U125, ADD_515_U126, ADD_515_U127, ADD_515_U128, ADD_515_U129, ADD_515_U130, ADD_515_U131, ADD_515_U132, ADD_515_U133, ADD_515_U134, ADD_515_U135, ADD_515_U136, ADD_515_U137, ADD_515_U138, ADD_515_U139, ADD_515_U140, ADD_515_U141, ADD_515_U142, ADD_515_U143, ADD_515_U144, ADD_515_U145, ADD_515_U146, ADD_515_U147, ADD_515_U148, ADD_515_U149, ADD_515_U150, ADD_515_U151, ADD_515_U152, ADD_515_U153, ADD_515_U154, ADD_515_U155, ADD_515_U156, ADD_515_U157, ADD_515_U158, ADD_515_U159, ADD_515_U160, ADD_515_U161, ADD_515_U162, ADD_515_U163, ADD_515_U164, ADD_515_U165, ADD_515_U166, ADD_515_U167, ADD_515_U168, ADD_515_U169, ADD_515_U170, ADD_515_U171, ADD_515_U172, ADD_515_U173, ADD_515_U174, ADD_515_U175, ADD_515_U176, ADD_515_U177, ADD_515_U178, ADD_515_U179, ADD_515_U180, ADD_515_U181, ADD_515_U182; 
assign U2352 = ~(STATE2_REG_2__SCAN_IN | STATEBS16_REG_SCAN_IN); 
assign U2427 = ~(STATE2_REG_3__SCAN_IN | STATE2_REG_1__SCAN_IN); 
assign U2428 = STATE2_REG_2__SCAN_IN & STATE2_REG_1__SCAN_IN; 
assign U2453 = INSTQUEUERD_ADDR_REG_3__SCAN_IN & INSTQUEUERD_ADDR_REG_2__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign U2469 = ~(INSTQUEUERD_ADDR_REG_3__SCAN_IN | INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign U2478 = INSTQUEUEWR_ADDR_REG_3__SCAN_IN & INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign U2488 = ~(INSTQUEUEWR_ADDR_REG_1__SCAN_IN | INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign U2510 = ~(INSTQUEUEWR_ADDR_REG_3__SCAN_IN | INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign U3234 = ~REQUESTPENDING_REG_SCAN_IN; 
assign U3235 = ~STATE_REG_1__SCAN_IN; 
assign U3238 = ~STATE_REG_2__SCAN_IN; 
assign U3240 = ~REIP_REG_1__SCAN_IN; 
assign U3242 = STATE_REG_2__SCAN_IN | STATE_REG_1__SCAN_IN; 
assign U3243 = ~HOLD; 
assign U3244 = ~READY_N; 
assign U3245 = ~STATE_REG_0__SCAN_IN; 
assign U3248 = HOLD | REQUESTPENDING_REG_SCAN_IN; 
assign U3249 = ~STATE2_REG_1__SCAN_IN; 
assign U3250 = ~STATE2_REG_2__SCAN_IN; 
assign U3251 = ~INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign U3252 = ~INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign U3253 = ~INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign U3255 = INSTQUEUERD_ADDR_REG_2__SCAN_IN | INSTQUEUERD_ADDR_REG_1__SCAN_IN | INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign U3256 = INSTQUEUERD_ADDR_REG_1__SCAN_IN | INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign U3257 = ~INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign U3262 = ~(INSTQUEUERD_ADDR_REG_1__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U3267 = READY_N | STATEBS16_REG_SCAN_IN; 
assign U3281 = ~STATE2_REG_0__SCAN_IN; 
assign U3283 = ~STATE2_REG_3__SCAN_IN; 
assign U3285 = STATE2_REG_2__SCAN_IN | STATE2_REG_1__SCAN_IN; 
assign U3288 = ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN; 
assign U3289 = ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign U3290 = ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign U3291 = ~INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign U3292 = ~(INSTQUEUEWR_ADDR_REG_1__SCAN_IN & INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign U3294 = STATE2_REG_3__SCAN_IN | STATE2_REG_2__SCAN_IN; 
assign U3295 = ~STATEBS16_REG_SCAN_IN; 
assign U3374 = ~FLUSH_REG_SCAN_IN; 
assign U3400 = ~REIP_REG_0__SCAN_IN; 
assign U3416 = ~EBX_REG_31__SCAN_IN; 
assign U3422 = ~CODEFETCH_REG_SCAN_IN; 
assign U3423 = ~READREQUEST_REG_SCAN_IN; 
assign U3467 = ~(DATAWIDTH_REG_1__SCAN_IN | REIP_REG_1__SCAN_IN); 
assign U3481 = READY_N & STATE_REG_1__SCAN_IN; 
assign U3484 = STATE_REG_0__SCAN_IN & REQUESTPENDING_REG_SCAN_IN; 
assign U3485 = ~(INSTQUEUERD_ADDR_REG_3__SCAN_IN | INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign U3486 = INSTQUEUERD_ADDR_REG_1__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign U3487 = ~(INSTQUEUERD_ADDR_REG_3__SCAN_IN | INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U3488 = INSTQUEUERD_ADDR_REG_2__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign U3489 = ~(INSTQUEUERD_ADDR_REG_3__SCAN_IN | INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U3490 = INSTQUEUERD_ADDR_REG_2__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign U3491 = ~(INSTQUEUERD_ADDR_REG_2__SCAN_IN | INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U3492 = INSTQUEUERD_ADDR_REG_3__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign U3493 = ~(INSTQUEUERD_ADDR_REG_2__SCAN_IN | INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U3494 = INSTQUEUERD_ADDR_REG_3__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign U3495 = INSTQUEUERD_ADDR_REG_3__SCAN_IN & INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign U3508 = ~(INSTQUEUERD_ADDR_REG_3__SCAN_IN | INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U3509 = INSTQUEUE_REG_5__5__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign U3510 = ~(INSTQUEUERD_ADDR_REG_3__SCAN_IN | INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U3511 = INSTQUEUE_REG_6__5__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign U3512 = INSTQUEUE_REG_8__5__SCAN_IN & INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign U3513 = ~(INSTQUEUERD_ADDR_REG_2__SCAN_IN | INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U3514 = INSTQUEUE_REG_10__5__SCAN_IN & INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign U3515 = INSTQUEUE_REG_12__5__SCAN_IN & INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign U3516 = ~(INSTQUEUERD_ADDR_REG_2__SCAN_IN | INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U3517 = INSTQUEUE_REG_9__5__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign U3522 = ~(INSTQUEUERD_ADDR_REG_3__SCAN_IN | INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign U3523 = INSTQUEUE_REG_3__6__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign U3528 = ~(INSTQUEUERD_ADDR_REG_3__SCAN_IN | INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign U3529 = INSTQUEUE_REG_1__4__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign U3530 = ~(INSTQUEUERD_ADDR_REG_1__SCAN_IN | INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U3531 = INSTQUEUE_REG_4__4__SCAN_IN & INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign U3532 = ~(INSTQUEUERD_ADDR_REG_1__SCAN_IN | INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U3533 = INSTQUEUE_REG_12__4__SCAN_IN & INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign U3534 = INSTQUEUERD_ADDR_REG_2__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign U3535 = INSTQUEUE_REG_13__4__SCAN_IN & INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign U3536 = ~(INSTQUEUERD_ADDR_REG_3__SCAN_IN | INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U3537 = INSTQUEUE_REG_6__4__SCAN_IN & INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign U3538 = INSTQUEUERD_ADDR_REG_2__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign U3539 = INSTQUEUE_REG_14__4__SCAN_IN & INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign U3540 = ~(INSTQUEUERD_ADDR_REG_2__SCAN_IN | INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U3541 = INSTQUEUE_REG_9__4__SCAN_IN & INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign U3572 = STATE2_REG_3__SCAN_IN & STATE2_REG_0__SCAN_IN; 
assign U3719 = STATE2_REG_0__SCAN_IN & FLUSH_REG_SCAN_IN; 
assign U3852 = STATE2_REG_1__SCAN_IN & STATEBS16_REG_SCAN_IN; 
assign U3876 = ~(READY_N | STATEBS16_REG_SCAN_IN); 
assign U3938 = ~(DATAWIDTH_REG_2__SCAN_IN | DATAWIDTH_REG_3__SCAN_IN | DATAWIDTH_REG_4__SCAN_IN | DATAWIDTH_REG_5__SCAN_IN); 
assign U3939 = ~(DATAWIDTH_REG_6__SCAN_IN | DATAWIDTH_REG_7__SCAN_IN | DATAWIDTH_REG_8__SCAN_IN | DATAWIDTH_REG_9__SCAN_IN); 
assign U3941 = ~(DATAWIDTH_REG_10__SCAN_IN | DATAWIDTH_REG_11__SCAN_IN | DATAWIDTH_REG_12__SCAN_IN | DATAWIDTH_REG_13__SCAN_IN); 
assign U3942 = ~(DATAWIDTH_REG_14__SCAN_IN | DATAWIDTH_REG_15__SCAN_IN | DATAWIDTH_REG_16__SCAN_IN | DATAWIDTH_REG_17__SCAN_IN); 
assign U3944 = ~(DATAWIDTH_REG_18__SCAN_IN | DATAWIDTH_REG_19__SCAN_IN | DATAWIDTH_REG_20__SCAN_IN | DATAWIDTH_REG_21__SCAN_IN); 
assign U3945 = ~(DATAWIDTH_REG_22__SCAN_IN | DATAWIDTH_REG_23__SCAN_IN | DATAWIDTH_REG_24__SCAN_IN | DATAWIDTH_REG_25__SCAN_IN); 
assign U3947 = ~(DATAWIDTH_REG_26__SCAN_IN | DATAWIDTH_REG_27__SCAN_IN); 
assign U3948 = ~(DATAWIDTH_REG_28__SCAN_IN | DATAWIDTH_REG_29__SCAN_IN); 
assign U3949 = ~(DATAWIDTH_REG_30__SCAN_IN | DATAWIDTH_REG_31__SCAN_IN); 
assign U3951 = ~(DATAWIDTH_REG_0__SCAN_IN | DATAWIDTH_REG_1__SCAN_IN | REIP_REG_0__SCAN_IN); 
assign U3954 = ~(READY_N | STATE2_REG_0__SCAN_IN); 
assign U4162 = ~INSTADDRPOINTER_REG_31__SCAN_IN; 
assign U4167 = ~BS16_N; 
assign U4350 = NA_N | STATE_REG_0__SCAN_IN; 
assign U4402 = ~(INSTQUEUE_REG_15__5__SCAN_IN & INSTQUEUERD_ADDR_REG_3__SCAN_IN & INSTQUEUERD_ADDR_REG_2__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U4498 = FLUSH_REG_SCAN_IN | MORE_REG_SCAN_IN; 
assign U4501 = ~(READY_N & STATE2_REG_1__SCAN_IN); 
assign U5465 = ~(INSTQUEUERD_ADDR_REG_2__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U6355 = READY_N | STATEBS16_REG_SCAN_IN; 
assign U6586 = ~(DATAWIDTH_REG_0__SCAN_IN & DATAWIDTH_REG_1__SCAN_IN); 
assign U6587 = REIP_REG_0__SCAN_IN | REIP_REG_1__SCAN_IN; 
assign U6601 = ~(STATE_REG_0__SCAN_IN & ADS_N_REG_SCAN_IN); 
assign U7457 = READY_N | STATE2_REG_2__SCAN_IN; 
assign U7636 = STATE_REG_1__SCAN_IN | STATE_REG_0__SCAN_IN; 
assign U7652 = ~(INSTQUEUE_REG_15__4__SCAN_IN & INSTQUEUERD_ADDR_REG_3__SCAN_IN & INSTQUEUERD_ADDR_REG_2__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U7675 = STATE2_REG_0__SCAN_IN | STATEBS16_REG_SCAN_IN; 
assign U7702 = ~(INSTADDRPOINTER_REG_0__SCAN_IN & INSTADDRPOINTER_REG_31__SCAN_IN); 
assign U7736 = DATAWIDTH_REG_0__SCAN_IN | DATAWIDTH_REG_1__SCAN_IN; 
assign U7740 = ~(REIP_REG_0__SCAN_IN & REIP_REG_1__SCAN_IN); 
assign R2027_U5 = ~INSTADDRPOINTER_REG_0__SCAN_IN; 
assign R2027_U6 = ~INSTADDRPOINTER_REG_2__SCAN_IN; 
assign R2027_U7 = ~INSTADDRPOINTER_REG_1__SCAN_IN; 
assign R2027_U8 = ~INSTADDRPOINTER_REG_4__SCAN_IN; 
assign R2027_U9 = ~INSTADDRPOINTER_REG_3__SCAN_IN; 
assign R2027_U10 = ~(INSTADDRPOINTER_REG_0__SCAN_IN & INSTADDRPOINTER_REG_1__SCAN_IN & INSTADDRPOINTER_REG_2__SCAN_IN); 
assign R2027_U11 = ~INSTADDRPOINTER_REG_6__SCAN_IN; 
assign R2027_U12 = ~INSTADDRPOINTER_REG_5__SCAN_IN; 
assign R2027_U14 = ~INSTADDRPOINTER_REG_8__SCAN_IN; 
assign R2027_U15 = ~INSTADDRPOINTER_REG_7__SCAN_IN; 
assign R2027_U18 = ~INSTADDRPOINTER_REG_9__SCAN_IN; 
assign R2027_U19 = ~INSTADDRPOINTER_REG_10__SCAN_IN; 
assign R2027_U20 = ~INSTADDRPOINTER_REG_12__SCAN_IN; 
assign R2027_U21 = ~INSTADDRPOINTER_REG_11__SCAN_IN; 
assign R2027_U23 = ~INSTADDRPOINTER_REG_14__SCAN_IN; 
assign R2027_U24 = ~INSTADDRPOINTER_REG_13__SCAN_IN; 
assign R2027_U26 = ~INSTADDRPOINTER_REG_15__SCAN_IN; 
assign R2027_U28 = ~INSTADDRPOINTER_REG_16__SCAN_IN; 
assign R2027_U29 = ~INSTADDRPOINTER_REG_18__SCAN_IN; 
assign R2027_U30 = ~INSTADDRPOINTER_REG_17__SCAN_IN; 
assign R2027_U32 = ~INSTADDRPOINTER_REG_20__SCAN_IN; 
assign R2027_U33 = ~INSTADDRPOINTER_REG_19__SCAN_IN; 
assign R2027_U35 = ~INSTADDRPOINTER_REG_21__SCAN_IN; 
assign R2027_U37 = ~INSTADDRPOINTER_REG_22__SCAN_IN; 
assign R2027_U38 = ~INSTADDRPOINTER_REG_24__SCAN_IN; 
assign R2027_U39 = ~INSTADDRPOINTER_REG_23__SCAN_IN; 
assign R2027_U41 = ~INSTADDRPOINTER_REG_26__SCAN_IN; 
assign R2027_U42 = ~INSTADDRPOINTER_REG_25__SCAN_IN; 
assign R2027_U44 = ~INSTADDRPOINTER_REG_27__SCAN_IN; 
assign R2027_U45 = ~INSTADDRPOINTER_REG_28__SCAN_IN; 
assign R2027_U47 = ~INSTADDRPOINTER_REG_29__SCAN_IN; 
assign R2027_U50 = ~INSTADDRPOINTER_REG_30__SCAN_IN; 
assign R2027_U82 = INSTADDRPOINTER_REG_3__SCAN_IN & INSTADDRPOINTER_REG_4__SCAN_IN; 
assign R2027_U83 = INSTADDRPOINTER_REG_5__SCAN_IN & INSTADDRPOINTER_REG_6__SCAN_IN; 
assign R2027_U84 = INSTADDRPOINTER_REG_7__SCAN_IN & INSTADDRPOINTER_REG_8__SCAN_IN; 
assign R2027_U85 = INSTADDRPOINTER_REG_9__SCAN_IN & INSTADDRPOINTER_REG_10__SCAN_IN; 
assign R2027_U86 = INSTADDRPOINTER_REG_11__SCAN_IN & INSTADDRPOINTER_REG_12__SCAN_IN; 
assign R2027_U87 = INSTADDRPOINTER_REG_13__SCAN_IN & INSTADDRPOINTER_REG_14__SCAN_IN; 
assign R2027_U88 = INSTADDRPOINTER_REG_15__SCAN_IN & INSTADDRPOINTER_REG_16__SCAN_IN; 
assign R2027_U89 = INSTADDRPOINTER_REG_17__SCAN_IN & INSTADDRPOINTER_REG_18__SCAN_IN; 
assign R2027_U90 = INSTADDRPOINTER_REG_19__SCAN_IN & INSTADDRPOINTER_REG_20__SCAN_IN; 
assign R2027_U91 = INSTADDRPOINTER_REG_21__SCAN_IN & INSTADDRPOINTER_REG_22__SCAN_IN; 
assign R2027_U92 = INSTADDRPOINTER_REG_23__SCAN_IN & INSTADDRPOINTER_REG_24__SCAN_IN; 
assign R2027_U93 = INSTADDRPOINTER_REG_25__SCAN_IN & INSTADDRPOINTER_REG_26__SCAN_IN; 
assign R2027_U94 = INSTADDRPOINTER_REG_27__SCAN_IN & INSTADDRPOINTER_REG_28__SCAN_IN; 
assign R2027_U98 = ~INSTADDRPOINTER_REG_31__SCAN_IN; 
assign R2027_U100 = ~(INSTADDRPOINTER_REG_0__SCAN_IN & INSTADDRPOINTER_REG_1__SCAN_IN); 
assign R2278_U21 = ~INSTADDRPOINTER_REG_30__SCAN_IN; 
assign R2278_U32 = ~INSTADDRPOINTER_REG_29__SCAN_IN; 
assign R2278_U34 = ~INSTADDRPOINTER_REG_28__SCAN_IN; 
assign R2278_U94 = ~INSTADDRPOINTER_REG_31__SCAN_IN; 
assign R2337_U5 = ~PHYADDRPOINTER_REG_1__SCAN_IN; 
assign R2337_U6 = ~PHYADDRPOINTER_REG_5__SCAN_IN; 
assign R2337_U7 = ~PHYADDRPOINTER_REG_4__SCAN_IN; 
assign R2337_U8 = ~PHYADDRPOINTER_REG_3__SCAN_IN; 
assign R2337_U9 = ~PHYADDRPOINTER_REG_2__SCAN_IN; 
assign R2337_U10 = ~(PHYADDRPOINTER_REG_1__SCAN_IN & PHYADDRPOINTER_REG_2__SCAN_IN & PHYADDRPOINTER_REG_3__SCAN_IN & PHYADDRPOINTER_REG_4__SCAN_IN & PHYADDRPOINTER_REG_5__SCAN_IN); 
assign R2337_U11 = ~PHYADDRPOINTER_REG_7__SCAN_IN; 
assign R2337_U12 = ~PHYADDRPOINTER_REG_6__SCAN_IN; 
assign R2337_U14 = ~PHYADDRPOINTER_REG_8__SCAN_IN; 
assign R2337_U15 = ~PHYADDRPOINTER_REG_9__SCAN_IN; 
assign R2337_U16 = ~(PHYADDRPOINTER_REG_1__SCAN_IN & PHYADDRPOINTER_REG_2__SCAN_IN & PHYADDRPOINTER_REG_3__SCAN_IN); 
assign R2337_U18 = ~PHYADDRPOINTER_REG_11__SCAN_IN; 
assign R2337_U19 = ~PHYADDRPOINTER_REG_10__SCAN_IN; 
assign R2337_U21 = ~PHYADDRPOINTER_REG_13__SCAN_IN; 
assign R2337_U22 = ~PHYADDRPOINTER_REG_12__SCAN_IN; 
assign R2337_U24 = ~PHYADDRPOINTER_REG_15__SCAN_IN; 
assign R2337_U25 = ~PHYADDRPOINTER_REG_14__SCAN_IN; 
assign R2337_U27 = ~PHYADDRPOINTER_REG_17__SCAN_IN; 
assign R2337_U28 = ~PHYADDRPOINTER_REG_16__SCAN_IN; 
assign R2337_U30 = ~PHYADDRPOINTER_REG_19__SCAN_IN; 
assign R2337_U31 = ~PHYADDRPOINTER_REG_18__SCAN_IN; 
assign R2337_U33 = ~PHYADDRPOINTER_REG_21__SCAN_IN; 
assign R2337_U34 = ~PHYADDRPOINTER_REG_20__SCAN_IN; 
assign R2337_U36 = ~PHYADDRPOINTER_REG_23__SCAN_IN; 
assign R2337_U37 = ~PHYADDRPOINTER_REG_22__SCAN_IN; 
assign R2337_U39 = ~PHYADDRPOINTER_REG_25__SCAN_IN; 
assign R2337_U40 = ~PHYADDRPOINTER_REG_24__SCAN_IN; 
assign R2337_U42 = ~PHYADDRPOINTER_REG_26__SCAN_IN; 
assign R2337_U44 = ~PHYADDRPOINTER_REG_27__SCAN_IN; 
assign R2337_U46 = ~PHYADDRPOINTER_REG_28__SCAN_IN; 
assign R2337_U48 = ~PHYADDRPOINTER_REG_29__SCAN_IN; 
assign R2337_U50 = ~PHYADDRPOINTER_REG_30__SCAN_IN; 
assign R2337_U81 = PHYADDRPOINTER_REG_6__SCAN_IN & PHYADDRPOINTER_REG_7__SCAN_IN; 
assign R2337_U82 = PHYADDRPOINTER_REG_8__SCAN_IN & PHYADDRPOINTER_REG_9__SCAN_IN; 
assign R2337_U83 = PHYADDRPOINTER_REG_10__SCAN_IN & PHYADDRPOINTER_REG_11__SCAN_IN; 
assign R2337_U84 = PHYADDRPOINTER_REG_12__SCAN_IN & PHYADDRPOINTER_REG_13__SCAN_IN; 
assign R2337_U85 = PHYADDRPOINTER_REG_14__SCAN_IN & PHYADDRPOINTER_REG_15__SCAN_IN; 
assign R2337_U86 = PHYADDRPOINTER_REG_16__SCAN_IN & PHYADDRPOINTER_REG_17__SCAN_IN; 
assign R2337_U87 = PHYADDRPOINTER_REG_18__SCAN_IN & PHYADDRPOINTER_REG_19__SCAN_IN; 
assign R2337_U88 = PHYADDRPOINTER_REG_20__SCAN_IN & PHYADDRPOINTER_REG_21__SCAN_IN; 
assign R2337_U89 = PHYADDRPOINTER_REG_22__SCAN_IN & PHYADDRPOINTER_REG_23__SCAN_IN; 
assign R2337_U90 = PHYADDRPOINTER_REG_24__SCAN_IN & PHYADDRPOINTER_REG_25__SCAN_IN; 
assign R2337_U94 = ~(PHYADDRPOINTER_REG_1__SCAN_IN & PHYADDRPOINTER_REG_2__SCAN_IN); 
assign R2337_U95 = ~PHYADDRPOINTER_REG_31__SCAN_IN; 
assign R2167_U16 = ~STATE2_REG_0__SCAN_IN; 
assign SUB_580_U7 = ~INSTADDRPOINTER_REG_1__SCAN_IN; 
assign SUB_580_U8 = ~INSTADDRPOINTER_REG_0__SCAN_IN; 
assign R2096_U4 = ~REIP_REG_1__SCAN_IN; 
assign R2096_U5 = ~REIP_REG_2__SCAN_IN; 
assign R2096_U6 = ~(REIP_REG_1__SCAN_IN & REIP_REG_2__SCAN_IN); 
assign R2096_U7 = ~REIP_REG_3__SCAN_IN; 
assign R2096_U9 = ~REIP_REG_4__SCAN_IN; 
assign R2096_U11 = ~REIP_REG_5__SCAN_IN; 
assign R2096_U13 = ~REIP_REG_6__SCAN_IN; 
assign R2096_U15 = ~REIP_REG_7__SCAN_IN; 
assign R2096_U17 = ~REIP_REG_8__SCAN_IN; 
assign R2096_U18 = ~REIP_REG_9__SCAN_IN; 
assign R2096_U21 = ~REIP_REG_10__SCAN_IN; 
assign R2096_U23 = ~REIP_REG_11__SCAN_IN; 
assign R2096_U25 = ~REIP_REG_12__SCAN_IN; 
assign R2096_U27 = ~REIP_REG_13__SCAN_IN; 
assign R2096_U29 = ~REIP_REG_14__SCAN_IN; 
assign R2096_U31 = ~REIP_REG_15__SCAN_IN; 
assign R2096_U33 = ~REIP_REG_16__SCAN_IN; 
assign R2096_U35 = ~REIP_REG_17__SCAN_IN; 
assign R2096_U37 = ~REIP_REG_18__SCAN_IN; 
assign R2096_U39 = ~REIP_REG_19__SCAN_IN; 
assign R2096_U41 = ~REIP_REG_20__SCAN_IN; 
assign R2096_U43 = ~REIP_REG_21__SCAN_IN; 
assign R2096_U45 = ~REIP_REG_22__SCAN_IN; 
assign R2096_U47 = ~REIP_REG_23__SCAN_IN; 
assign R2096_U49 = ~REIP_REG_24__SCAN_IN; 
assign R2096_U51 = ~REIP_REG_25__SCAN_IN; 
assign R2096_U53 = ~REIP_REG_26__SCAN_IN; 
assign R2096_U55 = ~REIP_REG_27__SCAN_IN; 
assign R2096_U57 = ~REIP_REG_28__SCAN_IN; 
assign R2096_U59 = ~REIP_REG_29__SCAN_IN; 
assign R2096_U61 = ~REIP_REG_30__SCAN_IN; 
assign R2096_U92 = ~REIP_REG_31__SCAN_IN; 
assign LT_563_U7 = ~INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign LT_563_U10 = ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign LT_563_U11 = ~INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign R2238_U8 = ~INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign R2238_U10 = ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign R2238_U11 = ~INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign R2238_U12 = ~INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign R2238_U13 = ~INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign R2238_U14 = ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign R2238_U15 = ~INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign R2238_U17 = ~INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign R2238_U18 = ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN; 
assign R2238_U29 = ~INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign SUB_450_U8 = ~INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign SUB_450_U10 = ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN; 
assign SUB_450_U11 = ~INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign SUB_450_U12 = ~INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign SUB_450_U13 = ~INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign SUB_450_U14 = ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN; 
assign SUB_450_U15 = ~INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign SUB_450_U17 = ~INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign SUB_450_U18 = ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN; 
assign SUB_450_U29 = ~INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign ADD_405_U4 = ~INSTADDRPOINTER_REG_0__SCAN_IN; 
assign ADD_405_U6 = ~INSTADDRPOINTER_REG_1__SCAN_IN; 
assign ADD_405_U7 = ~INSTADDRPOINTER_REG_3__SCAN_IN; 
assign ADD_405_U9 = ~INSTADDRPOINTER_REG_4__SCAN_IN; 
assign ADD_405_U11 = ~INSTADDRPOINTER_REG_5__SCAN_IN; 
assign ADD_405_U13 = ~INSTADDRPOINTER_REG_6__SCAN_IN; 
assign ADD_405_U15 = ~INSTADDRPOINTER_REG_7__SCAN_IN; 
assign ADD_405_U17 = ~INSTADDRPOINTER_REG_8__SCAN_IN; 
assign ADD_405_U18 = ~INSTADDRPOINTER_REG_9__SCAN_IN; 
assign ADD_405_U21 = ~INSTADDRPOINTER_REG_10__SCAN_IN; 
assign ADD_405_U23 = ~INSTADDRPOINTER_REG_11__SCAN_IN; 
assign ADD_405_U25 = ~INSTADDRPOINTER_REG_12__SCAN_IN; 
assign ADD_405_U27 = ~INSTADDRPOINTER_REG_13__SCAN_IN; 
assign ADD_405_U29 = ~INSTADDRPOINTER_REG_14__SCAN_IN; 
assign ADD_405_U31 = ~INSTADDRPOINTER_REG_15__SCAN_IN; 
assign ADD_405_U33 = ~INSTADDRPOINTER_REG_16__SCAN_IN; 
assign ADD_405_U35 = ~INSTADDRPOINTER_REG_17__SCAN_IN; 
assign ADD_405_U37 = ~INSTADDRPOINTER_REG_18__SCAN_IN; 
assign ADD_405_U39 = ~INSTADDRPOINTER_REG_19__SCAN_IN; 
assign ADD_405_U41 = ~INSTADDRPOINTER_REG_20__SCAN_IN; 
assign ADD_405_U43 = ~INSTADDRPOINTER_REG_21__SCAN_IN; 
assign ADD_405_U45 = ~INSTADDRPOINTER_REG_22__SCAN_IN; 
assign ADD_405_U47 = ~INSTADDRPOINTER_REG_23__SCAN_IN; 
assign ADD_405_U49 = ~INSTADDRPOINTER_REG_24__SCAN_IN; 
assign ADD_405_U51 = ~INSTADDRPOINTER_REG_25__SCAN_IN; 
assign ADD_405_U53 = ~INSTADDRPOINTER_REG_26__SCAN_IN; 
assign ADD_405_U55 = ~INSTADDRPOINTER_REG_27__SCAN_IN; 
assign ADD_405_U57 = ~INSTADDRPOINTER_REG_28__SCAN_IN; 
assign ADD_405_U59 = ~INSTADDRPOINTER_REG_29__SCAN_IN; 
assign ADD_405_U61 = ~INSTADDRPOINTER_REG_30__SCAN_IN; 
assign ADD_405_U62 = ~INSTADDRPOINTER_REG_2__SCAN_IN; 
assign ADD_405_U94 = ~INSTADDRPOINTER_REG_31__SCAN_IN; 
assign ADD_405_U96 = ~(INSTADDRPOINTER_REG_0__SCAN_IN & INSTADDRPOINTER_REG_1__SCAN_IN); 
assign ADD_405_U126 = ~(INSTADDRPOINTER_REG_0__SCAN_IN & INSTADDRPOINTER_REG_1__SCAN_IN & INSTADDRPOINTER_REG_2__SCAN_IN); 
assign ADD_515_U4 = ~INSTADDRPOINTER_REG_1__SCAN_IN; 
assign ADD_515_U5 = ~INSTADDRPOINTER_REG_2__SCAN_IN; 
assign ADD_515_U6 = ~(INSTADDRPOINTER_REG_1__SCAN_IN & INSTADDRPOINTER_REG_2__SCAN_IN); 
assign ADD_515_U7 = ~INSTADDRPOINTER_REG_3__SCAN_IN; 
assign ADD_515_U9 = ~INSTADDRPOINTER_REG_4__SCAN_IN; 
assign ADD_515_U11 = ~INSTADDRPOINTER_REG_5__SCAN_IN; 
assign ADD_515_U13 = ~INSTADDRPOINTER_REG_6__SCAN_IN; 
assign ADD_515_U15 = ~INSTADDRPOINTER_REG_7__SCAN_IN; 
assign ADD_515_U17 = ~INSTADDRPOINTER_REG_8__SCAN_IN; 
assign ADD_515_U18 = ~INSTADDRPOINTER_REG_9__SCAN_IN; 
assign ADD_515_U21 = ~INSTADDRPOINTER_REG_10__SCAN_IN; 
assign ADD_515_U23 = ~INSTADDRPOINTER_REG_11__SCAN_IN; 
assign ADD_515_U25 = ~INSTADDRPOINTER_REG_12__SCAN_IN; 
assign ADD_515_U27 = ~INSTADDRPOINTER_REG_13__SCAN_IN; 
assign ADD_515_U29 = ~INSTADDRPOINTER_REG_14__SCAN_IN; 
assign ADD_515_U31 = ~INSTADDRPOINTER_REG_15__SCAN_IN; 
assign ADD_515_U33 = ~INSTADDRPOINTER_REG_16__SCAN_IN; 
assign ADD_515_U35 = ~INSTADDRPOINTER_REG_17__SCAN_IN; 
assign ADD_515_U37 = ~INSTADDRPOINTER_REG_18__SCAN_IN; 
assign ADD_515_U39 = ~INSTADDRPOINTER_REG_19__SCAN_IN; 
assign ADD_515_U41 = ~INSTADDRPOINTER_REG_20__SCAN_IN; 
assign ADD_515_U43 = ~INSTADDRPOINTER_REG_21__SCAN_IN; 
assign ADD_515_U45 = ~INSTADDRPOINTER_REG_22__SCAN_IN; 
assign ADD_515_U47 = ~INSTADDRPOINTER_REG_23__SCAN_IN; 
assign ADD_515_U49 = ~INSTADDRPOINTER_REG_24__SCAN_IN; 
assign ADD_515_U51 = ~INSTADDRPOINTER_REG_25__SCAN_IN; 
assign ADD_515_U53 = ~INSTADDRPOINTER_REG_26__SCAN_IN; 
assign ADD_515_U55 = ~INSTADDRPOINTER_REG_27__SCAN_IN; 
assign ADD_515_U57 = ~INSTADDRPOINTER_REG_28__SCAN_IN; 
assign ADD_515_U59 = ~INSTADDRPOINTER_REG_29__SCAN_IN; 
assign ADD_515_U61 = ~INSTADDRPOINTER_REG_30__SCAN_IN; 
assign ADD_515_U92 = ~INSTADDRPOINTER_REG_31__SCAN_IN; 
assign U2430 = U3374 & STATE2_REG_1__SCAN_IN; 
assign U2454 = U3253 & INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign U2455 = U3253 & INSTQUEUERD_ADDR_REG_3__SCAN_IN & INSTQUEUERD_ADDR_REG_2__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign U2456 = U3252 & INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign U2457 = U3252 & INSTQUEUERD_ADDR_REG_3__SCAN_IN & INSTQUEUERD_ADDR_REG_2__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign U2459 = U3251 & INSTQUEUERD_ADDR_REG_3__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign U2460 = U3251 & U3253 & INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign U2461 = U3494 & U3493; 
assign U2462 = U3251 & U3252 & INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign U2463 = U3492 & U3491; 
assign U2465 = U3490 & U3489; 
assign U2466 = U3488 & U3487; 
assign U2468 = U3486 & U3485; 
assign U2470 = U3253 & U2469 & INSTQUEUERD_ADDR_REG_1__SCAN_IN; 
assign U2471 = U3252 & U2469 & INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign U2479 = U3290 & INSTQUEUEWR_ADDR_REG_2__SCAN_IN; 
assign U3236 = ~(U3245 & STATE_REG_1__SCAN_IN); 
assign U3241 = ~(U3238 & STATE_REG_1__SCAN_IN); 
assign U3247 = ~(U3243 & REQUESTPENDING_REG_SCAN_IN); 
assign U3254 = ~(U3257 & INSTQUEUERD_ADDR_REG_2__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U3261 = ~(U3257 & INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign U3284 = ~(U3249 & STATE2_REG_2__SCAN_IN); 
assign U3310 = ~(U3288 & INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign U3316 = ~(U3289 & INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign U3324 = ~(U2488 & U2478); 
assign U3327 = ~(U3291 & INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign U3371 = ~(U2510 & U2488); 
assign U3389 = ~(U3256 & U3262); 
assign U3395 = ~(U2427 & U3281); 
assign U3427 = ~(U3250 & STATEBS16_REG_SCAN_IN); 
assign U3431 = ~(U3251 & INSTQUEUERD_ADDR_REG_1__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U3450 = U3242 & U4167; 
assign U3571 = U2427 & U3244; 
assign U3940 = U3939 & U3938; 
assign U3943 = U3942 & U3941; 
assign U3946 = U3945 & U3944; 
assign U3950 = U3949 & U6586 & U3948 & U3947; 
assign U3952 = U3244 & STATE2_REG_2__SCAN_IN; 
assign U4145 = U2427 & STATE2_REG_0__SCAN_IN; 
assign U4171 = ~(U3256 & INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign U4173 = ~(HOLD & U3244); 
assign U4197 = ~U3294; 
assign U4230 = ~(U3719 & U2428); 
assign U4232 = ~(U3281 & U2352 & STATE2_REG_1__SCAN_IN); 
assign U4234 = ~(READY_N & U3250 & STATE2_REG_0__SCAN_IN); 
assign U4249 = ~U3285; 
assign U4348 = ~U3248; 
assign U4352 = ~U3242; 
assign U4354 = ~(U3481 & U3248); 
assign U4361 = ~(NA_N & U3245); 
assign U4364 = ~(U4167 & U3242); 
assign U4365 = ~U3267; 
assign U4366 = ~U3256; 
assign U4368 = ~U3255; 
assign U4386 = ~(U2453 & INSTQUEUE_REG_15__3__SCAN_IN); 
assign U4389 = ~(U3257 & INSTQUEUE_REG_7__5__SCAN_IN & INSTQUEUERD_ADDR_REG_2__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U4391 = ~(U2469 & U3252 & INSTQUEUE_REG_1__5__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U4392 = ~(U2469 & U3253 & INSTQUEUE_REG_2__5__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U4394 = ~(U3508 & U3509 & INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign U4395 = ~(U3510 & U3511 & INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign U4397 = ~(U3513 & U3514 & INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U4398 = ~(U3251 & INSTQUEUE_REG_11__5__SCAN_IN & INSTQUEUERD_ADDR_REG_3__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U4400 = ~(U3252 & INSTQUEUE_REG_13__5__SCAN_IN & INSTQUEUERD_ADDR_REG_3__SCAN_IN & INSTQUEUERD_ADDR_REG_2__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U4401 = ~(U3253 & INSTQUEUE_REG_14__5__SCAN_IN & INSTQUEUERD_ADDR_REG_3__SCAN_IN & INSTQUEUERD_ADDR_REG_2__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U4419 = ~(U2453 & INSTQUEUE_REG_15__2__SCAN_IN); 
assign U4436 = ~(U2453 & INSTQUEUE_REG_15__7__SCAN_IN); 
assign U4447 = ~(U3495 & U3486 & INSTQUEUE_REG_15__6__SCAN_IN); 
assign U4464 = ~(U2453 & INSTQUEUE_REG_15__1__SCAN_IN); 
assign U4481 = ~(U2453 & INSTQUEUE_REG_15__0__SCAN_IN); 
assign U4483 = ~(U3235 & STATE_REG_2__SCAN_IN); 
assign U4521 = ~U3292; 
assign U4527 = ~(U3292 & INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign U4534 = ~(U3250 & STATE2_REG_1__SCAN_IN); 
assign U5463 = ~(U3281 & STATE2_REG_3__SCAN_IN); 
assign U5466 = ~(U5465 & INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign U5469 = ~(U3486 & INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign U5472 = ~(U3262 & U3251); 
assign U5474 = ~(U2469 & U3262); 
assign U5498 = ~(U3262 & INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign U5526 = ~(U3283 & STATE2_REG_1__SCAN_IN); 
assign U5784 = ~(U3281 & STATE2_REG_2__SCAN_IN); 
assign U5785 = ~(U3295 & STATE2_REG_1__SCAN_IN); 
assign U6042 = ~(U2428 & U3281); 
assign U6590 = ~(U3954 & U2428); 
assign U6850 = ~(R2337_U5 & U2352); 
assign U6855 = ~(U2352 & PHYADDRPOINTER_REG_0__SCAN_IN); 
assign U7052 = ~(U3251 & INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign U7365 = ~(U3281 & INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign U7367 = ~(U3281 & INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign U7371 = ~(U3281 & INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign U7374 = ~(U3281 & INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U7377 = ~(U3281 & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U7629 = ~(U3238 & STATE_REG_0__SCAN_IN & REQUESTPENDING_REG_SCAN_IN); 
assign U7643 = ~(U3529 & U3528 & U3252); 
assign U7644 = ~(U3257 & INSTQUEUE_REG_7__4__SCAN_IN & INSTQUEUERD_ADDR_REG_2__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U7645 = ~(U3257 & U3252 & INSTQUEUE_REG_5__4__SCAN_IN & INSTQUEUERD_ADDR_REG_2__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U7646 = ~(U3257 & U3251 & U3253 & INSTQUEUE_REG_2__4__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U7647 = ~(U3531 & U3530 & U3257); 
assign U7648 = ~(U3533 & U3532 & INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign U7649 = ~(U3535 & U3534 & U3252); 
assign U7650 = ~(U3537 & U3536 & INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U7651 = ~(U3539 & U3538 & U3253); 
assign U7653 = ~(U3251 & U3252 & U3253 & U3257 & INSTQUEUE_REG_0__4__SCAN_IN); 
assign U7654 = ~(U3251 & U3252 & U3253 & INSTQUEUE_REG_8__4__SCAN_IN & INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign U7655 = ~(U3251 & U3253 & INSTQUEUE_REG_10__4__SCAN_IN & INSTQUEUERD_ADDR_REG_3__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U7656 = ~(U3541 & U3540 & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U7657 = ~(U3251 & U3257 & INSTQUEUE_REG_3__4__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U7658 = ~(U3251 & INSTQUEUE_REG_11__4__SCAN_IN & INSTQUEUERD_ADDR_REG_3__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U7659 = ~(U3251 & U3257 & INSTQUEUE_REG_3__5__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U7660 = ~(U3517 & U3516 & INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign U7661 = ~(U3251 & U3252 & INSTQUEUE_REG_9__6__SCAN_IN & INSTQUEUERD_ADDR_REG_3__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U7662 = ~(U3523 & U3522 & INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U7663 = ~(U3251 & U3253 & INSTQUEUE_REG_10__6__SCAN_IN & INSTQUEUERD_ADDR_REG_3__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U7664 = ~(U3251 & INSTQUEUE_REG_11__6__SCAN_IN & INSTQUEUERD_ADDR_REG_3__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U7665 = ~(U3251 & U3252 & U3253 & U3257 & INSTQUEUE_REG_0__6__SCAN_IN); 
assign U7666 = ~(U3251 & U3252 & U3253 & INSTQUEUE_REG_8__6__SCAN_IN & INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign U7672 = ~(U4501 & U3281); 
assign U7676 = ~(U7457 & STATE2_REG_0__SCAN_IN); 
assign U7682 = ~(U3292 & INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign U7698 = ~(U4162 & INSTADDRPOINTER_REG_1__SCAN_IN); 
assign U7701 = ~(U4162 & INSTADDRPOINTER_REG_0__SCAN_IN); 
assign U7706 = ~(U3251 & INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U7707 = ~(U3252 & INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign U7737 = ~(U3400 & DATAWIDTH_REG_0__SCAN_IN); 
assign R2027_U111 = ~R2027_U10; 
assign R2027_U130 = ~R2027_U100; 
assign R2027_U154 = ~(R2027_U10 & INSTADDRPOINTER_REG_3__SCAN_IN); 
assign R2027_U159 = ~(R2027_U100 & INSTADDRPOINTER_REG_2__SCAN_IN); 
assign R2027_U181 = ~(R2027_U7 & INSTADDRPOINTER_REG_0__SCAN_IN); 
assign R2027_U182 = ~(R2027_U5 & INSTADDRPOINTER_REG_1__SCAN_IN); 
assign R2358_U22 = ~U2352; 
assign R2337_U105 = ~R2337_U94; 
assign R2337_U106 = ~R2337_U16; 
assign R2337_U108 = ~R2337_U10; 
assign R2337_U140 = ~(R2337_U10 & PHYADDRPOINTER_REG_6__SCAN_IN); 
assign R2337_U144 = ~(R2337_U16 & PHYADDRPOINTER_REG_4__SCAN_IN); 
assign R2337_U146 = ~(R2337_U94 & PHYADDRPOINTER_REG_3__SCAN_IN); 
assign R2337_U152 = ~(R2337_U9 & PHYADDRPOINTER_REG_1__SCAN_IN); 
assign R2337_U153 = ~(R2337_U5 & PHYADDRPOINTER_REG_2__SCAN_IN); 
assign SUB_580_U9 = ~(SUB_580_U8 & INSTADDRPOINTER_REG_1__SCAN_IN); 
assign SUB_580_U10 = ~(SUB_580_U7 & INSTADDRPOINTER_REG_0__SCAN_IN); 
assign R2096_U94 = ~R2096_U6; 
assign R2096_U135 = ~(R2096_U6 & REIP_REG_3__SCAN_IN); 
assign R2096_U141 = ~(R2096_U4 & REIP_REG_2__SCAN_IN); 
assign R2096_U142 = ~(R2096_U5 & REIP_REG_1__SCAN_IN); 
assign R2238_U9 = ~(R2238_U18 & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign R2238_U35 = ~(R2238_U12 & INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign R2238_U37 = ~(R2238_U11 & INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign R2238_U39 = ~(R2238_U14 & INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign R2238_U41 = ~(R2238_U13 & INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign R2238_U43 = ~(R2238_U17 & INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign R2238_U45 = ~(R2238_U15 & INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign R2238_U46 = ~(R2238_U8 & INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign R2238_U47 = ~(R2238_U15 & INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign R2238_U48 = ~(R2238_U17 & INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign R2238_U52 = ~(R2238_U14 & INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign R2238_U53 = ~(R2238_U13 & INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign R2238_U57 = ~(R2238_U12 & INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign R2238_U58 = ~(R2238_U11 & INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign R2238_U62 = ~(R2238_U10 & INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign R2238_U63 = ~(R2238_U29 & INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign SUB_450_U9 = ~(SUB_450_U18 & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign SUB_450_U35 = ~(SUB_450_U12 & INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign SUB_450_U37 = ~(SUB_450_U11 & INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign SUB_450_U39 = ~(SUB_450_U14 & INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign SUB_450_U41 = ~(SUB_450_U13 & INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign SUB_450_U43 = ~(SUB_450_U17 & INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign SUB_450_U45 = ~(SUB_450_U15 & INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign SUB_450_U46 = ~(SUB_450_U8 & INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign SUB_450_U47 = ~(SUB_450_U15 & INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign SUB_450_U48 = ~(SUB_450_U17 & INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign SUB_450_U52 = ~(SUB_450_U14 & INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign SUB_450_U53 = ~(SUB_450_U13 & INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign SUB_450_U57 = ~(SUB_450_U12 & INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign SUB_450_U58 = ~(SUB_450_U11 & INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign SUB_450_U62 = ~(SUB_450_U10 & INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign SUB_450_U63 = ~(SUB_450_U29 & INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign ADD_405_U92 = ~(ADD_405_U62 & ADD_405_U96); 
assign ADD_405_U165 = ~(ADD_405_U4 & INSTADDRPOINTER_REG_1__SCAN_IN); 
assign ADD_405_U166 = ~(ADD_405_U6 & INSTADDRPOINTER_REG_0__SCAN_IN); 
assign ADD_515_U94 = ~ADD_515_U6; 
assign ADD_515_U135 = ~(ADD_515_U6 & INSTADDRPOINTER_REG_3__SCAN_IN); 
assign ADD_515_U141 = ~(ADD_515_U4 & INSTADDRPOINTER_REG_2__SCAN_IN); 
assign ADD_515_U142 = ~(ADD_515_U5 & INSTADDRPOINTER_REG_1__SCAN_IN); 
assign U2388 = U4197 & STATEBS16_REG_SCAN_IN; 
assign U2458 = U3495 & U4366; 
assign U2464 = U4368 & INSTQUEUERD_ADDR_REG_3__SCAN_IN; 
assign U2467 = U3257 & U4366 & INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign U2472 = U4368 & U3257; 
assign U2521 = U3389 & INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign U2524 = U3253 & U3389; 
assign U2607 = U7660 & U7659; 
assign U3222 = ~(U3316 & U3310); 
assign U3246 = ~(U3247 & STATE_REG_0__SCAN_IN); 
assign U3293 = ~(U4521 & U2478); 
assign U3307 = ~(U4197 & U3295); 
assign U3343 = ~(U2479 & U4521); 
assign U3357 = ~(U2488 & U2479); 
assign U3360 = ~(U2510 & U4521); 
assign U3388 = ~(U3431 & U5498); 
assign U3419 = ~(U4197 & U3249); 
assign U3420 = ~(U3950 & U3946 & U3943 & U3940); 
assign U3432 = ~(U3261 & U7052); 
assign U3439 = ~(U4171 & U3255); 
assign U3443 = ~(U7707 & U7706); 
assign U3458 = ~(U7702 & U7701); 
assign U3521 = U4402 & U4401; 
assign U3527 = U7666 & U7665 & U7664 & U7663; 
assign U3542 = U7646 & U7645 & U7644 & U7643; 
assign U3543 = U7650 & U7649 & U7648 & U7647; 
assign U3544 = U7654 & U7653 & U7652 & U7651; 
assign U3545 = U7658 & U7657 & U7656 & U7655; 
assign U3564 = U4402 & U4401; 
assign U3727 = U5463 & U4230; 
assign U3955 = U3294 & U3395 & U6590; 
assign U4059 = U4402 & U4401; 
assign U4158 = U7662 & U7661; 
assign U4175 = ~U3427; 
assign U4191 = ~U3395; 
assign U4209 = ~U3236; 
assign U4223 = ~U3284; 
assign U4229 = ~(U3572 & U4249); 
assign U4231 = ~(U4352 & U3245); 
assign U4246 = ~U3241; 
assign U4257 = ~(U3236 & ADDRESS_REG_29__SCAN_IN); 
assign U4260 = ~(U3236 & ADDRESS_REG_28__SCAN_IN); 
assign U4263 = ~(U3236 & ADDRESS_REG_27__SCAN_IN); 
assign U4266 = ~(U3236 & ADDRESS_REG_26__SCAN_IN); 
assign U4269 = ~(U3236 & ADDRESS_REG_25__SCAN_IN); 
assign U4272 = ~(U3236 & ADDRESS_REG_24__SCAN_IN); 
assign U4275 = ~(U3236 & ADDRESS_REG_23__SCAN_IN); 
assign U4278 = ~(U3236 & ADDRESS_REG_22__SCAN_IN); 
assign U4281 = ~(U3236 & ADDRESS_REG_21__SCAN_IN); 
assign U4284 = ~(U3236 & ADDRESS_REG_20__SCAN_IN); 
assign U4287 = ~(U3236 & ADDRESS_REG_19__SCAN_IN); 
assign U4290 = ~(U3236 & ADDRESS_REG_18__SCAN_IN); 
assign U4293 = ~(U3236 & ADDRESS_REG_17__SCAN_IN); 
assign U4296 = ~(U3236 & ADDRESS_REG_16__SCAN_IN); 
assign U4299 = ~(U3236 & ADDRESS_REG_15__SCAN_IN); 
assign U4302 = ~(U3236 & ADDRESS_REG_14__SCAN_IN); 
assign U4305 = ~(U3236 & ADDRESS_REG_13__SCAN_IN); 
assign U4308 = ~(U3236 & ADDRESS_REG_12__SCAN_IN); 
assign U4311 = ~(U3236 & ADDRESS_REG_11__SCAN_IN); 
assign U4314 = ~(U3236 & ADDRESS_REG_10__SCAN_IN); 
assign U4317 = ~(U3236 & ADDRESS_REG_9__SCAN_IN); 
assign U4320 = ~(U3236 & ADDRESS_REG_8__SCAN_IN); 
assign U4323 = ~(U3236 & ADDRESS_REG_7__SCAN_IN); 
assign U4326 = ~(U3236 & ADDRESS_REG_6__SCAN_IN); 
assign U4329 = ~(U3236 & ADDRESS_REG_5__SCAN_IN); 
assign U4332 = ~(U3236 & ADDRESS_REG_4__SCAN_IN); 
assign U4335 = ~(U3236 & ADDRESS_REG_3__SCAN_IN); 
assign U4338 = ~(U3236 & ADDRESS_REG_2__SCAN_IN); 
assign U4341 = ~(U3236 & ADDRESS_REG_1__SCAN_IN); 
assign U4344 = ~(U3236 & ADDRESS_REG_0__SCAN_IN); 
assign U4345 = ~U3247; 
assign U4349 = ~(U4348 & U3244); 
assign U4353 = ~(HOLD & U3234 & U4352); 
assign U4360 = ~(U3247 & STATE_REG_2__SCAN_IN); 
assign U4367 = ~U3431; 
assign U4369 = ~U3261; 
assign U4370 = ~U3254; 
assign U4373 = ~(U2471 & INSTQUEUE_REG_1__3__SCAN_IN); 
assign U4374 = ~(U2470 & INSTQUEUE_REG_2__3__SCAN_IN); 
assign U4375 = ~(U2468 & INSTQUEUE_REG_3__3__SCAN_IN); 
assign U4377 = ~(U2466 & INSTQUEUE_REG_5__3__SCAN_IN); 
assign U4378 = ~(U2465 & INSTQUEUE_REG_6__3__SCAN_IN); 
assign U4380 = ~(U2463 & INSTQUEUE_REG_9__3__SCAN_IN); 
assign U4381 = ~(U2461 & INSTQUEUE_REG_10__3__SCAN_IN); 
assign U4382 = ~(U2459 & INSTQUEUE_REG_11__3__SCAN_IN); 
assign U4384 = ~(U2457 & INSTQUEUE_REG_13__3__SCAN_IN); 
assign U4385 = ~(U2455 & INSTQUEUE_REG_14__3__SCAN_IN); 
assign U4390 = ~(U3257 & U4368 & INSTQUEUE_REG_0__5__SCAN_IN); 
assign U4393 = ~(U4366 & U3257 & INSTQUEUE_REG_4__5__SCAN_IN & INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign U4396 = ~(U3512 & U4368); 
assign U4399 = ~(U4366 & U3515 & INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign U4406 = ~(U2471 & INSTQUEUE_REG_1__2__SCAN_IN); 
assign U4407 = ~(U2470 & INSTQUEUE_REG_2__2__SCAN_IN); 
assign U4408 = ~(U2468 & INSTQUEUE_REG_3__2__SCAN_IN); 
assign U4410 = ~(U2466 & INSTQUEUE_REG_5__2__SCAN_IN); 
assign U4411 = ~(U2465 & INSTQUEUE_REG_6__2__SCAN_IN); 
assign U4413 = ~(U2463 & INSTQUEUE_REG_9__2__SCAN_IN); 
assign U4414 = ~(U2461 & INSTQUEUE_REG_10__2__SCAN_IN); 
assign U4415 = ~(U2459 & INSTQUEUE_REG_11__2__SCAN_IN); 
assign U4417 = ~(U2457 & INSTQUEUE_REG_13__2__SCAN_IN); 
assign U4418 = ~(U2455 & INSTQUEUE_REG_14__2__SCAN_IN); 
assign U4423 = ~(U2471 & INSTQUEUE_REG_1__7__SCAN_IN); 
assign U4424 = ~(U2470 & INSTQUEUE_REG_2__7__SCAN_IN); 
assign U4425 = ~(U2468 & INSTQUEUE_REG_3__7__SCAN_IN); 
assign U4427 = ~(U2466 & INSTQUEUE_REG_5__7__SCAN_IN); 
assign U4428 = ~(U2465 & INSTQUEUE_REG_6__7__SCAN_IN); 
assign U4430 = ~(U2463 & INSTQUEUE_REG_9__7__SCAN_IN); 
assign U4431 = ~(U2461 & INSTQUEUE_REG_10__7__SCAN_IN); 
assign U4432 = ~(U2459 & INSTQUEUE_REG_11__7__SCAN_IN); 
assign U4434 = ~(U2457 & INSTQUEUE_REG_13__7__SCAN_IN); 
assign U4435 = ~(U2455 & INSTQUEUE_REG_14__7__SCAN_IN); 
assign U4439 = ~(U2469 & U2456 & INSTQUEUE_REG_1__6__SCAN_IN); 
assign U4440 = ~(U2469 & U2454 & INSTQUEUE_REG_2__6__SCAN_IN); 
assign U4444 = ~(U4366 & U3495 & INSTQUEUE_REG_12__6__SCAN_IN); 
assign U4445 = ~(U3495 & U2456 & INSTQUEUE_REG_13__6__SCAN_IN); 
assign U4446 = ~(U3495 & U2454 & INSTQUEUE_REG_14__6__SCAN_IN); 
assign U4451 = ~(U2471 & INSTQUEUE_REG_1__1__SCAN_IN); 
assign U4452 = ~(U2470 & INSTQUEUE_REG_2__1__SCAN_IN); 
assign U4453 = ~(U2468 & INSTQUEUE_REG_3__1__SCAN_IN); 
assign U4455 = ~(U2466 & INSTQUEUE_REG_5__1__SCAN_IN); 
assign U4456 = ~(U2465 & INSTQUEUE_REG_6__1__SCAN_IN); 
assign U4458 = ~(U2463 & INSTQUEUE_REG_9__1__SCAN_IN); 
assign U4459 = ~(U2461 & INSTQUEUE_REG_10__1__SCAN_IN); 
assign U4460 = ~(U2459 & INSTQUEUE_REG_11__1__SCAN_IN); 
assign U4462 = ~(U2457 & INSTQUEUE_REG_13__1__SCAN_IN); 
assign U4463 = ~(U2455 & INSTQUEUE_REG_14__1__SCAN_IN); 
assign U4468 = ~(U2471 & INSTQUEUE_REG_1__0__SCAN_IN); 
assign U4469 = ~(U2470 & INSTQUEUE_REG_2__0__SCAN_IN); 
assign U4470 = ~(U2468 & INSTQUEUE_REG_3__0__SCAN_IN); 
assign U4472 = ~(U2466 & INSTQUEUE_REG_5__0__SCAN_IN); 
assign U4473 = ~(U2465 & INSTQUEUE_REG_6__0__SCAN_IN); 
assign U4475 = ~(U2463 & INSTQUEUE_REG_9__0__SCAN_IN); 
assign U4476 = ~(U2461 & INSTQUEUE_REG_10__0__SCAN_IN); 
assign U4477 = ~(U2459 & INSTQUEUE_REG_11__0__SCAN_IN); 
assign U4479 = ~(U2457 & INSTQUEUE_REG_13__0__SCAN_IN); 
assign U4480 = ~(U2455 & INSTQUEUE_REG_14__0__SCAN_IN); 
assign U4484 = ~(U3241 & U4483); 
assign U4503 = ~(U7676 & U7675 & STATE2_REG_1__SCAN_IN); 
assign U4526 = ~U3327; 
assign U4529 = ~U3316; 
assign U4530 = ~U3310; 
assign U4706 = ~U3324; 
assign U4714 = ~(U3324 & STATE2_REG_3__SCAN_IN); 
assign U5394 = ~U3371; 
assign U5402 = ~(U3371 & STATE2_REG_3__SCAN_IN); 
assign U5470 = ~(U5469 & INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign U5473 = ~(U5472 & INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign U5507 = ~U3389; 
assign U5782 = ~(U4197 & U3281); 
assign U5786 = ~(U5785 & U5784); 
assign U7083 = ~(U3284 & INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign U7203 = ~(U3284 & INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign U7205 = ~(U3284 & INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign U7207 = ~U4171; 
assign U7445 = ~(U2430 & INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign U7447 = ~(U2430 & INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign U7450 = ~(U2430 & INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign U7453 = ~(U2430 & INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U7455 = ~(U2430 & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U7456 = ~(U4173 & STATE_REG_0__SCAN_IN); 
assign U7621 = ~(U3236 & BE_N_REG_3__SCAN_IN); 
assign U7623 = ~(U3236 & BE_N_REG_2__SCAN_IN); 
assign U7625 = ~(U3236 & BE_N_REG_1__SCAN_IN); 
assign U7627 = ~(U3236 & BE_N_REG_0__SCAN_IN); 
assign U7634 = ~(U3247 & STATE_REG_2__SCAN_IN & STATE_REG_0__SCAN_IN); 
assign U7683 = ~(U4521 & U3291); 
assign U7738 = ~(U7737 & U7736); 
assign U7749 = ~(U3236 & W_R_N_REG_SCAN_IN); 
assign U7757 = ~(U3236 & D_C_N_REG_SCAN_IN); 
assign U7758 = ~(U3236 & M_IO_N_REG_SCAN_IN); 
assign U7775 = ~(U3284 & INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign U7776 = ~(U4171 & INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign R2027_U13 = ~(R2027_U82 & R2027_U111); 
assign R2027_U71 = ~(R2027_U182 & R2027_U181); 
assign R2027_U97 = ~(R2027_U111 & INSTADDRPOINTER_REG_3__SCAN_IN); 
assign R2027_U153 = ~(R2027_U111 & R2027_U9); 
assign R2027_U160 = ~(R2027_U130 & R2027_U6); 
assign R2337_U13 = ~(R2337_U81 & R2337_U108); 
assign R2337_U60 = ~(R2337_U153 & R2337_U152); 
assign R2337_U92 = ~(R2337_U108 & PHYADDRPOINTER_REG_6__SCAN_IN); 
assign R2337_U93 = ~(R2337_U106 & PHYADDRPOINTER_REG_4__SCAN_IN); 
assign R2337_U141 = ~(R2337_U108 & R2337_U12); 
assign R2337_U145 = ~(R2337_U106 & R2337_U7); 
assign R2337_U147 = ~(R2337_U105 & R2337_U8); 
assign SUB_580_U6 = ~(SUB_580_U10 & SUB_580_U9); 
assign R2096_U8 = ~(R2096_U94 & REIP_REG_3__SCAN_IN); 
assign R2096_U71 = ~(R2096_U142 & R2096_U141); 
assign R2096_U136 = ~(R2096_U94 & R2096_U7); 
assign R2238_U7 = ~(R2238_U9 & R2238_U46); 
assign R2238_U23 = ~(R2238_U48 & R2238_U47); 
assign R2238_U24 = ~(R2238_U53 & R2238_U52); 
assign R2238_U25 = ~(R2238_U58 & R2238_U57); 
assign R2238_U26 = ~(R2238_U63 & R2238_U62); 
assign R2238_U30 = ~R2238_U9; 
assign R2238_U33 = ~(R2238_U9 & INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign SUB_450_U7 = ~(SUB_450_U9 & SUB_450_U46); 
assign SUB_450_U23 = ~(SUB_450_U48 & SUB_450_U47); 
assign SUB_450_U24 = ~(SUB_450_U53 & SUB_450_U52); 
assign SUB_450_U25 = ~(SUB_450_U58 & SUB_450_U57); 
assign SUB_450_U26 = ~(SUB_450_U63 & SUB_450_U62); 
assign SUB_450_U30 = ~SUB_450_U9; 
assign SUB_450_U33 = ~(SUB_450_U9 & INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign ADD_405_U5 = ~(ADD_405_U92 & ADD_405_U126); 
assign ADD_405_U8 = ~(ADD_405_U92 & INSTADDRPOINTER_REG_3__SCAN_IN); 
assign ADD_405_U81 = ~(ADD_405_U166 & ADD_405_U165); 
assign ADD_405_U97 = ~ADD_405_U92; 
assign ADD_405_U139 = ~(ADD_405_U92 & INSTADDRPOINTER_REG_3__SCAN_IN); 
assign ADD_515_U8 = ~(ADD_515_U94 & INSTADDRPOINTER_REG_3__SCAN_IN); 
assign ADD_515_U71 = ~(ADD_515_U142 & ADD_515_U141); 
assign ADD_515_U136 = ~(ADD_515_U94 & ADD_515_U7); 
assign U2368 = U4223 & STATE2_REG_0__SCAN_IN; 
assign U2436 = U3222 & U3288; 
assign U2446 = U3458 & STATE2_REG_1__SCAN_IN; 
assign U2526 = U5507 & INSTQUEUERD_ADDR_REG_0__SCAN_IN; 
assign U2528 = U5507 & U3253; 
assign U2574 = U4367 & U3432; 
assign U2575 = U2460 & U3432; 
assign U2576 = U2462 & U3432; 
assign U2577 = U4368 & U3432; 
assign U2578 = U3432 & INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign U3237 = ~(U4209 & U3238); 
assign U3239 = ~(U4209 & STATE_REG_2__SCAN_IN); 
assign U3259 = ~(U4484 & U3245); 
assign U3265 = ~(U3545 & U3544 & U3543 & U3542); 
assign U3311 = ~(U4530 & U2478); 
assign U3317 = ~(U4529 & U2478); 
assign U3328 = ~(U4526 & U4521); 
assign U3333 = ~(U4526 & U4530); 
assign U3336 = ~(U4526 & U4529); 
assign U3340 = ~(U4526 & U2488); 
assign U3347 = ~(U3327 & U4527 & U3343); 
assign U3350 = ~(U4530 & U2479); 
assign U3353 = ~(U4529 & U2479); 
assign U3364 = ~(U2510 & U4530); 
assign U3367 = ~(U2510 & U4529); 
assign U3425 = ~(U3254 & U5470); 
assign U3442 = ~(U7683 & U7682); 
assign U3518 = U4392 & U4391 & U4390 & U4389; 
assign U3519 = U4396 & U4395 & U4394 & U4393; 
assign U3520 = U4400 & U4399 & U4398 & U4397; 
assign U3526 = U4446 & U4445 & U4447; 
assign U3561 = U4392 & U4391 & U4390 & U4389; 
assign U3562 = U4396 & U4395 & U4394 & U4393; 
assign U3563 = U4400 & U4399 & U4398 & U4397; 
assign U3570 = U4503 & U3284; 
assign U3573 = U4234 & U4229; 
assign U3728 = U5474 & U5473; 
assign U3851 = U5782 & U3395; 
assign U4056 = U4393 & U4392 & U4391 & U4389; 
assign U4057 = U4395 & U4394 & U4396; 
assign U4058 = U4400 & U4399 & U4398 & U4397; 
assign U4096 = U7203 & U3251; 
assign U4098 = U7205 & U3252; 
assign U4172 = ~U3439; 
assign U4208 = ~U3420; 
assign U4214 = ~U3307; 
assign U4243 = ~U3419; 
assign U4346 = ~(U4345 & U3244); 
assign U4347 = ~(NA_N & U4246); 
assign U4355 = ~(U4354 & U4353); 
assign U4358 = ~(READY_N & U4209); 
assign U4362 = ~(U4361 & U4360); 
assign U4371 = ~(U4370 & INSTQUEUE_REG_7__3__SCAN_IN); 
assign U4372 = ~(U2472 & INSTQUEUE_REG_0__3__SCAN_IN); 
assign U4376 = ~(U2467 & INSTQUEUE_REG_4__3__SCAN_IN); 
assign U4379 = ~(U2464 & INSTQUEUE_REG_8__3__SCAN_IN); 
assign U4383 = ~(U2458 & INSTQUEUE_REG_12__3__SCAN_IN); 
assign U4404 = ~(U4370 & INSTQUEUE_REG_7__2__SCAN_IN); 
assign U4405 = ~(U2472 & INSTQUEUE_REG_0__2__SCAN_IN); 
assign U4409 = ~(U2467 & INSTQUEUE_REG_4__2__SCAN_IN); 
assign U4412 = ~(U2464 & INSTQUEUE_REG_8__2__SCAN_IN); 
assign U4416 = ~(U2458 & INSTQUEUE_REG_12__2__SCAN_IN); 
assign U4421 = ~(U4370 & INSTQUEUE_REG_7__7__SCAN_IN); 
assign U4422 = ~(U2472 & INSTQUEUE_REG_0__7__SCAN_IN); 
assign U4426 = ~(U2467 & INSTQUEUE_REG_4__7__SCAN_IN); 
assign U4429 = ~(U2464 & INSTQUEUE_REG_8__7__SCAN_IN); 
assign U4433 = ~(U2458 & INSTQUEUE_REG_12__7__SCAN_IN); 
assign U4438 = ~(U3486 & U4369 & INSTQUEUE_REG_7__6__SCAN_IN); 
assign U4441 = ~(U4366 & U4369 & INSTQUEUE_REG_4__6__SCAN_IN); 
assign U4442 = ~(U2456 & U4369 & INSTQUEUE_REG_5__6__SCAN_IN); 
assign U4443 = ~(U2454 & U4369 & INSTQUEUE_REG_6__6__SCAN_IN); 
assign U4449 = ~(U4370 & INSTQUEUE_REG_7__1__SCAN_IN); 
assign U4450 = ~(U2472 & INSTQUEUE_REG_0__1__SCAN_IN); 
assign U4454 = ~(U2467 & INSTQUEUE_REG_4__1__SCAN_IN); 
assign U4457 = ~(U2464 & INSTQUEUE_REG_8__1__SCAN_IN); 
assign U4461 = ~(U2458 & INSTQUEUE_REG_12__1__SCAN_IN); 
assign U4466 = ~(U4370 & INSTQUEUE_REG_7__0__SCAN_IN); 
assign U4467 = ~(U2472 & INSTQUEUE_REG_0__0__SCAN_IN); 
assign U4471 = ~(U2467 & INSTQUEUE_REG_4__0__SCAN_IN); 
assign U4474 = ~(U2464 & INSTQUEUE_REG_8__0__SCAN_IN); 
assign U4478 = ~(U2458 & INSTQUEUE_REG_12__0__SCAN_IN); 
assign U4522 = ~U3293; 
assign U4525 = ~U3343; 
assign U4531 = ~U3222; 
assign U4540 = ~(U3293 & STATE2_REG_3__SCAN_IN); 
assign U5000 = ~(U3343 & STATE2_REG_3__SCAN_IN); 
assign U5164 = ~U3357; 
assign U5172 = ~(U3357 & STATE2_REG_3__SCAN_IN); 
assign U5221 = ~U3360; 
assign U5230 = ~(U3360 & STATE2_REG_3__SCAN_IN); 
assign U5467 = ~(U4369 & INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U5499 = ~U3388; 
assign U5551 = ~(U4191 & U3250); 
assign U6350 = ~(U4191 & U3250); 
assign U6736 = ~(U4175 & PHYADDRPOINTER_REG_9__SCAN_IN); 
assign U6739 = ~(U4175 & PHYADDRPOINTER_REG_8__SCAN_IN); 
assign U6742 = ~(U4175 & PHYADDRPOINTER_REG_7__SCAN_IN); 
assign U6745 = ~(U4175 & PHYADDRPOINTER_REG_6__SCAN_IN); 
assign U6749 = ~(U4175 & PHYADDRPOINTER_REG_5__SCAN_IN); 
assign U6753 = ~(U4175 & PHYADDRPOINTER_REG_4__SCAN_IN); 
assign U6757 = ~(U4175 & PHYADDRPOINTER_REG_31__SCAN_IN); 
assign U6761 = ~(U4175 & PHYADDRPOINTER_REG_30__SCAN_IN); 
assign U6765 = ~(U4175 & PHYADDRPOINTER_REG_3__SCAN_IN); 
assign U6770 = ~(U4175 & PHYADDRPOINTER_REG_29__SCAN_IN); 
assign U6774 = ~(U4175 & PHYADDRPOINTER_REG_28__SCAN_IN); 
assign U6778 = ~(U4175 & PHYADDRPOINTER_REG_27__SCAN_IN); 
assign U6782 = ~(U4175 & PHYADDRPOINTER_REG_26__SCAN_IN); 
assign U6786 = ~(U4175 & PHYADDRPOINTER_REG_25__SCAN_IN); 
assign U6790 = ~(U4175 & PHYADDRPOINTER_REG_24__SCAN_IN); 
assign U6794 = ~(U4175 & PHYADDRPOINTER_REG_23__SCAN_IN); 
assign U6798 = ~(U4175 & PHYADDRPOINTER_REG_22__SCAN_IN); 
assign U6802 = ~(U4175 & PHYADDRPOINTER_REG_21__SCAN_IN); 
assign U6806 = ~(U4175 & PHYADDRPOINTER_REG_20__SCAN_IN); 
assign U6810 = ~(U4175 & PHYADDRPOINTER_REG_2__SCAN_IN); 
assign U6811 = ~(R2337_U60 & U2352); 
assign U6815 = ~(U4175 & PHYADDRPOINTER_REG_19__SCAN_IN); 
assign U6819 = ~(U4175 & PHYADDRPOINTER_REG_18__SCAN_IN); 
assign U6823 = ~(U4175 & PHYADDRPOINTER_REG_17__SCAN_IN); 
assign U6827 = ~(U4175 & PHYADDRPOINTER_REG_16__SCAN_IN); 
assign U6830 = ~(U4175 & PHYADDRPOINTER_REG_15__SCAN_IN); 
assign U6833 = ~(U4175 & PHYADDRPOINTER_REG_14__SCAN_IN); 
assign U6836 = ~(U4175 & PHYADDRPOINTER_REG_13__SCAN_IN); 
assign U6839 = ~(U4175 & PHYADDRPOINTER_REG_12__SCAN_IN); 
assign U6842 = ~(U4175 & PHYADDRPOINTER_REG_11__SCAN_IN); 
assign U6845 = ~(U4175 & PHYADDRPOINTER_REG_10__SCAN_IN); 
assign U6849 = ~(U4175 & PHYADDRPOINTER_REG_1__SCAN_IN); 
assign U6854 = ~(U4175 & PHYADDRPOINTER_REG_0__SCAN_IN); 
assign U7053 = ~U3432; 
assign U7206 = ~(U4191 & U3222); 
assign U7609 = ~U3246; 
assign U7612 = ~(U7456 & STATE_REG_2__SCAN_IN); 
assign U7622 = ~(U4209 & BYTEENABLE_REG_3__SCAN_IN); 
assign U7624 = ~(U4209 & BYTEENABLE_REG_2__SCAN_IN); 
assign U7626 = ~(U4209 & BYTEENABLE_REG_1__SCAN_IN); 
assign U7628 = ~(U4209 & BYTEENABLE_REG_0__SCAN_IN); 
assign U7630 = ~(U3246 & STATE_REG_2__SCAN_IN); 
assign U7637 = ~(U4246 & STATE_REG_0__SCAN_IN); 
assign U7699 = ~(SUB_580_U6 & INSTADDRPOINTER_REG_31__SCAN_IN); 
assign U7703 = ~U3458; 
assign U7708 = ~U3443; 
assign U7734 = ~(U3420 & BYTEENABLE_REG_3__SCAN_IN); 
assign U7739 = ~(U7738 & U3240); 
assign U7742 = ~(U3420 & BYTEENABLE_REG_2__SCAN_IN); 
assign U7744 = ~(U3420 & BYTEENABLE_REG_1__SCAN_IN); 
assign U7746 = ~(U3420 & BYTEENABLE_REG_0__SCAN_IN); 
assign U7748 = ~(U4209 & U3423); 
assign U7756 = ~(U4209 & U3422); 
assign U7759 = ~(U4209 & MEMORYFETCH_REG_SCAN_IN); 
assign U7774 = ~(U4191 & U3288); 
assign U7777 = ~(U7207 & U3257); 
assign R2027_U57 = ~(R2027_U154 & R2027_U153); 
assign R2027_U60 = ~(R2027_U160 & R2027_U159); 
assign R2027_U112 = ~R2027_U13; 
assign R2027_U127 = ~R2027_U97; 
assign R2027_U150 = ~(R2027_U13 & INSTADDRPOINTER_REG_5__SCAN_IN); 
assign R2027_U151 = ~(R2027_U97 & INSTADDRPOINTER_REG_4__SCAN_IN); 
assign R2337_U54 = ~(R2337_U141 & R2337_U140); 
assign R2337_U56 = ~(R2337_U145 & R2337_U144); 
assign R2337_U57 = ~(R2337_U147 & R2337_U146); 
assign R2337_U107 = ~R2337_U93; 
assign R2337_U109 = ~R2337_U92; 
assign R2337_U110 = ~R2337_U13; 
assign R2337_U136 = ~(R2337_U13 & PHYADDRPOINTER_REG_8__SCAN_IN); 
assign R2337_U138 = ~(R2337_U92 & PHYADDRPOINTER_REG_7__SCAN_IN); 
assign R2337_U142 = ~(R2337_U93 & PHYADDRPOINTER_REG_5__SCAN_IN); 
assign R2096_U68 = ~(R2096_U136 & R2096_U135); 
assign R2096_U95 = ~R2096_U8; 
assign R2096_U133 = ~(R2096_U8 & REIP_REG_4__SCAN_IN); 
assign R2238_U31 = ~(R2238_U30 & R2238_U10); 
assign R2238_U49 = ~R2238_U23; 
assign R2238_U54 = ~R2238_U24; 
assign R2238_U59 = ~R2238_U25; 
assign R2238_U64 = ~R2238_U26; 
assign R2238_U66 = ~(R2238_U26 & R2238_U9); 
assign SUB_450_U31 = ~(SUB_450_U30 & SUB_450_U10); 
assign SUB_450_U49 = ~SUB_450_U23; 
assign SUB_450_U54 = ~SUB_450_U24; 
assign SUB_450_U59 = ~SUB_450_U25; 
assign SUB_450_U64 = ~SUB_450_U26; 
assign SUB_450_U66 = ~(SUB_450_U26 & SUB_450_U9); 
assign ADD_405_U98 = ~ADD_405_U8; 
assign ADD_405_U137 = ~(ADD_405_U8 & INSTADDRPOINTER_REG_4__SCAN_IN); 
assign ADD_405_U140 = ~(ADD_405_U97 & ADD_405_U7); 
assign ADD_515_U68 = ~(ADD_515_U136 & ADD_515_U135); 
assign ADD_515_U95 = ~ADD_515_U8; 
assign ADD_515_U133 = ~(ADD_515_U8 & INSTADDRPOINTER_REG_4__SCAN_IN); 
assign U2432 = U3442 & U3347; 
assign U2437 = U4531 & U3288; 
assign U2535 = U5499 & U3425; 
assign U2540 = U3425 & U3388; 
assign U2565 = U7053 & U4367; 
assign U2566 = U7053 & U2460; 
assign U2567 = U7053 & U2462; 
assign U2568 = U7053 & U4368; 
assign U2569 = U7053 & INSTQUEUERD_ADDR_REG_2__SCAN_IN; 
assign U2579 = U2578 & U3486; 
assign U2580 = U2578 & U2454; 
assign U2581 = U2578 & U2456; 
assign U2582 = U2578 & U4366; 
assign U2605 = U3521 & U2607 & U3520 & U3519 & U3518; 
assign U2608 = U7775 & U7774; 
assign U2791 = ~(U7757 & U7756 & U4231); 
assign U3429 = ~(U5467 & U5466); 
assign U3444 = ~(U7777 & U7776); 
assign U3445 = ~(U7622 & U7621); 
assign U3446 = ~(U7624 & U7623); 
assign U3447 = ~(U7626 & U7625); 
assign U3448 = ~(U7628 & U7627); 
assign U3449 = ~(U7637 & U7636); 
assign U3457 = ~(U7699 & U7698); 
assign U3470 = ~(U7749 & U7748); 
assign U3473 = ~(U7759 & U7758); 
assign U3483 = U4358 & U3237; 
assign U3496 = U4374 & U4373 & U4372 & U4371; 
assign U3497 = U4378 & U4377 & U4376 & U4375; 
assign U3498 = U4382 & U4381 & U4380 & U4379; 
assign U3499 = U4386 & U4385 & U4384 & U4383; 
assign U3500 = U4424 & U4423 & U4422 & U4421; 
assign U3501 = U4428 & U4427 & U4426 & U4425; 
assign U3502 = U4432 & U4431 & U4430 & U4429; 
assign U3503 = U4436 & U4435 & U4434 & U4433; 
assign U3504 = U4407 & U4406 & U4405 & U4404; 
assign U3505 = U4411 & U4410 & U4409 & U4408; 
assign U3506 = U4415 & U4414 & U4413 & U4412; 
assign U3507 = U4419 & U4418 & U4417 & U4416; 
assign U3524 = U4441 & U4440 & U4439 & U4438; 
assign U3525 = U4443 & U4442 & U4444; 
assign U3548 = U4469 & U4468 & U4467 & U4466; 
assign U3549 = U4473 & U4472 & U4471 & U4470; 
assign U3550 = U4477 & U4476 & U4475 & U4474; 
assign U3551 = U4481 & U4480 & U4479 & U4478; 
assign U3552 = U4452 & U4451 & U4450 & U4449; 
assign U3553 = U4456 & U4455 & U4454 & U4453; 
assign U3554 = U4460 & U4459 & U4458 & U4457; 
assign U3555 = U4464 & U4463 & U4462 & U4461; 
assign U3557 = U4407 & U4406 & U4405 & U4404; 
assign U3558 = U4411 & U4410 & U4409 & U4408; 
assign U3559 = U4415 & U4414 & U4413 & U4412; 
assign U3560 = U4419 & U4418 & U4417 & U4416; 
assign U3875 = U4229 & U4232 & U6350; 
assign U4100 = U7206 & U7205; 
assign U4161 = ~(U3564 & U2607 & U3563 & U3562 & U3561); 
assign U4220 = ~U3239; 
assign U4221 = ~U3237; 
assign U4228 = ~(U3951 & U4208); 
assign U4356 = ~(U4347 & U4355 & STATE_REG_0__SCAN_IN); 
assign U4363 = ~(U4362 & U3235); 
assign U4388 = ~U3265; 
assign U4485 = ~U3259; 
assign U4528 = ~U3347; 
assign U4590 = ~U3311; 
assign U4598 = ~(U3311 & STATE2_REG_3__SCAN_IN); 
assign U4648 = ~U3317; 
assign U4657 = ~(U3317 & STATE2_REG_3__SCAN_IN); 
assign U4763 = ~U3328; 
assign U4772 = ~(U3328 & STATE2_REG_3__SCAN_IN); 
assign U4821 = ~U3333; 
assign U4829 = ~(U3333 & STATE2_REG_3__SCAN_IN); 
assign U4878 = ~U3336; 
assign U4887 = ~(U3336 & STATE2_REG_3__SCAN_IN); 
assign U4936 = ~U3340; 
assign U4944 = ~(U3340 & STATE2_REG_3__SCAN_IN); 
assign U5049 = ~U3350; 
assign U5057 = ~(U3350 & STATE2_REG_3__SCAN_IN); 
assign U5106 = ~U3353; 
assign U5115 = ~(U3353 & STATE2_REG_3__SCAN_IN); 
assign U5279 = ~U3364; 
assign U5287 = ~(U3364 & STATE2_REG_3__SCAN_IN); 
assign U5336 = ~U3367; 
assign U5345 = ~(U3367 & STATE2_REG_3__SCAN_IN); 
assign U5471 = ~U3425; 
assign U5522 = ~(U7703 & STATE2_REG_1__SCAN_IN); 
assign U6600 = ~(U4243 & STATE2_REG_0__SCAN_IN); 
assign U6746 = ~(R2337_U54 & U2352); 
assign U6754 = ~(R2337_U56 & U2352); 
assign U6766 = ~(R2337_U57 & U2352); 
assign U7058 = ~(U2577 & INSTQUEUE_REG_12__7__SCAN_IN); 
assign U7059 = ~(U2576 & INSTQUEUE_REG_13__7__SCAN_IN); 
assign U7060 = ~(U2575 & INSTQUEUE_REG_14__7__SCAN_IN); 
assign U7061 = ~(U2574 & INSTQUEUE_REG_15__7__SCAN_IN); 
assign U7085 = ~(U4191 & U3347); 
assign U7090 = ~(U2577 & INSTQUEUE_REG_12__6__SCAN_IN); 
assign U7091 = ~(U2576 & INSTQUEUE_REG_13__6__SCAN_IN); 
assign U7092 = ~(U2575 & INSTQUEUE_REG_14__6__SCAN_IN); 
assign U7093 = ~(U2574 & INSTQUEUE_REG_15__6__SCAN_IN); 
assign U7107 = ~(U2577 & INSTQUEUE_REG_12__5__SCAN_IN); 
assign U7108 = ~(U2576 & INSTQUEUE_REG_13__5__SCAN_IN); 
assign U7109 = ~(U2575 & INSTQUEUE_REG_14__5__SCAN_IN); 
assign U7110 = ~(U2574 & INSTQUEUE_REG_15__5__SCAN_IN); 
assign U7124 = ~(U2577 & INSTQUEUE_REG_12__4__SCAN_IN); 
assign U7125 = ~(U2576 & INSTQUEUE_REG_13__4__SCAN_IN); 
assign U7126 = ~(U2575 & INSTQUEUE_REG_14__4__SCAN_IN); 
assign U7127 = ~(U2574 & INSTQUEUE_REG_15__4__SCAN_IN); 
assign U7139 = ~(U2577 & INSTQUEUE_REG_12__3__SCAN_IN); 
assign U7140 = ~(U2576 & INSTQUEUE_REG_13__3__SCAN_IN); 
assign U7141 = ~(U2575 & INSTQUEUE_REG_14__3__SCAN_IN); 
assign U7142 = ~(U2574 & INSTQUEUE_REG_15__3__SCAN_IN); 
assign U7156 = ~(U2577 & INSTQUEUE_REG_12__2__SCAN_IN); 
assign U7157 = ~(U2576 & INSTQUEUE_REG_13__2__SCAN_IN); 
assign U7158 = ~(U2575 & INSTQUEUE_REG_14__2__SCAN_IN); 
assign U7159 = ~(U2574 & INSTQUEUE_REG_15__2__SCAN_IN); 
assign U7173 = ~(U2577 & INSTQUEUE_REG_12__1__SCAN_IN); 
assign U7174 = ~(U2576 & INSTQUEUE_REG_13__1__SCAN_IN); 
assign U7175 = ~(U2575 & INSTQUEUE_REG_14__1__SCAN_IN); 
assign U7176 = ~(U2574 & INSTQUEUE_REG_15__1__SCAN_IN); 
assign U7190 = ~(U2577 & INSTQUEUE_REG_12__0__SCAN_IN); 
assign U7191 = ~(U2576 & INSTQUEUE_REG_13__0__SCAN_IN); 
assign U7192 = ~(U2575 & INSTQUEUE_REG_14__0__SCAN_IN); 
assign U7193 = ~(U2574 & INSTQUEUE_REG_15__0__SCAN_IN); 
assign U7204 = ~(U4191 & U3442); 
assign U7458 = ~(U4098 & U7206); 
assign U7483 = ~(U4059 & U2607 & U4058 & U4057 & U4056); 
assign U7610 = ~(U7609 & U3248); 
assign U7611 = ~(U4349 & U4346 & STATE_REG_1__SCAN_IN); 
assign U7613 = ~(U4346 & STATE_REG_1__SCAN_IN); 
assign U7631 = ~(U7630 & U7629); 
assign U7632 = ~(U7612 & U4349 & STATE_REG_1__SCAN_IN); 
assign U7684 = ~U3442; 
assign U7735 = ~(U3467 & U4208); 
assign U7741 = ~(U7740 & U7739); 
assign U7745 = ~(U4208 & REIP_REG_1__SCAN_IN); 
assign U7747 = ~(U4208 & U6587); 
assign U7782 = ~(U7703 & STATE2_REG_1__SCAN_IN & FLUSH_REG_SCAN_IN); 
assign R2027_U16 = ~(R2027_U83 & R2027_U112); 
assign R2027_U96 = ~(R2027_U112 & INSTADDRPOINTER_REG_5__SCAN_IN); 
assign R2027_U149 = ~(R2027_U112 & R2027_U12); 
assign R2027_U152 = ~(R2027_U127 & R2027_U8); 
assign R2337_U17 = ~(R2337_U82 & R2337_U110); 
assign R2337_U91 = ~(R2337_U110 & PHYADDRPOINTER_REG_8__SCAN_IN); 
assign R2337_U137 = ~(R2337_U110 & R2337_U14); 
assign R2337_U139 = ~(R2337_U109 & R2337_U11); 
assign R2337_U143 = ~(R2337_U107 & R2337_U6); 
assign R2096_U10 = ~(R2096_U95 & REIP_REG_4__SCAN_IN); 
assign R2096_U134 = ~(R2096_U95 & R2096_U9); 
assign R2238_U32 = ~(R2238_U31 & R2238_U29); 
assign R2238_U65 = ~(R2238_U64 & R2238_U30); 
assign SUB_450_U32 = ~(SUB_450_U31 & SUB_450_U29); 
assign SUB_450_U65 = ~(SUB_450_U64 & SUB_450_U30); 
assign ADD_405_U10 = ~(ADD_405_U98 & INSTADDRPOINTER_REG_4__SCAN_IN); 
assign ADD_405_U93 = ADD_405_U140 & ADD_405_U139; 
assign ADD_405_U138 = ~(ADD_405_U98 & ADD_405_U9); 
assign ADD_515_U10 = ~(ADD_515_U95 & INSTADDRPOINTER_REG_4__SCAN_IN); 
assign ADD_515_U134 = ~(ADD_515_U95 & ADD_515_U9); 
assign U2433 = U4528 & U3442; 
assign U2434 = U7684 & U3347; 
assign U2435 = U4528 & U7684; 
assign U2450 = U4388 & STATE2_REG_0__SCAN_IN; 
assign U2522 = U5471 & U5499; 
assign U2530 = U5471 & U3388; 
assign U2536 = U2535 & U2521; 
assign U2537 = U2535 & U2524; 
assign U2538 = U2535 & U2526; 
assign U2539 = U2535 & U2528; 
assign U2541 = U2521 & U2540; 
assign U2542 = U2524 & U2540; 
assign U2543 = U2526 & U2540; 
assign U2544 = U2528 & U2540; 
assign U2555 = U7708 & U3429; 
assign U2560 = U3443 & U3429; 
assign U2570 = U2569 & U3486; 
assign U2571 = U2569 & U2454; 
assign U2572 = U2569 & U2456; 
assign U2573 = U2569 & U4366; 
assign U2593 = U4172 & U3444; 
assign U2598 = U3444 & U3439; 
assign U2794 = ~(U7745 & U7744 & U4228); 
assign U2795 = ~(U7735 & U7734 & U4228); 
assign U3223 = ~(U2432 & U3222); 
assign U3224 = ~(U2432 & U4531); 
assign U3258 = ~(U3555 & U3554 & U3553 & U3552); 
assign U3263 = ~(U3507 & U3506 & U3505 & U3504); 
assign U3264 = ~(U3527 & U4158 & U3526 & U3525 & U3524); 
assign U3270 = ~(U3499 & U3498 & U3497 & U3496); 
assign U3271 = ~(U3551 & U3550 & U3549 & U3548); 
assign U3378 = ~(U3503 & U3502 & U3501 & U3500); 
assign U3402 = ~(U4388 & U4161); 
assign U3440 = ~(U2605 & STATE2_REG_0__SCAN_IN); 
assign U3469 = ~(U7747 & U7746); 
assign U3482 = U4356 & U3239; 
assign U3721 = U4485 & U3244; 
assign U3993 = U6746 & U6745; 
assign U4052 = U7061 & U7060 & U7059 & U7058; 
assign U4066 = U7085 & U7083; 
assign U4068 = U7093 & U7092 & U7091 & U7090; 
assign U4072 = U7110 & U7109 & U7108 & U7107; 
assign U4076 = U7127 & U7126 & U7125 & U7124; 
assign U4081 = U7142 & U7141 & U7140 & U7139; 
assign U4085 = U7159 & U7158 & U7157 & U7156; 
assign U4089 = U7176 & U7175 & U7174 & U7173; 
assign U4093 = U7193 & U7192 & U7191 & U7190; 
assign U4097 = U7204 & U7203; 
assign U4148 = U4161 & STATE2_REG_0__SCAN_IN; 
assign U4159 = ~(U3560 & U3559 & U3558 & U3557); 
assign U4255 = ~(U4221 & REIP_REG_31__SCAN_IN); 
assign U4256 = ~(U4220 & REIP_REG_30__SCAN_IN); 
assign U4258 = ~(U4221 & REIP_REG_30__SCAN_IN); 
assign U4259 = ~(U4220 & REIP_REG_29__SCAN_IN); 
assign U4261 = ~(U4221 & REIP_REG_29__SCAN_IN); 
assign U4262 = ~(U4220 & REIP_REG_28__SCAN_IN); 
assign U4264 = ~(U4221 & REIP_REG_28__SCAN_IN); 
assign U4265 = ~(U4220 & REIP_REG_27__SCAN_IN); 
assign U4267 = ~(U4221 & REIP_REG_27__SCAN_IN); 
assign U4268 = ~(U4220 & REIP_REG_26__SCAN_IN); 
assign U4270 = ~(U4221 & REIP_REG_26__SCAN_IN); 
assign U4271 = ~(U4220 & REIP_REG_25__SCAN_IN); 
assign U4273 = ~(U4221 & REIP_REG_25__SCAN_IN); 
assign U4274 = ~(U4220 & REIP_REG_24__SCAN_IN); 
assign U4276 = ~(U4221 & REIP_REG_24__SCAN_IN); 
assign U4277 = ~(U4220 & REIP_REG_23__SCAN_IN); 
assign U4279 = ~(U4221 & REIP_REG_23__SCAN_IN); 
assign U4280 = ~(U4220 & REIP_REG_22__SCAN_IN); 
assign U4282 = ~(U4221 & REIP_REG_22__SCAN_IN); 
assign U4283 = ~(U4220 & REIP_REG_21__SCAN_IN); 
assign U4285 = ~(U4221 & REIP_REG_21__SCAN_IN); 
assign U4286 = ~(U4220 & REIP_REG_20__SCAN_IN); 
assign U4288 = ~(U4221 & REIP_REG_20__SCAN_IN); 
assign U4289 = ~(U4220 & REIP_REG_19__SCAN_IN); 
assign U4291 = ~(U4221 & REIP_REG_19__SCAN_IN); 
assign U4292 = ~(U4220 & REIP_REG_18__SCAN_IN); 
assign U4294 = ~(U4221 & REIP_REG_18__SCAN_IN); 
assign U4295 = ~(U4220 & REIP_REG_17__SCAN_IN); 
assign U4297 = ~(U4221 & REIP_REG_17__SCAN_IN); 
assign U4298 = ~(U4220 & REIP_REG_16__SCAN_IN); 
assign U4300 = ~(U4221 & REIP_REG_16__SCAN_IN); 
assign U4301 = ~(U4220 & REIP_REG_15__SCAN_IN); 
assign U4303 = ~(U4221 & REIP_REG_15__SCAN_IN); 
assign U4304 = ~(U4220 & REIP_REG_14__SCAN_IN); 
assign U4306 = ~(U4221 & REIP_REG_14__SCAN_IN); 
assign U4307 = ~(U4220 & REIP_REG_13__SCAN_IN); 
assign U4309 = ~(U4221 & REIP_REG_13__SCAN_IN); 
assign U4310 = ~(U4220 & REIP_REG_12__SCAN_IN); 
assign U4312 = ~(U4221 & REIP_REG_12__SCAN_IN); 
assign U4313 = ~(U4220 & REIP_REG_11__SCAN_IN); 
assign U4315 = ~(U4221 & REIP_REG_11__SCAN_IN); 
assign U4316 = ~(U4220 & REIP_REG_10__SCAN_IN); 
assign U4318 = ~(U4221 & REIP_REG_10__SCAN_IN); 
assign U4319 = ~(U4220 & REIP_REG_9__SCAN_IN); 
assign U4321 = ~(U4221 & REIP_REG_9__SCAN_IN); 
assign U4322 = ~(U4220 & REIP_REG_8__SCAN_IN); 
assign U4324 = ~(U4221 & REIP_REG_8__SCAN_IN); 
assign U4325 = ~(U4220 & REIP_REG_7__SCAN_IN); 
assign U4327 = ~(U4221 & REIP_REG_7__SCAN_IN); 
assign U4328 = ~(U4220 & REIP_REG_6__SCAN_IN); 
assign U4330 = ~(U4221 & REIP_REG_6__SCAN_IN); 
assign U4331 = ~(U4220 & REIP_REG_5__SCAN_IN); 
assign U4333 = ~(U4221 & REIP_REG_5__SCAN_IN); 
assign U4334 = ~(U4220 & REIP_REG_4__SCAN_IN); 
assign U4336 = ~(U4221 & REIP_REG_4__SCAN_IN); 
assign U4337 = ~(U4220 & REIP_REG_3__SCAN_IN); 
assign U4339 = ~(U4221 & REIP_REG_3__SCAN_IN); 
assign U4340 = ~(U4220 & REIP_REG_2__SCAN_IN); 
assign U4342 = ~(U4221 & REIP_REG_2__SCAN_IN); 
assign U4343 = ~(U4220 & REIP_REG_1__SCAN_IN); 
assign U4351 = ~(U7610 & U4350 & U7611); 
assign U4359 = ~(U3484 & U7613); 
assign U4403 = ~U4161; 
assign U4532 = ~(U2432 & U2436); 
assign U4651 = ~(U2437 & U2432); 
assign U5468 = ~U3429; 
assign U5476 = ~(U4388 & U2605); 
assign U5503 = ~(U2446 & U3457); 
assign U6592 = ~(U4485 & STATEBS16_REG_SCAN_IN); 
assign U7054 = ~(U2582 & INSTQUEUE_REG_8__7__SCAN_IN); 
assign U7055 = ~(U2581 & INSTQUEUE_REG_9__7__SCAN_IN); 
assign U7056 = ~(U2580 & INSTQUEUE_REG_10__7__SCAN_IN); 
assign U7057 = ~(U2579 & INSTQUEUE_REG_11__7__SCAN_IN); 
assign U7066 = ~(U2568 & INSTQUEUE_REG_4__7__SCAN_IN); 
assign U7067 = ~(U2567 & INSTQUEUE_REG_5__7__SCAN_IN); 
assign U7068 = ~(U2566 & INSTQUEUE_REG_6__7__SCAN_IN); 
assign U7069 = ~(U2565 & INSTQUEUE_REG_7__7__SCAN_IN); 
assign U7086 = ~(U2582 & INSTQUEUE_REG_8__6__SCAN_IN); 
assign U7087 = ~(U2581 & INSTQUEUE_REG_9__6__SCAN_IN); 
assign U7088 = ~(U2580 & INSTQUEUE_REG_10__6__SCAN_IN); 
assign U7089 = ~(U2579 & INSTQUEUE_REG_11__6__SCAN_IN); 
assign U7098 = ~(U2568 & INSTQUEUE_REG_4__6__SCAN_IN); 
assign U7099 = ~(U2567 & INSTQUEUE_REG_5__6__SCAN_IN); 
assign U7100 = ~(U2566 & INSTQUEUE_REG_6__6__SCAN_IN); 
assign U7101 = ~(U2565 & INSTQUEUE_REG_7__6__SCAN_IN); 
assign U7103 = ~(U2582 & INSTQUEUE_REG_8__5__SCAN_IN); 
assign U7104 = ~(U2581 & INSTQUEUE_REG_9__5__SCAN_IN); 
assign U7105 = ~(U2580 & INSTQUEUE_REG_10__5__SCAN_IN); 
assign U7106 = ~(U2579 & INSTQUEUE_REG_11__5__SCAN_IN); 
assign U7115 = ~(U2568 & INSTQUEUE_REG_4__5__SCAN_IN); 
assign U7116 = ~(U2567 & INSTQUEUE_REG_5__5__SCAN_IN); 
assign U7117 = ~(U2566 & INSTQUEUE_REG_6__5__SCAN_IN); 
assign U7118 = ~(U2565 & INSTQUEUE_REG_7__5__SCAN_IN); 
assign U7120 = ~(U2582 & INSTQUEUE_REG_8__4__SCAN_IN); 
assign U7121 = ~(U2581 & INSTQUEUE_REG_9__4__SCAN_IN); 
assign U7122 = ~(U2580 & INSTQUEUE_REG_10__4__SCAN_IN); 
assign U7123 = ~(U2579 & INSTQUEUE_REG_11__4__SCAN_IN); 
assign U7131 = ~(U2568 & INSTQUEUE_REG_4__4__SCAN_IN); 
assign U7132 = ~(U2567 & INSTQUEUE_REG_5__4__SCAN_IN); 
assign U7133 = ~(U2566 & INSTQUEUE_REG_6__4__SCAN_IN); 
assign U7134 = ~(U2565 & INSTQUEUE_REG_7__4__SCAN_IN); 
assign U7135 = ~(U2582 & INSTQUEUE_REG_8__3__SCAN_IN); 
assign U7136 = ~(U2581 & INSTQUEUE_REG_9__3__SCAN_IN); 
assign U7137 = ~(U2580 & INSTQUEUE_REG_10__3__SCAN_IN); 
assign U7138 = ~(U2579 & INSTQUEUE_REG_11__3__SCAN_IN); 
assign U7147 = ~(U2568 & INSTQUEUE_REG_4__3__SCAN_IN); 
assign U7148 = ~(U2567 & INSTQUEUE_REG_5__3__SCAN_IN); 
assign U7149 = ~(U2566 & INSTQUEUE_REG_6__3__SCAN_IN); 
assign U7150 = ~(U2565 & INSTQUEUE_REG_7__3__SCAN_IN); 
assign U7152 = ~(U2582 & INSTQUEUE_REG_8__2__SCAN_IN); 
assign U7153 = ~(U2581 & INSTQUEUE_REG_9__2__SCAN_IN); 
assign U7154 = ~(U2580 & INSTQUEUE_REG_10__2__SCAN_IN); 
assign U7155 = ~(U2579 & INSTQUEUE_REG_11__2__SCAN_IN); 
assign U7164 = ~(U2568 & INSTQUEUE_REG_4__2__SCAN_IN); 
assign U7165 = ~(U2567 & INSTQUEUE_REG_5__2__SCAN_IN); 
assign U7166 = ~(U2566 & INSTQUEUE_REG_6__2__SCAN_IN); 
assign U7167 = ~(U2565 & INSTQUEUE_REG_7__2__SCAN_IN); 
assign U7169 = ~(U2582 & INSTQUEUE_REG_8__1__SCAN_IN); 
assign U7170 = ~(U2581 & INSTQUEUE_REG_9__1__SCAN_IN); 
assign U7171 = ~(U2580 & INSTQUEUE_REG_10__1__SCAN_IN); 
assign U7172 = ~(U2579 & INSTQUEUE_REG_11__1__SCAN_IN); 
assign U7181 = ~(U2568 & INSTQUEUE_REG_4__1__SCAN_IN); 
assign U7182 = ~(U2567 & INSTQUEUE_REG_5__1__SCAN_IN); 
assign U7183 = ~(U2566 & INSTQUEUE_REG_6__1__SCAN_IN); 
assign U7184 = ~(U2565 & INSTQUEUE_REG_7__1__SCAN_IN); 
assign U7186 = ~(U2582 & INSTQUEUE_REG_8__0__SCAN_IN); 
assign U7187 = ~(U2581 & INSTQUEUE_REG_9__0__SCAN_IN); 
assign U7188 = ~(U2580 & INSTQUEUE_REG_10__0__SCAN_IN); 
assign U7189 = ~(U2579 & INSTQUEUE_REG_11__0__SCAN_IN); 
assign U7198 = ~(U2568 & INSTQUEUE_REG_4__0__SCAN_IN); 
assign U7199 = ~(U2567 & INSTQUEUE_REG_5__0__SCAN_IN); 
assign U7200 = ~(U2566 & INSTQUEUE_REG_6__0__SCAN_IN); 
assign U7201 = ~(U2565 & INSTQUEUE_REG_7__0__SCAN_IN); 
assign U7368 = ~(U4161 & STATE2_REG_0__SCAN_IN); 
assign U7449 = ~(U2446 & U3457 & FLUSH_REG_SCAN_IN); 
assign U7466 = ~(U2608 & U3253); 
assign U7479 = ~(U4096 & U7204); 
assign U7633 = ~(U7631 & U3235); 
assign U7638 = ~U3449; 
assign U7640 = ~(U3450 & U3449); 
assign U7641 = ~(U3449 & U4364); 
assign U7700 = ~U3457; 
assign U7743 = ~(U7741 & U4208); 
assign U7753 = ~(BS16_N & U3449); 
assign U7778 = ~U3444; 
assign R2027_U55 = ~(R2027_U150 & R2027_U149); 
assign R2027_U56 = ~(R2027_U152 & R2027_U151); 
assign R2027_U118 = ~R2027_U16; 
assign R2027_U126 = ~R2027_U96; 
assign R2027_U146 = ~(R2027_U16 & INSTADDRPOINTER_REG_7__SCAN_IN); 
assign R2027_U147 = ~(R2027_U96 & INSTADDRPOINTER_REG_6__SCAN_IN); 
assign R2337_U52 = ~(R2337_U137 & R2337_U136); 
assign R2337_U53 = ~(R2337_U139 & R2337_U138); 
assign R2337_U55 = ~(R2337_U143 & R2337_U142); 
assign R2337_U111 = ~R2337_U91; 
assign R2337_U112 = ~R2337_U17; 
assign R2337_U134 = ~(R2337_U91 & PHYADDRPOINTER_REG_9__SCAN_IN); 
assign R2337_U192 = ~(R2337_U17 & PHYADDRPOINTER_REG_10__SCAN_IN); 
assign R2096_U67 = ~(R2096_U134 & R2096_U133); 
assign R2096_U96 = ~R2096_U10; 
assign R2096_U131 = ~(R2096_U10 & REIP_REG_5__SCAN_IN); 
assign R2238_U22 = ~(R2238_U66 & R2238_U65); 
assign R2238_U28 = ~(R2238_U33 & R2238_U32); 
assign SUB_450_U22 = ~(SUB_450_U66 & SUB_450_U65); 
assign SUB_450_U28 = ~(SUB_450_U33 & SUB_450_U32); 
assign ADD_405_U68 = ~(ADD_405_U138 & ADD_405_U137); 
assign ADD_405_U99 = ~ADD_405_U10; 
assign ADD_405_U135 = ~(ADD_405_U10 & INSTADDRPOINTER_REG_5__SCAN_IN); 
assign ADD_515_U67 = ~(ADD_515_U134 & ADD_515_U133); 
assign ADD_515_U96 = ~ADD_515_U10; 
assign ADD_515_U131 = ~(ADD_515_U10 & INSTADDRPOINTER_REG_5__SCAN_IN); 
assign U2452 = U4388 & U3264 & U3378 & U4161; 
assign U2523 = U2522 & U2521; 
assign U2525 = U2522 & U2524; 
assign U2527 = U2522 & U2526; 
assign U2529 = U2522 & U2528; 
assign U2531 = U2530 & U2521; 
assign U2532 = U2530 & U2524; 
assign U2533 = U2530 & U2526; 
assign U2534 = U2530 & U2528; 
assign U2545 = U5468 & U7708; 
assign U2550 = U5468 & U3443; 
assign U2556 = U2555 & U2454; 
assign U2557 = U2555 & U3486; 
assign U2558 = U2555 & U4366; 
assign U2559 = U2555 & U2456; 
assign U2561 = U2560 & U2454; 
assign U2562 = U2560 & U3486; 
assign U2563 = U2560 & U4366; 
assign U2564 = U2560 & U2456; 
assign U2583 = U7778 & U4172; 
assign U2588 = U7778 & U3439; 
assign U2594 = U2593 & U2524; 
assign U2595 = U2593 & U2521; 
assign U2596 = U2593 & U2528; 
assign U2597 = U2593 & U2526; 
assign U2599 = U2598 & U2524; 
assign U2600 = U2598 & U2521; 
assign U2601 = U2598 & U2528; 
assign U2602 = U2598 & U2526; 
assign U2789 = ~(U7638 & U6601); 
assign U3151 = U7638 & DATAWIDTH_REG_31__SCAN_IN; 
assign U3152 = U7638 & DATAWIDTH_REG_30__SCAN_IN; 
assign U3153 = U7638 & DATAWIDTH_REG_29__SCAN_IN; 
assign U3154 = U7638 & DATAWIDTH_REG_28__SCAN_IN; 
assign U3155 = U7638 & DATAWIDTH_REG_27__SCAN_IN; 
assign U3156 = U7638 & DATAWIDTH_REG_26__SCAN_IN; 
assign U3157 = U7638 & DATAWIDTH_REG_25__SCAN_IN; 
assign U3158 = U7638 & DATAWIDTH_REG_24__SCAN_IN; 
assign U3159 = U7638 & DATAWIDTH_REG_23__SCAN_IN; 
assign U3160 = U7638 & DATAWIDTH_REG_22__SCAN_IN; 
assign U3161 = U7638 & DATAWIDTH_REG_21__SCAN_IN; 
assign U3162 = U7638 & DATAWIDTH_REG_20__SCAN_IN; 
assign U3163 = U7638 & DATAWIDTH_REG_19__SCAN_IN; 
assign U3164 = U7638 & DATAWIDTH_REG_18__SCAN_IN; 
assign U3165 = U7638 & DATAWIDTH_REG_17__SCAN_IN; 
assign U3166 = U7638 & DATAWIDTH_REG_16__SCAN_IN; 
assign U3167 = U7638 & DATAWIDTH_REG_15__SCAN_IN; 
assign U3168 = U7638 & DATAWIDTH_REG_14__SCAN_IN; 
assign U3169 = U7638 & DATAWIDTH_REG_13__SCAN_IN; 
assign U3170 = U7638 & DATAWIDTH_REG_12__SCAN_IN; 
assign U3171 = U7638 & DATAWIDTH_REG_11__SCAN_IN; 
assign U3172 = U7638 & DATAWIDTH_REG_10__SCAN_IN; 
assign U3173 = U7638 & DATAWIDTH_REG_9__SCAN_IN; 
assign U3174 = U7638 & DATAWIDTH_REG_8__SCAN_IN; 
assign U3175 = U7638 & DATAWIDTH_REG_7__SCAN_IN; 
assign U3176 = U7638 & DATAWIDTH_REG_6__SCAN_IN; 
assign U3177 = U7638 & DATAWIDTH_REG_5__SCAN_IN; 
assign U3178 = U7638 & DATAWIDTH_REG_4__SCAN_IN; 
assign U3179 = U7638 & DATAWIDTH_REG_3__SCAN_IN; 
assign U3180 = U7638 & DATAWIDTH_REG_2__SCAN_IN; 
assign U3182 = ~(U7633 & U7632 & U3483); 
assign U3184 = ~(U4343 & U4342 & U4344); 
assign U3185 = ~(U4340 & U4339 & U4341); 
assign U3186 = ~(U4337 & U4336 & U4338); 
assign U3187 = ~(U4334 & U4333 & U4335); 
assign U3188 = ~(U4331 & U4330 & U4332); 
assign U3189 = ~(U4328 & U4327 & U4329); 
assign U3190 = ~(U4325 & U4324 & U4326); 
assign U3191 = ~(U4322 & U4321 & U4323); 
assign U3192 = ~(U4319 & U4318 & U4320); 
assign U3193 = ~(U4316 & U4315 & U4317); 
assign U3194 = ~(U4313 & U4312 & U4314); 
assign U3195 = ~(U4310 & U4309 & U4311); 
assign U3196 = ~(U4307 & U4306 & U4308); 
assign U3197 = ~(U4304 & U4303 & U4305); 
assign U3198 = ~(U4301 & U4300 & U4302); 
assign U3199 = ~(U4298 & U4297 & U4299); 
assign U3200 = ~(U4295 & U4294 & U4296); 
assign U3201 = ~(U4292 & U4291 & U4293); 
assign U3202 = ~(U4289 & U4288 & U4290); 
assign U3203 = ~(U4286 & U4285 & U4287); 
assign U3204 = ~(U4283 & U4282 & U4284); 
assign U3205 = ~(U4280 & U4279 & U4281); 
assign U3206 = ~(U4277 & U4276 & U4278); 
assign U3207 = ~(U4274 & U4273 & U4275); 
assign U3208 = ~(U4271 & U4270 & U4272); 
assign U3209 = ~(U4268 & U4267 & U4269); 
assign U3210 = ~(U4265 & U4264 & U4266); 
assign U3211 = ~(U4262 & U4261 & U4263); 
assign U3212 = ~(U4259 & U4258 & U4260); 
assign U3213 = ~(U4256 & U4255 & U4257); 
assign U3225 = ~(U2434 & U3222); 
assign U3226 = ~(U2434 & U4531); 
assign U3227 = ~(U2433 & U3222); 
assign U3228 = ~(U2433 & U4531); 
assign U3229 = ~(U2435 & U3222); 
assign U3230 = ~(U2435 & U4531); 
assign U3277 = ~(U3258 & U3270); 
assign U3309 = ~(U3293 & U4532); 
assign U3323 = ~(U3317 & U4651); 
assign U3376 = ~(U3271 & U3265); 
assign U3377 = ~(U3271 & U3258); 
assign U3381 = ~(U2605 & U3264); 
assign U3392 = ~(U3265 & U3271 & STATE2_REG_0__SCAN_IN); 
assign U3394 = ~(U3264 & U3378); 
assign U3399 = ~(U3258 & STATE2_REG_2__SCAN_IN); 
assign U3468 = ~(U7743 & U7742); 
assign U3853 = U2368 & U3271; 
assign U3872 = U2605 & U3378; 
assign U4051 = U7057 & U7056 & U7055 & U7054; 
assign U4054 = U7069 & U7068 & U7067 & U7066; 
assign U4060 = U4388 & U3378; 
assign U4061 = U3271 & STATE2_REG_0__SCAN_IN; 
assign U4067 = U7089 & U7088 & U7087 & U7086; 
assign U4070 = U7101 & U7100 & U7099 & U7098; 
assign U4071 = U7106 & U7105 & U7104 & U7103; 
assign U4074 = U7118 & U7117 & U7116 & U7115; 
assign U4075 = U7123 & U7122 & U7121 & U7120; 
assign U4078 = U7133 & U7132; 
assign U4080 = U7138 & U7137 & U7136 & U7135; 
assign U4083 = U7150 & U7149 & U7148 & U7147; 
assign U4084 = U7155 & U7154 & U7153 & U7152; 
assign U4087 = U7167 & U7166 & U7165 & U7164; 
assign U4088 = U7172 & U7171 & U7170 & U7169; 
assign U4091 = U7184 & U7183 & U7182 & U7181; 
assign U4092 = U7189 & U7188 & U7187 & U7186; 
assign U4095 = U7201 & U7200 & U7199 & U7198; 
assign U4142 = U3270 & U3378; 
assign U4147 = U3258 & U4161; 
assign U4156 = U7450 & U7449; 
assign U4239 = ~U3402; 
assign U4253 = ~U3440; 
assign U4357 = ~(U4351 & STATE_REG_2__SCAN_IN); 
assign U4387 = ~U3270; 
assign U4420 = ~U4159; 
assign U4437 = ~U3378; 
assign U4448 = ~U3264; 
assign U4465 = ~U3258; 
assign U4482 = ~U3271; 
assign U4593 = ~U3223; 
assign U4599 = ~(U3223 & STATE2_REG_2__SCAN_IN); 
assign U4709 = ~U3224; 
assign U4715 = ~(U3224 & STATE2_REG_2__SCAN_IN); 
assign U4766 = ~(U2434 & U2436); 
assign U4881 = ~(U2434 & U2437); 
assign U4995 = ~(U2433 & U2436); 
assign U5109 = ~(U2433 & U2437); 
assign U5224 = ~(U2435 & U2436); 
assign U5339 = ~(U2435 & U2437); 
assign U5514 = ~(U7700 & U2446); 
assign U6606 = ~(U2544 & INSTQUEUE_REG_15__7__SCAN_IN); 
assign U6607 = ~(U2543 & INSTQUEUE_REG_14__7__SCAN_IN); 
assign U6608 = ~(U2542 & INSTQUEUE_REG_13__7__SCAN_IN); 
assign U6609 = ~(U2541 & INSTQUEUE_REG_12__7__SCAN_IN); 
assign U6610 = ~(U2539 & INSTQUEUE_REG_11__7__SCAN_IN); 
assign U6611 = ~(U2538 & INSTQUEUE_REG_10__7__SCAN_IN); 
assign U6612 = ~(U2537 & INSTQUEUE_REG_9__7__SCAN_IN); 
assign U6613 = ~(U2536 & INSTQUEUE_REG_8__7__SCAN_IN); 
assign U6622 = ~(U2544 & INSTQUEUE_REG_15__6__SCAN_IN); 
assign U6623 = ~(U2543 & INSTQUEUE_REG_14__6__SCAN_IN); 
assign U6624 = ~(U2542 & INSTQUEUE_REG_13__6__SCAN_IN); 
assign U6625 = ~(U2541 & INSTQUEUE_REG_12__6__SCAN_IN); 
assign U6626 = ~(U2539 & INSTQUEUE_REG_11__6__SCAN_IN); 
assign U6627 = ~(U2538 & INSTQUEUE_REG_10__6__SCAN_IN); 
assign U6628 = ~(U2537 & INSTQUEUE_REG_9__6__SCAN_IN); 
assign U6629 = ~(U2536 & INSTQUEUE_REG_8__6__SCAN_IN); 
assign U6638 = ~(U2544 & INSTQUEUE_REG_15__5__SCAN_IN); 
assign U6639 = ~(U2543 & INSTQUEUE_REG_14__5__SCAN_IN); 
assign U6640 = ~(U2542 & INSTQUEUE_REG_13__5__SCAN_IN); 
assign U6641 = ~(U2541 & INSTQUEUE_REG_12__5__SCAN_IN); 
assign U6642 = ~(U2539 & INSTQUEUE_REG_11__5__SCAN_IN); 
assign U6643 = ~(U2538 & INSTQUEUE_REG_10__5__SCAN_IN); 
assign U6644 = ~(U2537 & INSTQUEUE_REG_9__5__SCAN_IN); 
assign U6645 = ~(U2536 & INSTQUEUE_REG_8__5__SCAN_IN); 
assign U6654 = ~(U2544 & INSTQUEUE_REG_15__4__SCAN_IN); 
assign U6655 = ~(U2543 & INSTQUEUE_REG_14__4__SCAN_IN); 
assign U6656 = ~(U2542 & INSTQUEUE_REG_13__4__SCAN_IN); 
assign U6657 = ~(U2541 & INSTQUEUE_REG_12__4__SCAN_IN); 
assign U6658 = ~(U2539 & INSTQUEUE_REG_11__4__SCAN_IN); 
assign U6659 = ~(U2538 & INSTQUEUE_REG_10__4__SCAN_IN); 
assign U6660 = ~(U2537 & INSTQUEUE_REG_9__4__SCAN_IN); 
assign U6661 = ~(U2536 & INSTQUEUE_REG_8__4__SCAN_IN); 
assign U6669 = ~(U2544 & INSTQUEUE_REG_15__3__SCAN_IN); 
assign U6670 = ~(U2543 & INSTQUEUE_REG_14__3__SCAN_IN); 
assign U6671 = ~(U2542 & INSTQUEUE_REG_13__3__SCAN_IN); 
assign U6672 = ~(U2541 & INSTQUEUE_REG_12__3__SCAN_IN); 
assign U6673 = ~(U2539 & INSTQUEUE_REG_11__3__SCAN_IN); 
assign U6674 = ~(U2538 & INSTQUEUE_REG_10__3__SCAN_IN); 
assign U6675 = ~(U2537 & INSTQUEUE_REG_9__3__SCAN_IN); 
assign U6676 = ~(U2536 & INSTQUEUE_REG_8__3__SCAN_IN); 
assign U6685 = ~(U2544 & INSTQUEUE_REG_15__2__SCAN_IN); 
assign U6686 = ~(U2543 & INSTQUEUE_REG_14__2__SCAN_IN); 
assign U6687 = ~(U2542 & INSTQUEUE_REG_13__2__SCAN_IN); 
assign U6688 = ~(U2541 & INSTQUEUE_REG_12__2__SCAN_IN); 
assign U6689 = ~(U2539 & INSTQUEUE_REG_11__2__SCAN_IN); 
assign U6690 = ~(U2538 & INSTQUEUE_REG_10__2__SCAN_IN); 
assign U6691 = ~(U2537 & INSTQUEUE_REG_9__2__SCAN_IN); 
assign U6692 = ~(U2536 & INSTQUEUE_REG_8__2__SCAN_IN); 
assign U6701 = ~(U2544 & INSTQUEUE_REG_15__1__SCAN_IN); 
assign U6702 = ~(U2543 & INSTQUEUE_REG_14__1__SCAN_IN); 
assign U6703 = ~(U2542 & INSTQUEUE_REG_13__1__SCAN_IN); 
assign U6704 = ~(U2541 & INSTQUEUE_REG_12__1__SCAN_IN); 
assign U6705 = ~(U2539 & INSTQUEUE_REG_11__1__SCAN_IN); 
assign U6706 = ~(U2538 & INSTQUEUE_REG_10__1__SCAN_IN); 
assign U6707 = ~(U2537 & INSTQUEUE_REG_9__1__SCAN_IN); 
assign U6708 = ~(U2536 & INSTQUEUE_REG_8__1__SCAN_IN); 
assign U6717 = ~(U2544 & INSTQUEUE_REG_15__0__SCAN_IN); 
assign U6718 = ~(U2543 & INSTQUEUE_REG_14__0__SCAN_IN); 
assign U6719 = ~(U2542 & INSTQUEUE_REG_13__0__SCAN_IN); 
assign U6720 = ~(U2541 & INSTQUEUE_REG_12__0__SCAN_IN); 
assign U6721 = ~(U2539 & INSTQUEUE_REG_11__0__SCAN_IN); 
assign U6722 = ~(U2538 & INSTQUEUE_REG_10__0__SCAN_IN); 
assign U6723 = ~(U2537 & INSTQUEUE_REG_9__0__SCAN_IN); 
assign U6724 = ~(U2536 & INSTQUEUE_REG_8__0__SCAN_IN); 
assign U6740 = ~(R2337_U52 & U2352); 
assign U6743 = ~(R2337_U53 & U2352); 
assign U6750 = ~(R2337_U55 & U2352); 
assign U6876 = ~(U2605 & U3271); 
assign U7062 = ~(U2573 & INSTQUEUE_REG_0__7__SCAN_IN); 
assign U7063 = ~(U2572 & INSTQUEUE_REG_1__7__SCAN_IN); 
assign U7064 = ~(U2571 & INSTQUEUE_REG_2__7__SCAN_IN); 
assign U7065 = ~(U2570 & INSTQUEUE_REG_3__7__SCAN_IN); 
assign U7094 = ~(U2573 & INSTQUEUE_REG_0__6__SCAN_IN); 
assign U7095 = ~(U2572 & INSTQUEUE_REG_1__6__SCAN_IN); 
assign U7096 = ~(U2571 & INSTQUEUE_REG_2__6__SCAN_IN); 
assign U7097 = ~(U2570 & INSTQUEUE_REG_3__6__SCAN_IN); 
assign U7111 = ~(U2573 & INSTQUEUE_REG_0__5__SCAN_IN); 
assign U7112 = ~(U2572 & INSTQUEUE_REG_1__5__SCAN_IN); 
assign U7113 = ~(U2571 & INSTQUEUE_REG_2__5__SCAN_IN); 
assign U7114 = ~(U2570 & INSTQUEUE_REG_3__5__SCAN_IN); 
assign U7128 = ~(U2572 & INSTQUEUE_REG_1__4__SCAN_IN); 
assign U7129 = ~(U2571 & INSTQUEUE_REG_2__4__SCAN_IN); 
assign U7130 = ~(U2570 & INSTQUEUE_REG_3__4__SCAN_IN); 
assign U7143 = ~(U2573 & INSTQUEUE_REG_0__3__SCAN_IN); 
assign U7144 = ~(U2572 & INSTQUEUE_REG_1__3__SCAN_IN); 
assign U7145 = ~(U2571 & INSTQUEUE_REG_2__3__SCAN_IN); 
assign U7146 = ~(U2570 & INSTQUEUE_REG_3__3__SCAN_IN); 
assign U7160 = ~(U2573 & INSTQUEUE_REG_0__2__SCAN_IN); 
assign U7161 = ~(U2572 & INSTQUEUE_REG_1__2__SCAN_IN); 
assign U7162 = ~(U2571 & INSTQUEUE_REG_2__2__SCAN_IN); 
assign U7163 = ~(U2570 & INSTQUEUE_REG_3__2__SCAN_IN); 
assign U7177 = ~(U2573 & INSTQUEUE_REG_0__1__SCAN_IN); 
assign U7178 = ~(U2572 & INSTQUEUE_REG_1__1__SCAN_IN); 
assign U7179 = ~(U2571 & INSTQUEUE_REG_2__1__SCAN_IN); 
assign U7180 = ~(U2570 & INSTQUEUE_REG_3__1__SCAN_IN); 
assign U7194 = ~(U2573 & INSTQUEUE_REG_0__0__SCAN_IN); 
assign U7195 = ~(U2572 & INSTQUEUE_REG_1__0__SCAN_IN); 
assign U7196 = ~(U2571 & INSTQUEUE_REG_2__0__SCAN_IN); 
assign U7197 = ~(U2570 & INSTQUEUE_REG_3__0__SCAN_IN); 
assign U7372 = ~(U2450 & U3258); 
assign U7452 = ~(U2446 & U7700 & FLUSH_REG_SCAN_IN); 
assign U7482 = ~U3263; 
assign U7605 = ~(U2573 & INSTQUEUE_REG_0__4__SCAN_IN); 
assign U7635 = ~(U4359 & U3238); 
assign U7639 = ~(U7638 & DATAWIDTH_REG_0__SCAN_IN); 
assign U7642 = ~(U7638 & DATAWIDTH_REG_1__SCAN_IN); 
assign U7692 = ~(U4403 & U3264); 
assign U7693 = ~(U3258 & U3402); 
assign U7752 = ~(U7638 & STATEBS16_REG_SCAN_IN); 
assign U7772 = ~(U2605 & U3264); 
assign U7779 = ~(U3263 & U3271); 
assign R2027_U17 = ~(R2027_U84 & R2027_U118); 
assign R2027_U95 = ~(R2027_U118 & INSTADDRPOINTER_REG_7__SCAN_IN); 
assign R2027_U145 = ~(R2027_U118 & R2027_U15); 
assign R2027_U148 = ~(R2027_U126 & R2027_U11); 
assign R2337_U20 = ~(R2337_U83 & R2337_U112); 
assign R2337_U104 = ~(R2337_U112 & PHYADDRPOINTER_REG_10__SCAN_IN); 
assign R2337_U135 = ~(R2337_U111 & R2337_U15); 
assign R2337_U193 = ~(R2337_U112 & R2337_U19); 
assign R2096_U12 = ~(R2096_U96 & REIP_REG_5__SCAN_IN); 
assign R2096_U132 = ~(R2096_U96 & R2096_U11); 
assign R2238_U34 = ~R2238_U28; 
assign R2238_U36 = ~(R2238_U35 & R2238_U28); 
assign R2238_U61 = ~(R2238_U25 & R2238_U28); 
assign SUB_450_U34 = ~SUB_450_U28; 
assign SUB_450_U36 = ~(SUB_450_U35 & SUB_450_U28); 
assign SUB_450_U61 = ~(SUB_450_U25 & SUB_450_U28); 
assign ADD_405_U12 = ~(ADD_405_U99 & INSTADDRPOINTER_REG_5__SCAN_IN); 
assign ADD_405_U136 = ~(ADD_405_U99 & ADD_405_U11); 
assign ADD_515_U12 = ~(ADD_515_U96 & INSTADDRPOINTER_REG_5__SCAN_IN); 
assign ADD_515_U132 = ~(ADD_515_U96 & ADD_515_U11); 
assign U2354 = U4253 & U4465; 
assign U2389 = U2452 & U7482; 
assign U2449 = U4482 & U3258; 
assign U2451 = U4239 & STATE2_REG_0__SCAN_IN; 
assign U2546 = U2545 & U2454; 
assign U2547 = U2545 & U3486; 
assign U2548 = U2545 & U4366; 
assign U2549 = U2545 & U2456; 
assign U2551 = U2550 & U2454; 
assign U2552 = U2550 & U3486; 
assign U2553 = U2550 & U4366; 
assign U2554 = U2550 & U2456; 
assign U2584 = U2583 & U2524; 
assign U2585 = U2583 & U2521; 
assign U2586 = U2583 & U2528; 
assign U2587 = U2583 & U2526; 
assign U2589 = U2588 & U2524; 
assign U2590 = U2588 & U2521; 
assign U2591 = U2588 & U2528; 
assign U2592 = U2588 & U2526; 
assign U2603 = U3376 & STATE2_REG_0__SCAN_IN; 
assign U2792 = ~(U7753 & U7752 & U4231); 
assign U3181 = ~(U7635 & U7634 & U4363); 
assign U3183 = ~(U3482 & U4357); 
assign U3269 = ~(U4465 & U3271); 
assign U3274 = ~(U4482 & U4465); 
assign U3276 = ~(U4448 & U3378 & U4161 & U3265); 
assign U3332 = ~(U3328 & U4766); 
assign U3339 = ~(U3336 & U4881); 
assign U3349 = ~(U3343 & U4995); 
assign U3356 = ~(U3353 & U5109); 
assign U3363 = ~(U3360 & U5224); 
assign U3370 = ~(U3367 & U5339); 
assign U3380 = ~(U4387 & U3271); 
assign U3382 = ~(U4387 & U7482 & U4482); 
assign U3384 = ~(U7482 & U4465 & U2605 & U4482 & U4387); 
assign U3385 = ~(U2605 & U4448 & U4159 & U4437 & U4388); 
assign U3396 = ~(U4448 & U3378); 
assign U3405 = ~(U4482 & STATE2_REG_0__SCAN_IN); 
assign U3406 = ~(U4387 & U7482); 
assign U3426 = ~(U4437 & STATE2_REG_2__SCAN_IN); 
assign U3436 = ~(U4465 & U4484); 
assign U3451 = ~(U7640 & U7639); 
assign U3452 = ~(U7642 & U7641); 
assign U3546 = U3378 & U3270 & U7482; 
assign U3547 = U4448 & U2605 & U4388; 
assign U3565 = U4387 & U4159; 
assign U3567 = U3271 & U3270 & U4388 & U7482; 
assign U3720 = U4482 & U4387; 
assign U3729 = U4437 & U4388; 
assign U3743 = U3271 & U3394; 
assign U3850 = U3270 & U3249 & U7482; 
assign U3873 = U3258 & U7482 & STATE2_REG_0__SCAN_IN; 
assign U3874 = U4387 & U4159; 
assign U3958 = U6609 & U6608 & U6607 & U6606; 
assign U3959 = U6613 & U6612 & U6611 & U6610; 
assign U3962 = U6625 & U6624 & U6623 & U6622; 
assign U3963 = U6629 & U6628 & U6627 & U6626; 
assign U3966 = U6641 & U6640 & U6639 & U6638; 
assign U3967 = U6645 & U6644 & U6643 & U6642; 
assign U3970 = U6657 & U6656 & U6655 & U6654; 
assign U3971 = U6661 & U6660 & U6659 & U6658; 
assign U3974 = U6672 & U6671 & U6670 & U6669; 
assign U3975 = U6676 & U6675 & U6674 & U6673; 
assign U3978 = U6688 & U6687 & U6686 & U6685; 
assign U3979 = U6692 & U6691 & U6690 & U6689; 
assign U3982 = U6704 & U6703 & U6702 & U6701; 
assign U3983 = U6708 & U6707 & U6706 & U6705; 
assign U3986 = U6720 & U6719 & U6718 & U6717; 
assign U3987 = U6724 & U6723 & U6722 & U6721; 
assign U3991 = U6740 & U6739; 
assign U3992 = U6743 & U6742; 
assign U3995 = U6750 & U6749; 
assign U4016 = U7482 & U6876 & U3270; 
assign U4053 = U7065 & U7064 & U7063 & U7062; 
assign U4069 = U7097 & U7096 & U7095 & U7094; 
assign U4073 = U7114 & U7113 & U7112 & U7111; 
assign U4077 = U7131 & U7130 & U7129 & U7128; 
assign U4079 = U7605 & U7134 & U4078; 
assign U4082 = U7146 & U7145 & U7144 & U7143; 
assign U4086 = U7163 & U7162 & U7161 & U7160; 
assign U4090 = U7180 & U7179 & U7178 & U7177; 
assign U4094 = U7197 & U7196 & U7195 & U7194; 
assign U4154 = U3440 & U7372; 
assign U4157 = U7453 & U7452; 
assign U4174 = ~U3399; 
assign U4178 = ~U3277; 
assign U4180 = ~U3392; 
assign U4183 = ~(U4253 & U3258); 
assign U4184 = ~(U4448 & U2605); 
assign U4198 = ~U3377; 
assign U4207 = ~(U4437 & U3258); 
assign U4219 = ~U3394; 
assign U4235 = ~U3381; 
assign U4245 = ~U3376; 
assign U4491 = ~(U4448 & U4161); 
assign U4533 = ~U3309; 
assign U4546 = ~(U3309 & STATE2_REG_2__SCAN_IN); 
assign U4604 = ~(U4593 & STATE2_REG_2__SCAN_IN); 
assign U4652 = ~U3323; 
assign U4663 = ~(U3323 & STATE2_REG_2__SCAN_IN); 
assign U4720 = ~(U4709 & STATE2_REG_2__SCAN_IN); 
assign U4824 = ~U3225; 
assign U4830 = ~(U3225 & STATE2_REG_2__SCAN_IN); 
assign U4939 = ~U3226; 
assign U4945 = ~(U3226 & STATE2_REG_2__SCAN_IN); 
assign U5052 = ~U3227; 
assign U5058 = ~(U3227 & STATE2_REG_2__SCAN_IN); 
assign U5167 = ~U3228; 
assign U5173 = ~(U3228 & STATE2_REG_2__SCAN_IN); 
assign U5282 = ~U3229; 
assign U5288 = ~(U3229 & STATE2_REG_2__SCAN_IN); 
assign U5397 = ~U3230; 
assign U5403 = ~(U3230 & STATE2_REG_2__SCAN_IN); 
assign U5451 = ~(U4388 & U4161 & U4448); 
assign U5475 = ~(U4482 & U3277); 
assign U5478 = ~(U4437 & U5476); 
assign U5482 = ~(U4448 & U4159); 
assign U5546 = ~(U4465 & U3259); 
assign U6614 = ~(U2534 & INSTQUEUE_REG_7__7__SCAN_IN); 
assign U6615 = ~(U2533 & INSTQUEUE_REG_6__7__SCAN_IN); 
assign U6616 = ~(U2532 & INSTQUEUE_REG_5__7__SCAN_IN); 
assign U6617 = ~(U2531 & INSTQUEUE_REG_4__7__SCAN_IN); 
assign U6618 = ~(U2529 & INSTQUEUE_REG_3__7__SCAN_IN); 
assign U6619 = ~(U2527 & INSTQUEUE_REG_2__7__SCAN_IN); 
assign U6620 = ~(U2525 & INSTQUEUE_REG_1__7__SCAN_IN); 
assign U6621 = ~(U2523 & INSTQUEUE_REG_0__7__SCAN_IN); 
assign U6630 = ~(U2534 & INSTQUEUE_REG_7__6__SCAN_IN); 
assign U6631 = ~(U2533 & INSTQUEUE_REG_6__6__SCAN_IN); 
assign U6632 = ~(U2532 & INSTQUEUE_REG_5__6__SCAN_IN); 
assign U6633 = ~(U2531 & INSTQUEUE_REG_4__6__SCAN_IN); 
assign U6634 = ~(U2529 & INSTQUEUE_REG_3__6__SCAN_IN); 
assign U6635 = ~(U2527 & INSTQUEUE_REG_2__6__SCAN_IN); 
assign U6636 = ~(U2525 & INSTQUEUE_REG_1__6__SCAN_IN); 
assign U6637 = ~(U2523 & INSTQUEUE_REG_0__6__SCAN_IN); 
assign U6646 = ~(U2534 & INSTQUEUE_REG_7__5__SCAN_IN); 
assign U6647 = ~(U2533 & INSTQUEUE_REG_6__5__SCAN_IN); 
assign U6648 = ~(U2532 & INSTQUEUE_REG_5__5__SCAN_IN); 
assign U6649 = ~(U2531 & INSTQUEUE_REG_4__5__SCAN_IN); 
assign U6650 = ~(U2529 & INSTQUEUE_REG_3__5__SCAN_IN); 
assign U6651 = ~(U2527 & INSTQUEUE_REG_2__5__SCAN_IN); 
assign U6652 = ~(U2525 & INSTQUEUE_REG_1__5__SCAN_IN); 
assign U6653 = ~(U2523 & INSTQUEUE_REG_0__5__SCAN_IN); 
assign U6662 = ~(U2534 & INSTQUEUE_REG_7__4__SCAN_IN); 
assign U6663 = ~(U2533 & INSTQUEUE_REG_6__4__SCAN_IN); 
assign U6664 = ~(U2532 & INSTQUEUE_REG_5__4__SCAN_IN); 
assign U6665 = ~(U2531 & INSTQUEUE_REG_4__4__SCAN_IN); 
assign U6666 = ~(U2529 & INSTQUEUE_REG_3__4__SCAN_IN); 
assign U6667 = ~(U2527 & INSTQUEUE_REG_2__4__SCAN_IN); 
assign U6668 = ~(U2525 & INSTQUEUE_REG_1__4__SCAN_IN); 
assign U6677 = ~(U2534 & INSTQUEUE_REG_7__3__SCAN_IN); 
assign U6678 = ~(U2533 & INSTQUEUE_REG_6__3__SCAN_IN); 
assign U6679 = ~(U2532 & INSTQUEUE_REG_5__3__SCAN_IN); 
assign U6680 = ~(U2531 & INSTQUEUE_REG_4__3__SCAN_IN); 
assign U6681 = ~(U2529 & INSTQUEUE_REG_3__3__SCAN_IN); 
assign U6682 = ~(U2527 & INSTQUEUE_REG_2__3__SCAN_IN); 
assign U6683 = ~(U2525 & INSTQUEUE_REG_1__3__SCAN_IN); 
assign U6684 = ~(U2523 & INSTQUEUE_REG_0__3__SCAN_IN); 
assign U6693 = ~(U2534 & INSTQUEUE_REG_7__2__SCAN_IN); 
assign U6694 = ~(U2533 & INSTQUEUE_REG_6__2__SCAN_IN); 
assign U6695 = ~(U2532 & INSTQUEUE_REG_5__2__SCAN_IN); 
assign U6696 = ~(U2531 & INSTQUEUE_REG_4__2__SCAN_IN); 
assign U6697 = ~(U2529 & INSTQUEUE_REG_3__2__SCAN_IN); 
assign U6698 = ~(U2527 & INSTQUEUE_REG_2__2__SCAN_IN); 
assign U6699 = ~(U2525 & INSTQUEUE_REG_1__2__SCAN_IN); 
assign U6700 = ~(U2523 & INSTQUEUE_REG_0__2__SCAN_IN); 
assign U6709 = ~(U2534 & INSTQUEUE_REG_7__1__SCAN_IN); 
assign U6710 = ~(U2533 & INSTQUEUE_REG_6__1__SCAN_IN); 
assign U6711 = ~(U2532 & INSTQUEUE_REG_5__1__SCAN_IN); 
assign U6712 = ~(U2531 & INSTQUEUE_REG_4__1__SCAN_IN); 
assign U6713 = ~(U2529 & INSTQUEUE_REG_3__1__SCAN_IN); 
assign U6714 = ~(U2527 & INSTQUEUE_REG_2__1__SCAN_IN); 
assign U6715 = ~(U2525 & INSTQUEUE_REG_1__1__SCAN_IN); 
assign U6716 = ~(U2523 & INSTQUEUE_REG_0__1__SCAN_IN); 
assign U6725 = ~(U2534 & INSTQUEUE_REG_7__0__SCAN_IN); 
assign U6726 = ~(U2533 & INSTQUEUE_REG_6__0__SCAN_IN); 
assign U6727 = ~(U2532 & INSTQUEUE_REG_5__0__SCAN_IN); 
assign U6728 = ~(U2531 & INSTQUEUE_REG_4__0__SCAN_IN); 
assign U6729 = ~(U2529 & INSTQUEUE_REG_3__0__SCAN_IN); 
assign U6730 = ~(U2527 & INSTQUEUE_REG_2__0__SCAN_IN); 
assign U6731 = ~(U2525 & INSTQUEUE_REG_1__0__SCAN_IN); 
assign U6732 = ~(U2523 & INSTQUEUE_REG_0__0__SCAN_IN); 
assign U6733 = ~(U4448 & STATE2_REG_2__SCAN_IN); 
assign U6873 = ~(U4482 & U3270); 
assign U6879 = ~(U4482 & U3270); 
assign U6880 = ~(U2564 & INSTQUEUE_REG_15__1__SCAN_IN); 
assign U6881 = ~(U2563 & INSTQUEUE_REG_14__1__SCAN_IN); 
assign U6882 = ~(U2562 & INSTQUEUE_REG_13__1__SCAN_IN); 
assign U6883 = ~(U2561 & INSTQUEUE_REG_12__1__SCAN_IN); 
assign U6884 = ~(U2559 & INSTQUEUE_REG_11__1__SCAN_IN); 
assign U6885 = ~(U2558 & INSTQUEUE_REG_10__1__SCAN_IN); 
assign U6886 = ~(U2557 & INSTQUEUE_REG_9__1__SCAN_IN); 
assign U6887 = ~(U2556 & INSTQUEUE_REG_8__1__SCAN_IN); 
assign U6898 = ~(U2564 & INSTQUEUE_REG_15__0__SCAN_IN); 
assign U6899 = ~(U2563 & INSTQUEUE_REG_14__0__SCAN_IN); 
assign U6900 = ~(U2562 & INSTQUEUE_REG_13__0__SCAN_IN); 
assign U6901 = ~(U2561 & INSTQUEUE_REG_12__0__SCAN_IN); 
assign U6902 = ~(U2559 & INSTQUEUE_REG_11__0__SCAN_IN); 
assign U6903 = ~(U2558 & INSTQUEUE_REG_10__0__SCAN_IN); 
assign U6904 = ~(U2557 & INSTQUEUE_REG_9__0__SCAN_IN); 
assign U6905 = ~(U2556 & INSTQUEUE_REG_8__0__SCAN_IN); 
assign U6929 = ~(U2564 & INSTQUEUE_REG_15__7__SCAN_IN); 
assign U6930 = ~(U2563 & INSTQUEUE_REG_14__7__SCAN_IN); 
assign U6931 = ~(U2562 & INSTQUEUE_REG_13__7__SCAN_IN); 
assign U6932 = ~(U2561 & INSTQUEUE_REG_12__7__SCAN_IN); 
assign U6933 = ~(U2559 & INSTQUEUE_REG_11__7__SCAN_IN); 
assign U6934 = ~(U2558 & INSTQUEUE_REG_10__7__SCAN_IN); 
assign U6935 = ~(U2557 & INSTQUEUE_REG_9__7__SCAN_IN); 
assign U6936 = ~(U2556 & INSTQUEUE_REG_8__7__SCAN_IN); 
assign U6946 = ~(U2564 & INSTQUEUE_REG_15__6__SCAN_IN); 
assign U6947 = ~(U2563 & INSTQUEUE_REG_14__6__SCAN_IN); 
assign U6948 = ~(U2562 & INSTQUEUE_REG_13__6__SCAN_IN); 
assign U6949 = ~(U2561 & INSTQUEUE_REG_12__6__SCAN_IN); 
assign U6950 = ~(U2559 & INSTQUEUE_REG_11__6__SCAN_IN); 
assign U6951 = ~(U2558 & INSTQUEUE_REG_10__6__SCAN_IN); 
assign U6952 = ~(U2557 & INSTQUEUE_REG_9__6__SCAN_IN); 
assign U6953 = ~(U2556 & INSTQUEUE_REG_8__6__SCAN_IN); 
assign U6963 = ~(U2564 & INSTQUEUE_REG_15__5__SCAN_IN); 
assign U6964 = ~(U2563 & INSTQUEUE_REG_14__5__SCAN_IN); 
assign U6965 = ~(U2562 & INSTQUEUE_REG_13__5__SCAN_IN); 
assign U6966 = ~(U2561 & INSTQUEUE_REG_12__5__SCAN_IN); 
assign U6967 = ~(U2559 & INSTQUEUE_REG_11__5__SCAN_IN); 
assign U6968 = ~(U2558 & INSTQUEUE_REG_10__5__SCAN_IN); 
assign U6969 = ~(U2557 & INSTQUEUE_REG_9__5__SCAN_IN); 
assign U6970 = ~(U2556 & INSTQUEUE_REG_8__5__SCAN_IN); 
assign U6980 = ~(U2564 & INSTQUEUE_REG_15__4__SCAN_IN); 
assign U6981 = ~(U2563 & INSTQUEUE_REG_14__4__SCAN_IN); 
assign U6982 = ~(U2562 & INSTQUEUE_REG_13__4__SCAN_IN); 
assign U6983 = ~(U2561 & INSTQUEUE_REG_12__4__SCAN_IN); 
assign U6984 = ~(U2559 & INSTQUEUE_REG_11__4__SCAN_IN); 
assign U6985 = ~(U2558 & INSTQUEUE_REG_10__4__SCAN_IN); 
assign U6986 = ~(U2557 & INSTQUEUE_REG_9__4__SCAN_IN); 
assign U6987 = ~(U2556 & INSTQUEUE_REG_8__4__SCAN_IN); 
assign U6995 = ~(U2564 & INSTQUEUE_REG_15__3__SCAN_IN); 
assign U6996 = ~(U2563 & INSTQUEUE_REG_14__3__SCAN_IN); 
assign U6997 = ~(U2562 & INSTQUEUE_REG_13__3__SCAN_IN); 
assign U6998 = ~(U2561 & INSTQUEUE_REG_12__3__SCAN_IN); 
assign U6999 = ~(U2559 & INSTQUEUE_REG_11__3__SCAN_IN); 
assign U7000 = ~(U2558 & INSTQUEUE_REG_10__3__SCAN_IN); 
assign U7001 = ~(U2557 & INSTQUEUE_REG_9__3__SCAN_IN); 
assign U7002 = ~(U2556 & INSTQUEUE_REG_8__3__SCAN_IN); 
assign U7012 = ~(U2564 & INSTQUEUE_REG_15__2__SCAN_IN); 
assign U7013 = ~(U2563 & INSTQUEUE_REG_14__2__SCAN_IN); 
assign U7014 = ~(U2562 & INSTQUEUE_REG_13__2__SCAN_IN); 
assign U7015 = ~(U2561 & INSTQUEUE_REG_12__2__SCAN_IN); 
assign U7016 = ~(U2559 & INSTQUEUE_REG_11__2__SCAN_IN); 
assign U7017 = ~(U2558 & INSTQUEUE_REG_10__2__SCAN_IN); 
assign U7018 = ~(U2557 & INSTQUEUE_REG_9__2__SCAN_IN); 
assign U7019 = ~(U2556 & INSTQUEUE_REG_8__2__SCAN_IN); 
assign U7208 = ~(U2602 & INSTQUEUE_REG_8__7__SCAN_IN); 
assign U7209 = ~(U2601 & INSTQUEUE_REG_9__7__SCAN_IN); 
assign U7210 = ~(U2600 & INSTQUEUE_REG_10__7__SCAN_IN); 
assign U7211 = ~(U2599 & INSTQUEUE_REG_11__7__SCAN_IN); 
assign U7212 = ~(U2597 & INSTQUEUE_REG_12__7__SCAN_IN); 
assign U7213 = ~(U2596 & INSTQUEUE_REG_13__7__SCAN_IN); 
assign U7214 = ~(U2595 & INSTQUEUE_REG_14__7__SCAN_IN); 
assign U7215 = ~(U2594 & INSTQUEUE_REG_15__7__SCAN_IN); 
assign U7225 = ~(U2602 & INSTQUEUE_REG_8__6__SCAN_IN); 
assign U7226 = ~(U2601 & INSTQUEUE_REG_9__6__SCAN_IN); 
assign U7227 = ~(U2600 & INSTQUEUE_REG_10__6__SCAN_IN); 
assign U7228 = ~(U2599 & INSTQUEUE_REG_11__6__SCAN_IN); 
assign U7229 = ~(U2597 & INSTQUEUE_REG_12__6__SCAN_IN); 
assign U7230 = ~(U2596 & INSTQUEUE_REG_13__6__SCAN_IN); 
assign U7231 = ~(U2595 & INSTQUEUE_REG_14__6__SCAN_IN); 
assign U7232 = ~(U2594 & INSTQUEUE_REG_15__6__SCAN_IN); 
assign U7242 = ~(U2602 & INSTQUEUE_REG_8__5__SCAN_IN); 
assign U7243 = ~(U2601 & INSTQUEUE_REG_9__5__SCAN_IN); 
assign U7244 = ~(U2600 & INSTQUEUE_REG_10__5__SCAN_IN); 
assign U7245 = ~(U2599 & INSTQUEUE_REG_11__5__SCAN_IN); 
assign U7246 = ~(U2597 & INSTQUEUE_REG_12__5__SCAN_IN); 
assign U7247 = ~(U2596 & INSTQUEUE_REG_13__5__SCAN_IN); 
assign U7248 = ~(U2595 & INSTQUEUE_REG_14__5__SCAN_IN); 
assign U7249 = ~(U2594 & INSTQUEUE_REG_15__5__SCAN_IN); 
assign U7259 = ~(U2602 & INSTQUEUE_REG_8__4__SCAN_IN); 
assign U7260 = ~(U2601 & INSTQUEUE_REG_9__4__SCAN_IN); 
assign U7261 = ~(U2600 & INSTQUEUE_REG_10__4__SCAN_IN); 
assign U7262 = ~(U2599 & INSTQUEUE_REG_11__4__SCAN_IN); 
assign U7263 = ~(U2597 & INSTQUEUE_REG_12__4__SCAN_IN); 
assign U7264 = ~(U2596 & INSTQUEUE_REG_13__4__SCAN_IN); 
assign U7265 = ~(U2595 & INSTQUEUE_REG_14__4__SCAN_IN); 
assign U7266 = ~(U2594 & INSTQUEUE_REG_15__4__SCAN_IN); 
assign U7274 = ~(U2602 & INSTQUEUE_REG_8__3__SCAN_IN); 
assign U7275 = ~(U2601 & INSTQUEUE_REG_9__3__SCAN_IN); 
assign U7276 = ~(U2600 & INSTQUEUE_REG_10__3__SCAN_IN); 
assign U7277 = ~(U2599 & INSTQUEUE_REG_11__3__SCAN_IN); 
assign U7278 = ~(U2597 & INSTQUEUE_REG_12__3__SCAN_IN); 
assign U7279 = ~(U2596 & INSTQUEUE_REG_13__3__SCAN_IN); 
assign U7280 = ~(U2595 & INSTQUEUE_REG_14__3__SCAN_IN); 
assign U7281 = ~(U2594 & INSTQUEUE_REG_15__3__SCAN_IN); 
assign U7291 = ~(U2602 & INSTQUEUE_REG_8__2__SCAN_IN); 
assign U7292 = ~(U2601 & INSTQUEUE_REG_9__2__SCAN_IN); 
assign U7293 = ~(U2600 & INSTQUEUE_REG_10__2__SCAN_IN); 
assign U7294 = ~(U2599 & INSTQUEUE_REG_11__2__SCAN_IN); 
assign U7295 = ~(U2597 & INSTQUEUE_REG_12__2__SCAN_IN); 
assign U7296 = ~(U2596 & INSTQUEUE_REG_13__2__SCAN_IN); 
assign U7297 = ~(U2595 & INSTQUEUE_REG_14__2__SCAN_IN); 
assign U7298 = ~(U2594 & INSTQUEUE_REG_15__2__SCAN_IN); 
assign U7308 = ~(U2602 & INSTQUEUE_REG_8__1__SCAN_IN); 
assign U7309 = ~(U2601 & INSTQUEUE_REG_9__1__SCAN_IN); 
assign U7310 = ~(U2600 & INSTQUEUE_REG_10__1__SCAN_IN); 
assign U7311 = ~(U2599 & INSTQUEUE_REG_11__1__SCAN_IN); 
assign U7312 = ~(U2597 & INSTQUEUE_REG_12__1__SCAN_IN); 
assign U7313 = ~(U2596 & INSTQUEUE_REG_13__1__SCAN_IN); 
assign U7314 = ~(U2595 & INSTQUEUE_REG_14__1__SCAN_IN); 
assign U7315 = ~(U2594 & INSTQUEUE_REG_15__1__SCAN_IN); 
assign U7325 = ~(U2602 & INSTQUEUE_REG_8__0__SCAN_IN); 
assign U7326 = ~(U2601 & INSTQUEUE_REG_9__0__SCAN_IN); 
assign U7327 = ~(U2600 & INSTQUEUE_REG_10__0__SCAN_IN); 
assign U7328 = ~(U2599 & INSTQUEUE_REG_11__0__SCAN_IN); 
assign U7329 = ~(U2597 & INSTQUEUE_REG_12__0__SCAN_IN); 
assign U7330 = ~(U2596 & INSTQUEUE_REG_13__0__SCAN_IN); 
assign U7331 = ~(U2595 & INSTQUEUE_REG_14__0__SCAN_IN); 
assign U7332 = ~(U2594 & INSTQUEUE_REG_15__0__SCAN_IN); 
assign U7444 = ~(U4465 & U4484); 
assign U7601 = ~(U2523 & INSTQUEUE_REG_0__4__SCAN_IN); 
assign U7691 = ~(U4448 & U3265); 
assign U7773 = ~(U4448 & U7483); 
assign R2027_U53 = ~(R2027_U146 & R2027_U145); 
assign R2027_U54 = ~(R2027_U148 & R2027_U147); 
assign R2027_U120 = ~R2027_U17; 
assign R2027_U125 = ~R2027_U95; 
assign R2027_U142 = ~(R2027_U17 & INSTADDRPOINTER_REG_9__SCAN_IN); 
assign R2027_U143 = ~(R2027_U95 & INSTADDRPOINTER_REG_8__SCAN_IN); 
assign R2337_U51 = ~(R2337_U135 & R2337_U134); 
assign R2337_U80 = ~(R2337_U193 & R2337_U192); 
assign R2337_U113 = ~R2337_U104; 
assign R2337_U114 = ~R2337_U20; 
assign R2337_U188 = ~(R2337_U20 & PHYADDRPOINTER_REG_12__SCAN_IN); 
assign R2337_U190 = ~(R2337_U104 & PHYADDRPOINTER_REG_11__SCAN_IN); 
assign R2096_U66 = ~(R2096_U132 & R2096_U131); 
assign R2096_U97 = ~R2096_U12; 
assign R2096_U129 = ~(R2096_U12 & REIP_REG_6__SCAN_IN); 
assign R2238_U27 = ~(R2238_U37 & R2238_U36); 
assign R2238_U60 = ~(R2238_U34 & R2238_U59); 
assign SUB_450_U27 = ~(SUB_450_U37 & SUB_450_U36); 
assign SUB_450_U60 = ~(SUB_450_U34 & SUB_450_U59); 
assign ADD_405_U67 = ~(ADD_405_U136 & ADD_405_U135); 
assign ADD_405_U100 = ~ADD_405_U12; 
assign ADD_405_U133 = ~(ADD_405_U12 & INSTADDRPOINTER_REG_6__SCAN_IN); 
assign ADD_515_U66 = ~(ADD_515_U132 & ADD_515_U131); 
assign ADD_515_U97 = ~ADD_515_U12; 
assign ADD_515_U129 = ~(ADD_515_U12 & INSTADDRPOINTER_REG_6__SCAN_IN); 
assign U2353 = U4219 & STATE2_REG_2__SCAN_IN; 
assign U2447 = U3565 & U2452; 
assign U2678 = ~(U7444 & U3271); 
assign U2722 = ~(U4147 & U4180); 
assign U3231 = ~(U3378 & U3381 & U5451); 
assign U3266 = ~(U3547 & U3546); 
assign U3273 = ~(U2389 & U3270); 
assign U3278 = ~(U4178 & U3271); 
assign U3383 = ~(U3729 & U4235); 
assign U3398 = ~(U4178 & U2452); 
assign U3409 = ~(U4198 & STATE2_REG_0__SCAN_IN); 
assign U3410 = ~(U4491 & U3378); 
assign U3722 = U4198 & U3244; 
assign U3742 = U5546 & U3244; 
assign U3747 = U4174 & U3271; 
assign U3854 = U2449 & STATE2_REG_0__SCAN_IN; 
assign U3877 = U4482 & U4174; 
assign U3956 = U3274 & STATE2_REG_2__SCAN_IN; 
assign U3960 = U6617 & U6616 & U6615 & U6614; 
assign U3961 = U6621 & U6620 & U6619 & U6618; 
assign U3964 = U6633 & U6632 & U6631 & U6630; 
assign U3965 = U6637 & U6636 & U6635 & U6634; 
assign U3968 = U6649 & U6648 & U6647 & U6646; 
assign U3969 = U6653 & U6652 & U6651 & U6650; 
assign U3972 = U6665 & U6664 & U6663 & U6662; 
assign U3973 = U7601 & U6668 & U6667 & U6666; 
assign U3976 = U6680 & U6679 & U6678 & U6677; 
assign U3977 = U6684 & U6683 & U6682 & U6681; 
assign U3980 = U6696 & U6695 & U6694 & U6693; 
assign U3981 = U6700 & U6699 & U6698 & U6697; 
assign U3984 = U6712 & U6711 & U6710 & U6709; 
assign U3985 = U6716 & U6715 & U6714 & U6713; 
assign U3988 = U6728 & U6727 & U6726 & U6725; 
assign U3989 = U6732 & U6731 & U6730 & U6729; 
assign U4017 = U6883 & U6882 & U6881 & U6880; 
assign U4018 = U6887 & U6886 & U6885 & U6884; 
assign U4021 = U6901 & U6900 & U6899 & U6898; 
assign U4022 = U6905 & U6904 & U6903 & U6902; 
assign U4025 = U6932 & U6931 & U6930 & U6929; 
assign U4026 = U6936 & U6935 & U6934 & U6933; 
assign U4029 = U6949 & U6948 & U6947 & U6946; 
assign U4030 = U6953 & U6952 & U6951 & U6950; 
assign U4033 = U6966 & U6965 & U6964 & U6963; 
assign U4034 = U6970 & U6969 & U6968 & U6967; 
assign U4037 = U6983 & U6982 & U6981 & U6980; 
assign U4038 = U6987 & U6986 & U6985 & U6984; 
assign U4041 = U6998 & U6997 & U6996 & U6995; 
assign U4042 = U7002 & U7001 & U7000 & U6999; 
assign U4045 = U7015 & U7014 & U7013 & U7012; 
assign U4046 = U7019 & U7018 & U7017 & U7016; 
assign U4109 = U7211 & U7210 & U7209 & U7208; 
assign U4110 = U7215 & U7214 & U7213 & U7212; 
assign U4113 = U7228 & U7227 & U7226 & U7225; 
assign U4114 = U7232 & U7231 & U7230 & U7229; 
assign U4117 = U7245 & U7244 & U7243 & U7242; 
assign U4118 = U7249 & U7248 & U7247 & U7246; 
assign U4121 = U7262 & U7261 & U7260 & U7259; 
assign U4122 = U7266 & U7265 & U7264 & U7263; 
assign U4125 = U7277 & U7276 & U7275 & U7274; 
assign U4126 = U7281 & U7280 & U7279 & U7278; 
assign U4129 = U7294 & U7293 & U7292 & U7291; 
assign U4130 = U7298 & U7297 & U7296 & U7295; 
assign U4133 = U7311 & U7310 & U7309 & U7308; 
assign U4134 = U7315 & U7314 & U7313 & U7312; 
assign U4137 = U7328 & U7327 & U7326 & U7325; 
assign U4138 = U7332 & U7331 & U7330 & U7329; 
assign U4141 = U3271 & U3406; 
assign U4176 = ~U3426; 
assign U4177 = ~U3380; 
assign U4179 = ~U3436; 
assign U4187 = ~U3276; 
assign U4194 = ~U3405; 
assign U4196 = ~U3269; 
assign U4222 = ~U3382; 
assign U4224 = ~U3385; 
assign U4237 = ~U3274; 
assign U4238 = ~U3384; 
assign U4241 = ~U3396; 
assign U4242 = ~U3406; 
assign U4488 = ~(U3259 & U3377 & U3274); 
assign U4541 = ~(U4533 & STATE2_REG_2__SCAN_IN); 
assign U4658 = ~(U4652 & STATE2_REG_2__SCAN_IN); 
assign U4767 = ~U3332; 
assign U4778 = ~(U3332 & STATE2_REG_2__SCAN_IN); 
assign U4835 = ~(U4824 & STATE2_REG_2__SCAN_IN); 
assign U4882 = ~U3339; 
assign U4893 = ~(U3339 & STATE2_REG_2__SCAN_IN); 
assign U4950 = ~(U4939 & STATE2_REG_2__SCAN_IN); 
assign U4996 = ~U3349; 
assign U5006 = ~(U3349 & STATE2_REG_2__SCAN_IN); 
assign U5063 = ~(U5052 & STATE2_REG_2__SCAN_IN); 
assign U5110 = ~U3356; 
assign U5121 = ~(U3356 & STATE2_REG_2__SCAN_IN); 
assign U5178 = ~(U5167 & STATE2_REG_2__SCAN_IN); 
assign U5225 = ~U3363; 
assign U5236 = ~(U3363 & STATE2_REG_2__SCAN_IN); 
assign U5293 = ~(U5282 & STATE2_REG_2__SCAN_IN); 
assign U5340 = ~U3370; 
assign U5351 = ~(U3370 & STATE2_REG_2__SCAN_IN); 
assign U5408 = ~(U5397 & STATE2_REG_2__SCAN_IN); 
assign U5450 = ~(U3378 & U3381 & U4491); 
assign U5453 = ~(U4482 & U3276); 
assign U5455 = ~(U3720 & U2452); 
assign U5459 = ~(U2449 & U7482); 
assign U5460 = ~(U4245 & U4491); 
assign U5477 = ~(U7692 & U7691 & U7482); 
assign U5479 = ~(U4388 & U3381 & U3396); 
assign U5483 = ~(U3382 & U5482); 
assign U5485 = ~(U4245 & U4491); 
assign U5549 = ~(U4223 & U4491 & U4180); 
assign U5947 = ~(READY_N & U3269); 
assign U6734 = ~(U3399 & U6733); 
assign U6737 = ~(R2337_U51 & U2352); 
assign U6846 = ~(R2337_U80 & U2352); 
assign U6888 = ~(U2554 & INSTQUEUE_REG_7__1__SCAN_IN); 
assign U6889 = ~(U2553 & INSTQUEUE_REG_6__1__SCAN_IN); 
assign U6890 = ~(U2552 & INSTQUEUE_REG_5__1__SCAN_IN); 
assign U6891 = ~(U2551 & INSTQUEUE_REG_4__1__SCAN_IN); 
assign U6892 = ~(U2549 & INSTQUEUE_REG_3__1__SCAN_IN); 
assign U6893 = ~(U2548 & INSTQUEUE_REG_2__1__SCAN_IN); 
assign U6894 = ~(U2547 & INSTQUEUE_REG_1__1__SCAN_IN); 
assign U6895 = ~(U2546 & INSTQUEUE_REG_0__1__SCAN_IN); 
assign U6897 = ~(U3392 & U3405); 
assign U6906 = ~(U2554 & INSTQUEUE_REG_7__0__SCAN_IN); 
assign U6907 = ~(U2553 & INSTQUEUE_REG_6__0__SCAN_IN); 
assign U6908 = ~(U2552 & INSTQUEUE_REG_5__0__SCAN_IN); 
assign U6909 = ~(U2551 & INSTQUEUE_REG_4__0__SCAN_IN); 
assign U6910 = ~(U2549 & INSTQUEUE_REG_3__0__SCAN_IN); 
assign U6911 = ~(U2548 & INSTQUEUE_REG_2__0__SCAN_IN); 
assign U6912 = ~(U2547 & INSTQUEUE_REG_1__0__SCAN_IN); 
assign U6913 = ~(U2546 & INSTQUEUE_REG_0__0__SCAN_IN); 
assign U6937 = ~(U2554 & INSTQUEUE_REG_7__7__SCAN_IN); 
assign U6938 = ~(U2553 & INSTQUEUE_REG_6__7__SCAN_IN); 
assign U6939 = ~(U2552 & INSTQUEUE_REG_5__7__SCAN_IN); 
assign U6940 = ~(U2551 & INSTQUEUE_REG_4__7__SCAN_IN); 
assign U6941 = ~(U2549 & INSTQUEUE_REG_3__7__SCAN_IN); 
assign U6942 = ~(U2548 & INSTQUEUE_REG_2__7__SCAN_IN); 
assign U6943 = ~(U2547 & INSTQUEUE_REG_1__7__SCAN_IN); 
assign U6944 = ~(U2546 & INSTQUEUE_REG_0__7__SCAN_IN); 
assign U6954 = ~(U2554 & INSTQUEUE_REG_7__6__SCAN_IN); 
assign U6955 = ~(U2553 & INSTQUEUE_REG_6__6__SCAN_IN); 
assign U6956 = ~(U2552 & INSTQUEUE_REG_5__6__SCAN_IN); 
assign U6957 = ~(U2551 & INSTQUEUE_REG_4__6__SCAN_IN); 
assign U6958 = ~(U2549 & INSTQUEUE_REG_3__6__SCAN_IN); 
assign U6959 = ~(U2548 & INSTQUEUE_REG_2__6__SCAN_IN); 
assign U6960 = ~(U2547 & INSTQUEUE_REG_1__6__SCAN_IN); 
assign U6961 = ~(U2546 & INSTQUEUE_REG_0__6__SCAN_IN); 
assign U6971 = ~(U2554 & INSTQUEUE_REG_7__5__SCAN_IN); 
assign U6972 = ~(U2553 & INSTQUEUE_REG_6__5__SCAN_IN); 
assign U6973 = ~(U2552 & INSTQUEUE_REG_5__5__SCAN_IN); 
assign U6974 = ~(U2551 & INSTQUEUE_REG_4__5__SCAN_IN); 
assign U6975 = ~(U2549 & INSTQUEUE_REG_3__5__SCAN_IN); 
assign U6976 = ~(U2548 & INSTQUEUE_REG_2__5__SCAN_IN); 
assign U6977 = ~(U2547 & INSTQUEUE_REG_1__5__SCAN_IN); 
assign U6978 = ~(U2546 & INSTQUEUE_REG_0__5__SCAN_IN); 
assign U6988 = ~(U2554 & INSTQUEUE_REG_7__4__SCAN_IN); 
assign U6989 = ~(U2553 & INSTQUEUE_REG_6__4__SCAN_IN); 
assign U6990 = ~(U2552 & INSTQUEUE_REG_5__4__SCAN_IN); 
assign U6991 = ~(U2551 & INSTQUEUE_REG_4__4__SCAN_IN); 
assign U6992 = ~(U2549 & INSTQUEUE_REG_3__4__SCAN_IN); 
assign U6993 = ~(U2548 & INSTQUEUE_REG_2__4__SCAN_IN); 
assign U6994 = ~(U2547 & INSTQUEUE_REG_1__4__SCAN_IN); 
assign U7003 = ~(U2554 & INSTQUEUE_REG_7__3__SCAN_IN); 
assign U7004 = ~(U2553 & INSTQUEUE_REG_6__3__SCAN_IN); 
assign U7005 = ~(U2552 & INSTQUEUE_REG_5__3__SCAN_IN); 
assign U7006 = ~(U2551 & INSTQUEUE_REG_4__3__SCAN_IN); 
assign U7007 = ~(U2549 & INSTQUEUE_REG_3__3__SCAN_IN); 
assign U7008 = ~(U2548 & INSTQUEUE_REG_2__3__SCAN_IN); 
assign U7009 = ~(U2547 & INSTQUEUE_REG_1__3__SCAN_IN); 
assign U7010 = ~(U2546 & INSTQUEUE_REG_0__3__SCAN_IN); 
assign U7020 = ~(U2554 & INSTQUEUE_REG_7__2__SCAN_IN); 
assign U7021 = ~(U2553 & INSTQUEUE_REG_6__2__SCAN_IN); 
assign U7022 = ~(U2552 & INSTQUEUE_REG_5__2__SCAN_IN); 
assign U7023 = ~(U2551 & INSTQUEUE_REG_4__2__SCAN_IN); 
assign U7024 = ~(U2549 & INSTQUEUE_REG_3__2__SCAN_IN); 
assign U7025 = ~(U2548 & INSTQUEUE_REG_2__2__SCAN_IN); 
assign U7026 = ~(U2547 & INSTQUEUE_REG_1__2__SCAN_IN); 
assign U7027 = ~(U2546 & INSTQUEUE_REG_0__2__SCAN_IN); 
assign U7036 = ~(U4180 & INSTQUEUE_REG_0__7__SCAN_IN); 
assign U7038 = ~(U4180 & INSTQUEUE_REG_0__6__SCAN_IN); 
assign U7040 = ~(U4180 & INSTQUEUE_REG_0__5__SCAN_IN); 
assign U7043 = ~(U4180 & INSTQUEUE_REG_0__3__SCAN_IN); 
assign U7045 = ~(U4180 & INSTQUEUE_REG_0__2__SCAN_IN); 
assign U7047 = ~(U4180 & INSTQUEUE_REG_0__1__SCAN_IN); 
assign U7050 = ~(U4180 & INSTQUEUE_REG_0__0__SCAN_IN); 
assign U7070 = ~(U4054 & U4053 & U4052 & U4051); 
assign U7074 = ~(U4491 & U3265); 
assign U7076 = ~(U4388 & U4491 & U4142 & U3381); 
assign U7102 = ~(U4070 & U4069 & U4068 & U4067); 
assign U7119 = ~(U4074 & U4073 & U4072 & U4071); 
assign U7151 = ~(U4083 & U4082 & U4081 & U4080); 
assign U7168 = ~(U4087 & U4086 & U4085 & U4084); 
assign U7185 = ~(U4091 & U4090 & U4089 & U4088); 
assign U7202 = ~(U4095 & U4094 & U4093 & U4092); 
assign U7216 = ~(U2592 & INSTQUEUE_REG_0__7__SCAN_IN); 
assign U7217 = ~(U2591 & INSTQUEUE_REG_1__7__SCAN_IN); 
assign U7218 = ~(U2590 & INSTQUEUE_REG_2__7__SCAN_IN); 
assign U7219 = ~(U2589 & INSTQUEUE_REG_3__7__SCAN_IN); 
assign U7220 = ~(U2587 & INSTQUEUE_REG_4__7__SCAN_IN); 
assign U7221 = ~(U2586 & INSTQUEUE_REG_5__7__SCAN_IN); 
assign U7222 = ~(U2585 & INSTQUEUE_REG_6__7__SCAN_IN); 
assign U7223 = ~(U2584 & INSTQUEUE_REG_7__7__SCAN_IN); 
assign U7233 = ~(U2592 & INSTQUEUE_REG_0__6__SCAN_IN); 
assign U7234 = ~(U2591 & INSTQUEUE_REG_1__6__SCAN_IN); 
assign U7235 = ~(U2590 & INSTQUEUE_REG_2__6__SCAN_IN); 
assign U7236 = ~(U2589 & INSTQUEUE_REG_3__6__SCAN_IN); 
assign U7237 = ~(U2587 & INSTQUEUE_REG_4__6__SCAN_IN); 
assign U7238 = ~(U2586 & INSTQUEUE_REG_5__6__SCAN_IN); 
assign U7239 = ~(U2585 & INSTQUEUE_REG_6__6__SCAN_IN); 
assign U7240 = ~(U2584 & INSTQUEUE_REG_7__6__SCAN_IN); 
assign U7250 = ~(U2592 & INSTQUEUE_REG_0__5__SCAN_IN); 
assign U7251 = ~(U2591 & INSTQUEUE_REG_1__5__SCAN_IN); 
assign U7252 = ~(U2590 & INSTQUEUE_REG_2__5__SCAN_IN); 
assign U7253 = ~(U2589 & INSTQUEUE_REG_3__5__SCAN_IN); 
assign U7254 = ~(U2587 & INSTQUEUE_REG_4__5__SCAN_IN); 
assign U7255 = ~(U2586 & INSTQUEUE_REG_5__5__SCAN_IN); 
assign U7256 = ~(U2585 & INSTQUEUE_REG_6__5__SCAN_IN); 
assign U7257 = ~(U2584 & INSTQUEUE_REG_7__5__SCAN_IN); 
assign U7267 = ~(U2591 & INSTQUEUE_REG_1__4__SCAN_IN); 
assign U7268 = ~(U2590 & INSTQUEUE_REG_2__4__SCAN_IN); 
assign U7269 = ~(U2589 & INSTQUEUE_REG_3__4__SCAN_IN); 
assign U7270 = ~(U2587 & INSTQUEUE_REG_4__4__SCAN_IN); 
assign U7271 = ~(U2586 & INSTQUEUE_REG_5__4__SCAN_IN); 
assign U7272 = ~(U2585 & INSTQUEUE_REG_6__4__SCAN_IN); 
assign U7273 = ~(U2584 & INSTQUEUE_REG_7__4__SCAN_IN); 
assign U7282 = ~(U2592 & INSTQUEUE_REG_0__3__SCAN_IN); 
assign U7283 = ~(U2591 & INSTQUEUE_REG_1__3__SCAN_IN); 
assign U7284 = ~(U2590 & INSTQUEUE_REG_2__3__SCAN_IN); 
assign U7285 = ~(U2589 & INSTQUEUE_REG_3__3__SCAN_IN); 
assign U7286 = ~(U2587 & INSTQUEUE_REG_4__3__SCAN_IN); 
assign U7287 = ~(U2586 & INSTQUEUE_REG_5__3__SCAN_IN); 
assign U7288 = ~(U2585 & INSTQUEUE_REG_6__3__SCAN_IN); 
assign U7289 = ~(U2584 & INSTQUEUE_REG_7__3__SCAN_IN); 
assign U7299 = ~(U2592 & INSTQUEUE_REG_0__2__SCAN_IN); 
assign U7300 = ~(U2591 & INSTQUEUE_REG_1__2__SCAN_IN); 
assign U7301 = ~(U2590 & INSTQUEUE_REG_2__2__SCAN_IN); 
assign U7302 = ~(U2589 & INSTQUEUE_REG_3__2__SCAN_IN); 
assign U7303 = ~(U2587 & INSTQUEUE_REG_4__2__SCAN_IN); 
assign U7304 = ~(U2586 & INSTQUEUE_REG_5__2__SCAN_IN); 
assign U7305 = ~(U2585 & INSTQUEUE_REG_6__2__SCAN_IN); 
assign U7306 = ~(U2584 & INSTQUEUE_REG_7__2__SCAN_IN); 
assign U7316 = ~(U2592 & INSTQUEUE_REG_0__1__SCAN_IN); 
assign U7317 = ~(U2591 & INSTQUEUE_REG_1__1__SCAN_IN); 
assign U7318 = ~(U2590 & INSTQUEUE_REG_2__1__SCAN_IN); 
assign U7319 = ~(U2589 & INSTQUEUE_REG_3__1__SCAN_IN); 
assign U7320 = ~(U2587 & INSTQUEUE_REG_4__1__SCAN_IN); 
assign U7321 = ~(U2586 & INSTQUEUE_REG_5__1__SCAN_IN); 
assign U7322 = ~(U2585 & INSTQUEUE_REG_6__1__SCAN_IN); 
assign U7323 = ~(U2584 & INSTQUEUE_REG_7__1__SCAN_IN); 
assign U7333 = ~(U2592 & INSTQUEUE_REG_0__0__SCAN_IN); 
assign U7334 = ~(U2591 & INSTQUEUE_REG_1__0__SCAN_IN); 
assign U7335 = ~(U2590 & INSTQUEUE_REG_2__0__SCAN_IN); 
assign U7336 = ~(U2589 & INSTQUEUE_REG_3__0__SCAN_IN); 
assign U7337 = ~(U2587 & INSTQUEUE_REG_4__0__SCAN_IN); 
assign U7338 = ~(U2586 & INSTQUEUE_REG_5__0__SCAN_IN); 
assign U7339 = ~(U2585 & INSTQUEUE_REG_6__0__SCAN_IN); 
assign U7340 = ~(U2584 & INSTQUEUE_REG_7__0__SCAN_IN); 
assign U7346 = ~(U4178 & U2452); 
assign U7350 = ~(U2451 & U4198); 
assign U7361 = ~(SUB_450_U22 & U2354); 
assign U7363 = ~(SUB_450_U7 & U2354); 
assign U7373 = ~(R2238_U22 & U4180); 
assign U7375 = ~(U2451 & U3271); 
assign U7376 = ~(R2238_U7 & U4180); 
assign U7378 = ~(U3380 & U3277); 
assign U7379 = ~(U3271 & U3436); 
assign U7478 = ~(U7773 & U7772 & U4060); 
assign U7602 = ~(U2546 & INSTQUEUE_REG_0__4__SCAN_IN); 
assign U7604 = ~(U4180 & INSTQUEUE_REG_0__4__SCAN_IN); 
assign U7606 = ~(U4079 & U4077 & U4076 & U4075); 
assign U7607 = ~(U2592 & INSTQUEUE_REG_0__4__SCAN_IN); 
assign U7615 = ~(U5475 & U4159); 
assign U7616 = ~(U3270 & U3276); 
assign U7619 = ~(U5475 & U4159); 
assign R2027_U22 = ~(R2027_U85 & R2027_U120); 
assign R2027_U110 = ~(R2027_U120 & INSTADDRPOINTER_REG_9__SCAN_IN); 
assign R2027_U141 = ~(R2027_U120 & R2027_U18); 
assign R2027_U144 = ~(R2027_U125 & R2027_U14); 
assign R2337_U23 = ~(R2337_U84 & R2337_U114); 
assign R2337_U103 = ~(R2337_U114 & PHYADDRPOINTER_REG_12__SCAN_IN); 
assign R2337_U189 = ~(R2337_U114 & R2337_U22); 
assign R2337_U191 = ~(R2337_U113 & R2337_U18); 
assign R2099_U4 = ~U4178; 
assign R2096_U14 = ~(R2096_U97 & REIP_REG_6__SCAN_IN); 
assign R2096_U130 = ~(R2096_U97 & R2096_U13); 
assign R2238_U21 = ~(R2238_U61 & R2238_U60); 
assign R2238_U38 = ~R2238_U27; 
assign R2238_U40 = ~(R2238_U39 & R2238_U27); 
assign R2238_U56 = ~(R2238_U24 & R2238_U27); 
assign SUB_450_U21 = ~(SUB_450_U61 & SUB_450_U60); 
assign SUB_450_U38 = ~SUB_450_U27; 
assign SUB_450_U40 = ~(SUB_450_U39 & SUB_450_U27); 
assign SUB_450_U56 = ~(SUB_450_U24 & SUB_450_U27); 
assign ADD_405_U14 = ~(ADD_405_U100 & INSTADDRPOINTER_REG_6__SCAN_IN); 
assign ADD_405_U134 = ~(ADD_405_U100 & ADD_405_U13); 
assign ADD_515_U14 = ~(ADD_515_U97 & INSTADDRPOINTER_REG_6__SCAN_IN); 
assign ADD_515_U130 = ~(ADD_515_U97 & ADD_515_U13); 
assign U2431 = U4187 & U7482; 
assign U3214 = ~(U3989 & U3988 & U3987 & U3986); 
assign U3215 = ~(U3985 & U3984 & U3983 & U3982); 
assign U3216 = ~(U3981 & U3980 & U3979 & U3978); 
assign U3217 = ~(U3977 & U3976 & U3975 & U3974); 
assign U3218 = ~(U3973 & U3972 & U3971 & U3970); 
assign U3219 = ~(U3969 & U3968 & U3967 & U3966); 
assign U3220 = ~(U3965 & U3964 & U3963 & U3962); 
assign U3221 = ~(U3961 & U3960 & U3959 & U3958); 
assign U3275 = ~(U4237 & U2447); 
assign U3379 = ~(U5478 & U5477 & U7616); 
assign U3386 = ~(U4187 & U4465 & U4222); 
assign U3387 = ~(U2449 & U2447); 
assign U3397 = ~(U4241 & U3265); 
assign U3407 = ~(U4194 & U4465); 
assign U3414 = ~(U4237 & U3874 & U2452 & STATE2_REG_0__SCAN_IN); 
assign U3415 = ~(U3854 & U2447); 
assign U3421 = ~(U4194 & U3258); 
assign U3434 = ~(U4219 & U4388 & U4238); 
assign U3435 = ~(U4219 & U3265 & U4238); 
assign U3556 = U4365 & U4196; 
assign U3566 = U4237 & U3270; 
assign U3724 = U5459 & U5460; 
assign U3744 = U5551 & U5549; 
assign U3855 = U4196 & U2368; 
assign U3957 = U4223 & U4194; 
assign U3990 = U6737 & U6736; 
assign U4014 = U6846 & U6845; 
assign U4019 = U6891 & U6890 & U6889 & U6888; 
assign U4020 = U6895 & U6894 & U6893 & U6892; 
assign U4023 = U6909 & U6908 & U6907 & U6906; 
assign U4024 = U6913 & U6912 & U6911 & U6910; 
assign U4027 = U6940 & U6939 & U6938 & U6937; 
assign U4028 = U6944 & U6943 & U6942 & U6941; 
assign U4031 = U6957 & U6956 & U6955 & U6954; 
assign U4032 = U6961 & U6960 & U6959 & U6958; 
assign U4035 = U6974 & U6973 & U6972 & U6971; 
assign U4036 = U6978 & U6977 & U6976 & U6975; 
assign U4039 = U6991 & U6990 & U6989 & U6988; 
assign U4040 = U7602 & U6994 & U6993 & U6992; 
assign U4043 = U7006 & U7005 & U7004 & U7003; 
assign U4044 = U7010 & U7009 & U7008 & U7007; 
assign U4047 = U7023 & U7022 & U7021 & U7020; 
assign U4048 = U7027 & U7026 & U7025 & U7024; 
assign U4050 = U7050 & STATE2_REG_0__SCAN_IN; 
assign U4111 = U7219 & U7218 & U7217 & U7216; 
assign U4112 = U7223 & U7222 & U7221 & U7220; 
assign U4115 = U7236 & U7235 & U7234 & U7233; 
assign U4116 = U7240 & U7239 & U7238 & U7237; 
assign U4119 = U7253 & U7252 & U7251 & U7250; 
assign U4120 = U7257 & U7256 & U7255 & U7254; 
assign U4123 = U7270 & U7269 & U7268 & U7267; 
assign U4124 = U7607 & U7273 & U7272 & U7271; 
assign U4127 = U7285 & U7284 & U7283 & U7282; 
assign U4128 = U7289 & U7288 & U7287 & U7286; 
assign U4131 = U7302 & U7301 & U7300 & U7299; 
assign U4132 = U7306 & U7305 & U7304 & U7303; 
assign U4135 = U7319 & U7318 & U7317 & U7316; 
assign U4136 = U7323 & U7322 & U7321 & U7320; 
assign U4139 = U7336 & U7335 & U7334 & U7333; 
assign U4140 = U7340 & U7339 & U7338 & U7337; 
assign U4151 = U7361 & STATE2_REG_0__SCAN_IN; 
assign U4152 = U7363 & U2603; 
assign U4155 = U7377 & U7376 & U7375; 
assign U4185 = ~U3383; 
assign U4189 = ~U3409; 
assign U4244 = ~U3278; 
assign U4250 = ~U3273; 
assign U4251 = ~(U4224 & U4387); 
assign U4252 = ~U3398; 
assign U4489 = ~(U4488 & U3244); 
assign U4492 = ~(U4184 & U3273); 
assign U4773 = ~(U4767 & STATE2_REG_2__SCAN_IN); 
assign U4888 = ~(U4882 & STATE2_REG_2__SCAN_IN); 
assign U5001 = ~(U4996 & STATE2_REG_2__SCAN_IN); 
assign U5116 = ~(U5110 & STATE2_REG_2__SCAN_IN); 
assign U5231 = ~(U5225 & STATE2_REG_2__SCAN_IN); 
assign U5346 = ~(U5340 & STATE2_REG_2__SCAN_IN); 
assign U5449 = ~U3410; 
assign U5452 = ~U3231; 
assign U5456 = ~(U4196 & U5450); 
assign U5480 = ~(U5479 & U4159); 
assign U5484 = ~(U4196 & U5450); 
assign U5486 = ~(U5483 & U3258); 
assign U5488 = ~(U4178 & U3231); 
assign U6352 = ~(U4237 & STATE2_REG_2__SCAN_IN); 
assign U6593 = ~(U4196 & U6592); 
assign U6603 = ~(U3956 & U3278); 
assign U6735 = ~(U4176 & EAX_REG_9__SCAN_IN); 
assign U6738 = ~(U4176 & EAX_REG_8__SCAN_IN); 
assign U6741 = ~(U4176 & EAX_REG_7__SCAN_IN); 
assign U6744 = ~(U4176 & EAX_REG_6__SCAN_IN); 
assign U6748 = ~(U4176 & EAX_REG_5__SCAN_IN); 
assign U6752 = ~(U4176 & EAX_REG_4__SCAN_IN); 
assign U6755 = ~(U2353 & INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign U6756 = ~(U4176 & EAX_REG_31__SCAN_IN); 
assign U6760 = ~(U4176 & EAX_REG_30__SCAN_IN); 
assign U6764 = ~(U4176 & EAX_REG_3__SCAN_IN); 
assign U6767 = ~(U2353 & INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign U6769 = ~(U4176 & EAX_REG_29__SCAN_IN); 
assign U6773 = ~(U4176 & EAX_REG_28__SCAN_IN); 
assign U6777 = ~(U4176 & EAX_REG_27__SCAN_IN); 
assign U6781 = ~(U4176 & EAX_REG_26__SCAN_IN); 
assign U6785 = ~(U4176 & EAX_REG_25__SCAN_IN); 
assign U6789 = ~(U4176 & EAX_REG_24__SCAN_IN); 
assign U6793 = ~(U4176 & EAX_REG_23__SCAN_IN); 
assign U6797 = ~(U4176 & EAX_REG_22__SCAN_IN); 
assign U6801 = ~(U4176 & EAX_REG_21__SCAN_IN); 
assign U6805 = ~(U4176 & EAX_REG_20__SCAN_IN); 
assign U6809 = ~(U4176 & EAX_REG_2__SCAN_IN); 
assign U6812 = ~(U2353 & INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign U6814 = ~(U4176 & EAX_REG_19__SCAN_IN); 
assign U6818 = ~(U4176 & EAX_REG_18__SCAN_IN); 
assign U6822 = ~(U4176 & EAX_REG_17__SCAN_IN); 
assign U6826 = ~(U4176 & EAX_REG_16__SCAN_IN); 
assign U6829 = ~(U4176 & EAX_REG_15__SCAN_IN); 
assign U6832 = ~(U4176 & EAX_REG_14__SCAN_IN); 
assign U6835 = ~(U4176 & EAX_REG_13__SCAN_IN); 
assign U6838 = ~(U4176 & EAX_REG_12__SCAN_IN); 
assign U6841 = ~(U4176 & EAX_REG_11__SCAN_IN); 
assign U6844 = ~(U4176 & EAX_REG_10__SCAN_IN); 
assign U6848 = ~(U4176 & EAX_REG_1__SCAN_IN); 
assign U6851 = ~(U2353 & INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U6853 = ~(U4176 & EAX_REG_0__SCAN_IN); 
assign U6856 = ~(U2353 & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U7072 = ~(U4061 & U4179); 
assign U7077 = ~(U4177 & STATE2_REG_0__SCAN_IN); 
assign U7342 = ~(U4219 & U2354 & U4222); 
assign U7348 = ~(U4196 & U7076); 
assign U7349 = ~(U4148 & U4196); 
assign U7359 = ~(SUB_450_U21 & U2354); 
assign U7370 = ~(R2238_U21 & U4180); 
assign U7380 = ~(U7379 & INSTADDRPOINTER_REG_9__SCAN_IN); 
assign U7381 = ~(U7378 & EBX_REG_9__SCAN_IN); 
assign U7382 = ~(U7379 & INSTADDRPOINTER_REG_8__SCAN_IN); 
assign U7383 = ~(U7378 & EBX_REG_8__SCAN_IN); 
assign U7384 = ~(U7379 & INSTADDRPOINTER_REG_7__SCAN_IN); 
assign U7385 = ~(U7378 & EBX_REG_7__SCAN_IN); 
assign U7386 = ~(U7379 & INSTADDRPOINTER_REG_6__SCAN_IN); 
assign U7387 = ~(U7378 & EBX_REG_6__SCAN_IN); 
assign U7388 = ~(U7379 & INSTADDRPOINTER_REG_5__SCAN_IN); 
assign U7389 = ~(U7378 & EBX_REG_5__SCAN_IN); 
assign U7390 = ~(U7379 & INSTADDRPOINTER_REG_4__SCAN_IN); 
assign U7391 = ~(U7378 & EBX_REG_4__SCAN_IN); 
assign U7392 = ~(U7379 & INSTADDRPOINTER_REG_31__SCAN_IN); 
assign U7393 = ~(U7378 & EBX_REG_31__SCAN_IN); 
assign U7394 = ~(U7379 & INSTADDRPOINTER_REG_30__SCAN_IN); 
assign U7395 = ~(U7378 & EBX_REG_30__SCAN_IN); 
assign U7396 = ~(U7379 & INSTADDRPOINTER_REG_3__SCAN_IN); 
assign U7397 = ~(U7378 & EBX_REG_3__SCAN_IN); 
assign U7398 = ~(U7379 & INSTADDRPOINTER_REG_29__SCAN_IN); 
assign U7399 = ~(U7378 & EBX_REG_29__SCAN_IN); 
assign U7400 = ~(U7379 & INSTADDRPOINTER_REG_28__SCAN_IN); 
assign U7401 = ~(U7378 & EBX_REG_28__SCAN_IN); 
assign U7402 = ~(U7379 & INSTADDRPOINTER_REG_27__SCAN_IN); 
assign U7403 = ~(U7378 & EBX_REG_27__SCAN_IN); 
assign U7404 = ~(U7379 & INSTADDRPOINTER_REG_26__SCAN_IN); 
assign U7405 = ~(U7378 & EBX_REG_26__SCAN_IN); 
assign U7406 = ~(U7379 & INSTADDRPOINTER_REG_25__SCAN_IN); 
assign U7407 = ~(U7378 & EBX_REG_25__SCAN_IN); 
assign U7408 = ~(U7379 & INSTADDRPOINTER_REG_24__SCAN_IN); 
assign U7409 = ~(U7378 & EBX_REG_24__SCAN_IN); 
assign U7410 = ~(U7379 & INSTADDRPOINTER_REG_23__SCAN_IN); 
assign U7411 = ~(U7378 & EBX_REG_23__SCAN_IN); 
assign U7412 = ~(U7379 & INSTADDRPOINTER_REG_22__SCAN_IN); 
assign U7413 = ~(U7378 & EBX_REG_22__SCAN_IN); 
assign U7414 = ~(U7379 & INSTADDRPOINTER_REG_21__SCAN_IN); 
assign U7415 = ~(U7378 & EBX_REG_21__SCAN_IN); 
assign U7416 = ~(U7379 & INSTADDRPOINTER_REG_20__SCAN_IN); 
assign U7417 = ~(U7378 & EBX_REG_20__SCAN_IN); 
assign U7418 = ~(U7379 & INSTADDRPOINTER_REG_2__SCAN_IN); 
assign U7419 = ~(U7378 & EBX_REG_2__SCAN_IN); 
assign U7420 = ~(U7379 & INSTADDRPOINTER_REG_19__SCAN_IN); 
assign U7421 = ~(U7378 & EBX_REG_19__SCAN_IN); 
assign U7422 = ~(U7379 & INSTADDRPOINTER_REG_18__SCAN_IN); 
assign U7423 = ~(U7378 & EBX_REG_18__SCAN_IN); 
assign U7424 = ~(U7379 & INSTADDRPOINTER_REG_17__SCAN_IN); 
assign U7425 = ~(U7378 & EBX_REG_17__SCAN_IN); 
assign U7426 = ~(U7379 & INSTADDRPOINTER_REG_16__SCAN_IN); 
assign U7427 = ~(U7378 & EBX_REG_16__SCAN_IN); 
assign U7428 = ~(U7379 & INSTADDRPOINTER_REG_15__SCAN_IN); 
assign U7429 = ~(U7378 & EBX_REG_15__SCAN_IN); 
assign U7430 = ~(U7379 & INSTADDRPOINTER_REG_14__SCAN_IN); 
assign U7431 = ~(U7378 & EBX_REG_14__SCAN_IN); 
assign U7432 = ~(U7379 & INSTADDRPOINTER_REG_13__SCAN_IN); 
assign U7433 = ~(U7378 & EBX_REG_13__SCAN_IN); 
assign U7434 = ~(U7379 & INSTADDRPOINTER_REG_12__SCAN_IN); 
assign U7435 = ~(U7378 & EBX_REG_12__SCAN_IN); 
assign U7436 = ~(U7379 & INSTADDRPOINTER_REG_11__SCAN_IN); 
assign U7437 = ~(U7378 & EBX_REG_11__SCAN_IN); 
assign U7438 = ~(U7379 & INSTADDRPOINTER_REG_10__SCAN_IN); 
assign U7439 = ~(U7378 & EBX_REG_10__SCAN_IN); 
assign U7440 = ~(U7379 & INSTADDRPOINTER_REG_1__SCAN_IN); 
assign U7441 = ~(U7378 & EBX_REG_1__SCAN_IN); 
assign U7442 = ~(U7379 & INSTADDRPOINTER_REG_0__SCAN_IN); 
assign U7443 = ~(U7378 & EBX_REG_0__SCAN_IN); 
assign U7463 = ~(U4224 & STATE2_REG_0__SCAN_IN); 
assign U7477 = ~(U4224 & STATE2_REG_0__SCAN_IN); 
assign U7481 = ~U3266; 
assign U7618 = ~(U4196 & U7478); 
assign U7688 = ~(U5455 & U4159); 
assign R2027_U51 = ~(R2027_U142 & R2027_U141); 
assign R2027_U52 = ~(R2027_U144 & R2027_U143); 
assign R2027_U113 = ~R2027_U22; 
assign R2027_U140 = ~R2027_U110; 
assign R2027_U200 = ~(R2027_U22 & INSTADDRPOINTER_REG_11__SCAN_IN); 
assign R2027_U201 = ~(R2027_U110 & INSTADDRPOINTER_REG_10__SCAN_IN); 
assign R2337_U78 = ~(R2337_U189 & R2337_U188); 
assign R2337_U79 = ~(R2337_U191 & R2337_U190); 
assign R2337_U115 = ~R2337_U103; 
assign R2337_U116 = ~R2337_U23; 
assign R2337_U184 = ~(R2337_U23 & PHYADDRPOINTER_REG_14__SCAN_IN); 
assign R2337_U186 = ~(R2337_U103 & PHYADDRPOINTER_REG_13__SCAN_IN); 
assign R2099_U5 = ~U4177; 
assign R2099_U6 = ~U2678; 
assign R2099_U146 = U4178 | U4177; 
assign R2099_U148 = ~(U4177 & U4178); 
assign R2099_U345 = ~(U4177 & R2099_U4); 
assign R2167_U23 = ~U2722; 
assign R2096_U65 = ~(R2096_U130 & R2096_U129); 
assign R2096_U98 = ~R2096_U14; 
assign R2096_U127 = ~(R2096_U14 & REIP_REG_7__SCAN_IN); 
assign R2238_U16 = ~(R2238_U41 & R2238_U40); 
assign R2238_U55 = ~(R2238_U38 & R2238_U54); 
assign SUB_450_U16 = ~(SUB_450_U41 & SUB_450_U40); 
assign SUB_450_U55 = ~(SUB_450_U38 & SUB_450_U54); 
assign ADD_405_U66 = ~(ADD_405_U134 & ADD_405_U133); 
assign ADD_405_U101 = ~ADD_405_U14; 
assign ADD_405_U131 = ~(ADD_405_U14 & INSTADDRPOINTER_REG_7__SCAN_IN); 
assign ADD_515_U65 = ~(ADD_515_U130 & ADD_515_U129); 
assign ADD_515_U98 = ~ADD_515_U14; 
assign ADD_515_U127 = ~(ADD_515_U14 & INSTADDRPOINTER_REG_7__SCAN_IN); 
assign U2355 = U3221 & U2450; 
assign U2609 = ~(U6744 & U3993); 
assign U2610 = ~(U6741 & U3992); 
assign U2611 = ~(U6738 & U3991); 
assign U2612 = ~(U6735 & U3990); 
assign U2613 = ~(U6844 & U4014); 
assign U2679 = ~(U7393 & U7392); 
assign U2680 = ~(U7395 & U7394); 
assign U2681 = ~(U7399 & U7398); 
assign U2682 = ~(U7401 & U7400); 
assign U2683 = ~(U7403 & U7402); 
assign U2684 = ~(U7405 & U7404); 
assign U2685 = ~(U7407 & U7406); 
assign U2686 = ~(U7409 & U7408); 
assign U2687 = ~(U7411 & U7410); 
assign U2688 = ~(U7413 & U7412); 
assign U2689 = ~(U7415 & U7414); 
assign U2690 = ~(U7417 & U7416); 
assign U2691 = ~(U7421 & U7420); 
assign U2692 = ~(U7423 & U7422); 
assign U2693 = ~(U7425 & U7424); 
assign U2694 = ~(U7427 & U7426); 
assign U2695 = ~(U7429 & U7428); 
assign U2696 = ~(U7431 & U7430); 
assign U2697 = ~(U7433 & U7432); 
assign U2698 = ~(U7435 & U7434); 
assign U2699 = ~(U7437 & U7436); 
assign U2700 = ~(U7439 & U7438); 
assign U2701 = ~(U7381 & U7380); 
assign U2702 = ~(U7383 & U7382); 
assign U2703 = ~(U7385 & U7384); 
assign U2704 = ~(U7387 & U7386); 
assign U2705 = ~(U7389 & U7388); 
assign U2706 = ~(U7391 & U7390); 
assign U2707 = ~(U7397 & U7396); 
assign U2708 = ~(U7419 & U7418); 
assign U2709 = ~(U7441 & U7440); 
assign U2710 = ~(U7443 & U7442); 
assign U2714 = ~(U7374 & U7373 & U4154 & U3421); 
assign U3232 = ~(U7074 & U5452); 
assign U3279 = ~(U4244 & U2431); 
assign U3428 = ~U3221; 
assign U3433 = ~(U4185 & U4222); 
assign U3730 = U5484 & U3380; 
assign U3731 = U5486 & U5485; 
assign U3733 = U4251 & U3384; 
assign U3994 = U6748 & U3995; 
assign U3996 = U6752 & U6753; 
assign U3998 = U6764 & U6765; 
assign U4009 = U6809 & U6810; 
assign U4015 = U6848 & U6849; 
assign U4055 = U4244 & STATE2_REG_0__SCAN_IN; 
assign U4099 = U7077 & U3414; 
assign U4146 = U4145 & U7348; 
assign U4150 = U7359 & U2603; 
assign U4153 = U7370 & U7371; 
assign U4181 = ~U3421; 
assign U4182 = ~U3407; 
assign U4190 = ~U3415; 
assign U4192 = ~U3414; 
assign U4193 = ~(U3873 & U4177 & U4185); 
assign U4200 = ~U3434; 
assign U4201 = ~U3435; 
assign U4202 = ~U3387; 
assign U4203 = ~U3275; 
assign U4205 = ~(U3566 & U2431); 
assign U4206 = ~U3386; 
assign U4254 = ~U3397; 
assign U4493 = ~(U4492 & U3567); 
assign U5454 = ~(U5453 & U3270 & U5452); 
assign U5508 = ~(U2431 & U4237); 
assign U5553 = ~(U4250 & U4196); 
assign U5554 = ~(U4244 & U2389); 
assign U5556 = ~(U4252 & U4482); 
assign U6594 = ~(U3952 & U6593); 
assign U6840 = ~(R2337_U78 & U2352); 
assign U6843 = ~(R2337_U79 & U2352); 
assign U6896 = ~(U4020 & U4019 & U4018 & U4017); 
assign U6914 = ~(U4024 & U4023 & U4022 & U4021); 
assign U6945 = ~(U4028 & U4027 & U4026 & U4025); 
assign U6962 = ~(U4032 & U4031 & U4030 & U4029); 
assign U6979 = ~(U4036 & U4035 & U4034 & U4033); 
assign U7011 = ~(U4044 & U4043 & U4042 & U4041); 
assign U7028 = ~(U4048 & U4047 & U4046 & U4045); 
assign U7035 = ~(U4194 & U3221); 
assign U7037 = ~(U4194 & U3220); 
assign U7039 = ~(U4194 & U3219); 
assign U7041 = ~(U4194 & U3218); 
assign U7042 = ~(U4194 & U3217); 
assign U7044 = ~(U4194 & U3216); 
assign U7046 = ~(U4194 & U3215); 
assign U7048 = ~(U4194 & U3214); 
assign U7049 = ~(U3221 & U4388); 
assign U7051 = ~(U3415 & U3414); 
assign U7073 = ~(U7072 & U3409); 
assign U7224 = ~(U4112 & U4111 & U4110 & U4109); 
assign U7241 = ~(U4116 & U4115 & U4114 & U4113); 
assign U7258 = ~(U4120 & U4119 & U4118 & U4117); 
assign U7290 = ~(U4128 & U4127 & U4126 & U4125); 
assign U7307 = ~(U4132 & U4131 & U4130 & U4129); 
assign U7324 = ~(U4136 & U4135 & U4134 & U4133); 
assign U7341 = ~(U4140 & U4139 & U4138 & U4137); 
assign U7344 = ~(U3383 & U3397); 
assign U7351 = ~(U3407 & U3421 & U4183 & U7350 & U7349); 
assign U7369 = ~(U3407 & U7368); 
assign U7459 = ~(U7072 & U3409); 
assign U7464 = ~(U4252 & STATE2_REG_0__SCAN_IN); 
assign U7484 = ~(U3722 & U7481); 
assign U7495 = ~(U3747 & U7481); 
assign U7593 = ~(U3855 & U7481); 
assign U7595 = ~(U4196 & U7481); 
assign U7597 = ~(U3266 & U3387); 
assign U7598 = ~(U3742 & U7481); 
assign U7603 = ~(U4040 & U4039 & U4038 & U4037); 
assign U7608 = ~(U4124 & U4123 & U4122 & U4121); 
assign U7617 = ~U3379; 
assign U7620 = ~(U7619 & U7618); 
assign R2027_U25 = ~(R2027_U86 & R2027_U113); 
assign R2027_U109 = ~(R2027_U113 & INSTADDRPOINTER_REG_11__SCAN_IN); 
assign R2027_U199 = ~(R2027_U113 & R2027_U21); 
assign R2027_U202 = ~(R2027_U140 & R2027_U19); 
assign R2337_U26 = ~(R2337_U85 & R2337_U116); 
assign R2337_U102 = ~(R2337_U116 & PHYADDRPOINTER_REG_14__SCAN_IN); 
assign R2337_U185 = ~(R2337_U116 & R2337_U25); 
assign R2337_U187 = ~(R2337_U115 & R2337_U21); 
assign R2099_U346 = ~(U4178 & R2099_U5); 
assign SUB_357_U6 = ~U3220; 
assign SUB_357_U7 = ~U3215; 
assign SUB_357_U8 = ~U3221; 
assign SUB_357_U9 = ~U3219; 
assign SUB_357_U10 = ~U3214; 
assign SUB_357_U11 = ~U3217; 
assign SUB_357_U12 = ~U3216; 
assign SUB_357_U13 = ~U3218; 
assign R2096_U16 = ~(R2096_U98 & REIP_REG_7__SCAN_IN); 
assign R2096_U128 = ~(R2096_U98 & R2096_U15); 
assign R2238_U20 = ~(R2238_U56 & R2238_U55); 
assign R2238_U42 = ~R2238_U16; 
assign R2238_U51 = ~(R2238_U23 & R2238_U16); 
assign SUB_450_U20 = ~(SUB_450_U56 & SUB_450_U55); 
assign SUB_450_U42 = ~SUB_450_U16; 
assign SUB_450_U51 = ~(SUB_450_U23 & SUB_450_U16); 
assign ADD_371_U4 = ~U3214; 
assign ADD_371_U7 = ~U3215; 
assign ADD_371_U8 = ~U3217; 
assign ADD_371_U10 = ~U3218; 
assign ADD_371_U12 = ~U3219; 
assign ADD_371_U14 = ~U3221; 
assign ADD_371_U15 = ~U3220; 
assign ADD_371_U16 = ~U3216; 
assign ADD_371_U22 = U3221 & U3220; 
assign ADD_371_U26 = ~(U3215 & U3214); 
assign ADD_371_U32 = ~(U3215 & U3214 & U3216); 
assign ADD_405_U16 = ~(ADD_405_U101 & INSTADDRPOINTER_REG_7__SCAN_IN); 
assign ADD_405_U132 = ~(ADD_405_U101 & ADD_405_U15); 
assign ADD_515_U16 = ~(ADD_515_U98 & INSTADDRPOINTER_REG_7__SCAN_IN); 
assign ADD_515_U128 = ~(ADD_515_U98 & ADD_515_U15); 
assign U2520 = U4207 & U3433; 
assign U2614 = ~(U6841 & U6842 & U6843); 
assign U2615 = ~(U6838 & U6839 & U6840); 
assign U2740 = U7051 & INSTQUEUERD_ADDR_REG_4__SCAN_IN; 
assign U2745 = ~(U7036 & U7035); 
assign U2746 = ~(U7038 & U7037); 
assign U2747 = ~(U7040 & U7039); 
assign U2748 = ~(U7604 & U7041); 
assign U2749 = ~(U7043 & U7042); 
assign U2750 = ~(U7045 & U7044); 
assign U2752 = ~(U4050 & U7048 & U7049); 
assign U2753 = U6945 & U6897; 
assign U2754 = U6962 & U6897; 
assign U2755 = U6979 & U6897; 
assign U2756 = U7603 & U6897; 
assign U2757 = U7011 & U6897; 
assign U2758 = U7028 & U6897; 
assign U2759 = U6897 & U6896; 
assign U2760 = U6914 & U6897; 
assign U3408 = ~(U4182 & U2431); 
assign U3430 = ~(U2450 & U3428); 
assign U3438 = ~(U4242 & U4254); 
assign U3568 = U4205 & U3387; 
assign U3723 = U7484 & U4205; 
assign U3732 = U5488 & U7615 & U3730 & U3731; 
assign U3748 = U3275 & U4205 & U3435; 
assign U3749 = U5554 & U7495; 
assign U4199 = ~U3433; 
assign U4204 = ~U3279; 
assign U4227 = ~(U4465 & U7369); 
assign U5457 = ~(U3721 & U7597); 
assign U5481 = ~(U7617 & U5480); 
assign U5489 = ~(U3279 & U4205); 
assign U5492 = ~(U4206 & U3425); 
assign U5493 = ~(U4202 & U3429); 
assign U5501 = ~(U4202 & U3443); 
assign U5509 = ~(U3279 & U5508); 
assign U5512 = ~(U4202 & U3252); 
assign U5555 = ~(U4254 & U4238); 
assign U6138 = ~(U4242 & U4185 & U4182); 
assign U6595 = ~(U6594 & STATE2_REG_0__SCAN_IN); 
assign U6596 = ~(U4181 & U3259); 
assign U6878 = ~(ADD_371_U4 & U4196); 
assign U6916 = ~(U2355 & SUB_357_U8); 
assign U6918 = ~(SUB_357_U6 & U2355); 
assign U6920 = ~(SUB_357_U9 & U2355); 
assign U6922 = ~(SUB_357_U13 & U2355); 
assign U6924 = ~(SUB_357_U11 & U2355); 
assign U6927 = ~(SUB_357_U12 & U2355); 
assign U7030 = ~(SUB_357_U7 & U2355); 
assign U7033 = ~(SUB_357_U10 & U2355); 
assign U7075 = ~U3232; 
assign U7078 = ~(U4055 & U3232); 
assign U7345 = ~(U4222 & U7344); 
assign U7356 = ~(R2238_U20 & U7351); 
assign U7357 = ~(SUB_450_U20 & U2354); 
assign U7358 = ~(R2238_U21 & U7351); 
assign U7360 = ~(R2238_U22 & U7351); 
assign U7362 = ~(R2238_U7 & U7351); 
assign U7366 = ~(R2238_U20 & U4180); 
assign U7461 = ~(U4200 & STATE2_REG_0__SCAN_IN); 
assign U7462 = ~(U4201 & STATE2_REG_0__SCAN_IN); 
assign U7465 = ~(U7620 & STATE2_REG_0__SCAN_IN); 
assign U7468 = ~(U7620 & STATE2_REG_0__SCAN_IN); 
assign U7474 = ~(U5479 & U4159 & U4182); 
assign U7476 = ~(U4182 & U3379); 
assign U7492 = ~(U7481 & U7073); 
assign U7493 = ~(U7481 & U7459); 
assign U7594 = ~(U7593 & U3415); 
assign U7596 = ~(U7595 & U3434); 
assign U7599 = ~(U3743 & U7598); 
assign U7687 = ~(U4420 & U5454); 
assign U7705 = ~(U4206 & U3388); 
assign U7713 = ~(U4202 & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign R2027_U80 = ~(R2027_U200 & R2027_U199); 
assign R2027_U81 = ~(R2027_U202 & R2027_U201); 
assign R2027_U119 = ~R2027_U25; 
assign R2027_U139 = ~R2027_U109; 
assign R2027_U196 = ~(R2027_U25 & INSTADDRPOINTER_REG_13__SCAN_IN); 
assign R2027_U197 = ~(R2027_U109 & INSTADDRPOINTER_REG_12__SCAN_IN); 
assign R2358_U164 = ~U2612; 
assign R2358_U166 = ~U2610; 
assign R2358_U167 = ~U2609; 
assign R2358_U174 = ~U2611; 
assign R2358_U181 = ~U2613; 
assign R2358_U441 = ~(U2612 & R2358_U22); 
assign R2358_U449 = ~(U2610 & R2358_U22); 
assign R2358_U452 = ~(U2610 & R2358_U22); 
assign R2358_U454 = ~(U2609 & R2358_U22); 
assign R2358_U487 = ~(U2611 & R2358_U22); 
assign R2358_U489 = ~(U2611 & R2358_U22); 
assign R2358_U510 = ~(U2613 & R2358_U22); 
assign R2358_U517 = ~(U2613 & R2358_U22); 
assign R2337_U76 = ~(R2337_U185 & R2337_U184); 
assign R2337_U77 = ~(R2337_U187 & R2337_U186); 
assign R2337_U117 = ~R2337_U102; 
assign R2337_U118 = ~R2337_U26; 
assign R2337_U180 = ~(R2337_U26 & PHYADDRPOINTER_REG_16__SCAN_IN); 
assign R2337_U182 = ~(R2337_U102 & PHYADDRPOINTER_REG_15__SCAN_IN); 
assign R2144_U12 = ~U2355; 
assign R2099_U98 = ~(R2099_U346 & R2099_U345); 
assign R2099_U99 = ~U2702; 
assign R2099_U100 = ~U2710; 
assign R2099_U101 = ~U2709; 
assign R2099_U102 = ~U2708; 
assign R2099_U103 = ~U2707; 
assign R2099_U104 = ~U2706; 
assign R2099_U105 = ~U2705; 
assign R2099_U106 = ~U2704; 
assign R2099_U107 = ~U2703; 
assign R2099_U108 = ~U2701; 
assign R2099_U113 = ~U2682; 
assign R2099_U114 = ~U2683; 
assign R2099_U115 = ~U2684; 
assign R2099_U116 = ~U2685; 
assign R2099_U117 = ~U2686; 
assign R2099_U118 = ~U2687; 
assign R2099_U119 = ~U2688; 
assign R2099_U120 = ~U2689; 
assign R2099_U121 = ~U2690; 
assign R2099_U122 = ~U2691; 
assign R2099_U123 = ~U2692; 
assign R2099_U124 = ~U2700; 
assign R2099_U125 = ~U2699; 
assign R2099_U126 = ~U2698; 
assign R2099_U127 = ~U2697; 
assign R2099_U128 = ~U2696; 
assign R2099_U129 = ~U2695; 
assign R2099_U130 = ~U2694; 
assign R2099_U131 = ~U2693; 
assign R2099_U132 = ~U2680; 
assign R2099_U133 = ~U2681; 
assign R2099_U134 = ~U2679; 
assign R2099_U183 = ~(U2702 & R2099_U4); 
assign R2099_U186 = ~(U2710 & R2099_U4); 
assign R2099_U189 = ~(U2709 & R2099_U4); 
assign R2099_U192 = ~(U2708 & R2099_U4); 
assign R2099_U195 = ~(U2707 & R2099_U4); 
assign R2099_U198 = ~(U2706 & R2099_U4); 
assign R2099_U201 = ~(U2705 & R2099_U4); 
assign R2099_U204 = ~(U2704 & R2099_U4); 
assign R2099_U207 = ~(U2703 & R2099_U4); 
assign R2099_U210 = ~(U2701 & R2099_U4); 
assign R2099_U227 = ~(U2682 & R2099_U4); 
assign R2099_U230 = ~(U2683 & R2099_U4); 
assign R2099_U233 = ~(U2684 & R2099_U4); 
assign R2099_U236 = ~(U2685 & R2099_U4); 
assign R2099_U239 = ~(U2686 & R2099_U4); 
assign R2099_U242 = ~(U2687 & R2099_U4); 
assign R2099_U245 = ~(U2688 & R2099_U4); 
assign R2099_U248 = ~(U2689 & R2099_U4); 
assign R2099_U251 = ~(U2690 & R2099_U4); 
assign R2099_U254 = ~(U2691 & R2099_U4); 
assign R2099_U257 = ~(U2692 & R2099_U4); 
assign R2099_U260 = ~(U2700 & R2099_U4); 
assign R2099_U263 = ~(U2699 & R2099_U4); 
assign R2099_U266 = ~(U2698 & R2099_U4); 
assign R2099_U269 = ~(U2697 & R2099_U4); 
assign R2099_U272 = ~(U2696 & R2099_U4); 
assign R2099_U275 = ~(U2695 & R2099_U4); 
assign R2099_U278 = ~(U2694 & R2099_U4); 
assign R2099_U281 = ~(U2693 & R2099_U4); 
assign R2099_U284 = ~(U2680 & R2099_U4); 
assign R2099_U287 = ~(U2681 & R2099_U4); 
assign R2099_U290 = ~(U2679 & R2099_U4); 
assign R2167_U7 = ~U2714; 
assign R2096_U64 = ~(R2096_U128 & R2096_U127); 
assign R2096_U99 = ~R2096_U16; 
assign R2096_U125 = ~(R2096_U16 & REIP_REG_8__SCAN_IN); 
assign R2238_U44 = ~(R2238_U42 & R2238_U43); 
assign R2238_U50 = ~(R2238_U49 & R2238_U42); 
assign SUB_450_U44 = ~(SUB_450_U42 & SUB_450_U43); 
assign SUB_450_U50 = ~(SUB_450_U49 & SUB_450_U42); 
assign ADD_371_U24 = ~(ADD_371_U16 & ADD_371_U26); 
assign ADD_371_U43 = ~(U3215 & ADD_371_U4); 
assign ADD_371_U44 = ~(U3214 & ADD_371_U7); 
assign ADD_405_U65 = ~(ADD_405_U132 & ADD_405_U131); 
assign ADD_405_U102 = ~ADD_405_U16; 
assign ADD_405_U129 = ~(ADD_405_U16 & INSTADDRPOINTER_REG_8__SCAN_IN); 
assign ADD_515_U64 = ~(ADD_515_U128 & ADD_515_U127); 
assign ADD_515_U99 = ~ADD_515_U16; 
assign ADD_515_U125 = ~(ADD_515_U16 & INSTADDRPOINTER_REG_8__SCAN_IN); 
assign U2518 = U7688 & U7687 & U5456; 
assign U2606 = U7492 & U3414; 
assign U2712 = ~(U7367 & U7366); 
assign U2713 = ~(U4153 & U4227); 
assign U2715 = ~(U4227 & U4155); 
assign U2719 = ~(U4150 & U7358); 
assign U2720 = ~(U4151 & U7360); 
assign U2721 = ~(U4152 & U7362); 
assign U3412 = ~(U4204 & STATE2_REG_0__SCAN_IN); 
assign U3734 = U3398 & U3275 & U3733 & U2520 & U3266; 
assign U3736 = U5493 & U5492; 
assign U3745 = U3385 & U3386 & U5555; 
assign U3953 = U6596 & U3285; 
assign U4049 = U7047 & U3430; 
assign U4062 = U7078 & U7077; 
assign U4064 = U7463 & U7464 & U7462; 
assign U4103 = U7474 & U7468 & U7464 & U7462; 
assign U4105 = U7078 & U7077; 
assign U4107 = U7463 & U7464 & U7462; 
assign U4143 = U7345 & U7346 & U4251; 
assign U4149 = U7357 & STATE2_REG_0__SCAN_IN; 
assign U4188 = ~U3408; 
assign U4195 = ~U3430; 
assign U4494 = ~(U3568 & U4493); 
assign U5490 = ~(U3728 & U5489); 
assign U5510 = ~(U5507 & U5509); 
assign U6834 = ~(R2337_U76 & U2352); 
assign U6837 = ~(R2337_U77 & U2352); 
assign U7079 = ~U3438; 
assign U7080 = ~(U3438 & U5480 & U7617); 
assign U7343 = ~(U4141 & U7075); 
assign U7460 = ~(U4199 & STATE2_REG_0__SCAN_IN); 
assign U7485 = ~(U3723 & U5457); 
assign U7496 = ~(U3749 & U5553 & U3748); 
assign U7694 = ~(U4465 & U5481); 
assign U7704 = ~(U5499 & U5489); 
assign U7714 = ~(U5509 & U3253); 
assign R2027_U27 = ~(R2027_U87 & R2027_U119); 
assign R2027_U108 = ~(R2027_U119 & INSTADDRPOINTER_REG_13__SCAN_IN); 
assign R2027_U195 = ~(R2027_U119 & R2027_U24); 
assign R2027_U198 = ~(R2027_U139 & R2027_U20); 
assign R2358_U182 = ~U2614; 
assign R2358_U184 = ~U2615; 
assign R2358_U440 = ~(U2352 & R2358_U164); 
assign R2358_U448 = ~(U2352 & R2358_U166); 
assign R2358_U451 = ~(U2352 & R2358_U166); 
assign R2358_U453 = ~(U2352 & R2358_U167); 
assign R2358_U486 = ~(U2352 & R2358_U174); 
assign R2358_U488 = ~(U2352 & R2358_U174); 
assign R2358_U509 = ~(U2352 & R2358_U181); 
assign R2358_U512 = ~(U2614 & R2358_U22); 
assign R2358_U514 = ~(U2614 & R2358_U22); 
assign R2358_U516 = ~(U2352 & R2358_U181); 
assign R2358_U523 = ~(U2615 & R2358_U22); 
assign R2358_U530 = ~(U2615 & R2358_U22); 
assign R2337_U29 = ~(R2337_U86 & R2337_U118); 
assign R2337_U101 = ~(R2337_U118 & PHYADDRPOINTER_REG_16__SCAN_IN); 
assign R2337_U181 = ~(R2337_U118 & R2337_U28); 
assign R2337_U183 = ~(R2337_U117 & R2337_U24); 
assign R2182_U12 = ~U2740; 
assign R2144_U13 = ~U2750; 
assign R2144_U15 = ~U2752; 
assign R2144_U16 = ~U2749; 
assign R2144_U17 = ~U2745; 
assign R2144_U18 = ~U2748; 
assign R2144_U20 = ~U2747; 
assign R2144_U22 = ~U2746; 
assign R2144_U76 = ~U2760; 
assign R2144_U77 = ~U2759; 
assign R2144_U85 = ~U2754; 
assign R2144_U86 = ~U2753; 
assign R2144_U87 = ~U2755; 
assign R2144_U88 = ~U2756; 
assign R2144_U89 = ~U2757; 
assign R2144_U90 = ~U2758; 
assign R2144_U203 = ~(U2760 & R2144_U12); 
assign R2144_U206 = ~(U2759 & R2144_U12); 
assign R2144_U221 = ~(U2754 & R2144_U12); 
assign R2144_U224 = ~(U2753 & R2144_U12); 
assign R2144_U227 = ~(U2755 & R2144_U12); 
assign R2144_U230 = ~(U2756 & R2144_U12); 
assign R2144_U233 = ~(U2757 & R2144_U12); 
assign R2144_U236 = ~(U2758 & R2144_U12); 
assign R2099_U182 = ~(U4178 & R2099_U99); 
assign R2099_U185 = ~(U4178 & R2099_U100); 
assign R2099_U188 = ~(U4178 & R2099_U101); 
assign R2099_U191 = ~(U4178 & R2099_U102); 
assign R2099_U194 = ~(U4178 & R2099_U103); 
assign R2099_U197 = ~(U4178 & R2099_U104); 
assign R2099_U200 = ~(U4178 & R2099_U105); 
assign R2099_U203 = ~(U4178 & R2099_U106); 
assign R2099_U206 = ~(U4178 & R2099_U107); 
assign R2099_U209 = ~(U4178 & R2099_U108); 
assign R2099_U226 = ~(U4178 & R2099_U113); 
assign R2099_U229 = ~(U4178 & R2099_U114); 
assign R2099_U232 = ~(U4178 & R2099_U115); 
assign R2099_U235 = ~(U4178 & R2099_U116); 
assign R2099_U238 = ~(U4178 & R2099_U117); 
assign R2099_U241 = ~(U4178 & R2099_U118); 
assign R2099_U244 = ~(U4178 & R2099_U119); 
assign R2099_U247 = ~(U4178 & R2099_U120); 
assign R2099_U250 = ~(U4178 & R2099_U121); 
assign R2099_U253 = ~(U4178 & R2099_U122); 
assign R2099_U256 = ~(U4178 & R2099_U123); 
assign R2099_U259 = ~(U4178 & R2099_U124); 
assign R2099_U262 = ~(U4178 & R2099_U125); 
assign R2099_U265 = ~(U4178 & R2099_U126); 
assign R2099_U268 = ~(U4178 & R2099_U127); 
assign R2099_U271 = ~(U4178 & R2099_U128); 
assign R2099_U274 = ~(U4178 & R2099_U129); 
assign R2099_U277 = ~(U4178 & R2099_U130); 
assign R2099_U280 = ~(U4178 & R2099_U131); 
assign R2099_U283 = ~(U4178 & R2099_U132); 
assign R2099_U286 = ~(U4178 & R2099_U133); 
assign R2099_U289 = ~(U4178 & R2099_U134); 
assign R2099_U347 = ~R2099_U98; 
assign R2096_U19 = ~(R2096_U99 & REIP_REG_8__SCAN_IN); 
assign R2096_U126 = ~(R2096_U99 & R2096_U17); 
assign R2238_U6 = ~(R2238_U45 & R2238_U44); 
assign R2238_U19 = ~(R2238_U51 & R2238_U50); 
assign SUB_450_U6 = ~(SUB_450_U45 & SUB_450_U44); 
assign SUB_450_U19 = ~(SUB_450_U51 & SUB_450_U50); 
assign ADD_371_U5 = ~(ADD_371_U24 & ADD_371_U32); 
assign ADD_371_U9 = ~(U3217 & ADD_371_U24); 
assign ADD_371_U21 = ~(ADD_371_U44 & ADD_371_U43); 
assign ADD_371_U27 = ~ADD_371_U24; 
assign ADD_371_U41 = ~(U3217 & ADD_371_U24); 
assign ADD_405_U19 = ~(ADD_405_U102 & INSTADDRPOINTER_REG_8__SCAN_IN); 
assign ADD_405_U130 = ~(ADD_405_U102 & ADD_405_U17); 
assign ADD_515_U19 = ~(ADD_515_U99 & INSTADDRPOINTER_REG_8__SCAN_IN); 
assign ADD_515_U126 = ~(ADD_515_U99 & ADD_515_U17); 
assign U2356 = R2238_U6 & U4180; 
assign U2616 = ~(U6835 & U6836 & U6837); 
assign U2617 = ~(U6832 & U6833 & U6834); 
assign U2718 = ~(U4149 & U7356); 
assign U2731 = ~(U2606 & U7342); 
assign U2751 = ~(U4049 & U7046); 
assign U3735 = U3736 & U5490; 
assign U3737 = U7705 & U7704 & U5501; 
assign U3738 = U5512 & U5510; 
assign U3746 = U2520 & U5556 & U3745; 
assign U3750 = U7496 & STATE2_REG_2__SCAN_IN; 
assign U4063 = U7460 & U3421 & U7461; 
assign U4065 = U2606 & U7465 & U4064; 
assign U4101 = U4100 & U7460 & U7461; 
assign U4106 = U7460 & U3421 & U7461; 
assign U4108 = U2608 & U7465 & U2606 & U4107; 
assign U4163 = U7714 & U7713; 
assign U4186 = ~U3412; 
assign U6597 = ~(U3953 & U6595); 
assign U6872 = ~(ADD_371_U5 & U4196); 
assign U6875 = ~(ADD_371_U21 & U4196); 
assign U6915 = ~(U4195 & U3221); 
assign U6917 = ~(U4195 & U3220); 
assign U6919 = ~(U4195 & U3219); 
assign U6921 = ~(U4195 & U3218); 
assign U6923 = ~(U4195 & U3217); 
assign U6926 = ~(U4195 & U3216); 
assign U7029 = ~(U4195 & U3215); 
assign U7032 = ~(U4195 & U3214); 
assign U7071 = ~(U3412 & U3408); 
assign U7081 = ~(U4182 & U7080); 
assign U7347 = ~(U7343 & U3258); 
assign U7352 = ~(R2238_U6 & U7351); 
assign U7353 = ~(SUB_450_U6 & U2354); 
assign U7354 = ~(R2238_U19 & U7351); 
assign U7355 = ~(SUB_450_U19 & U2354); 
assign U7364 = ~(R2238_U19 & U4180); 
assign U7475 = ~(U7079 & U4182); 
assign U7695 = ~(U7694 & U7693); 
assign R2027_U78 = ~(R2027_U196 & R2027_U195); 
assign R2027_U79 = ~(R2027_U198 & R2027_U197); 
assign R2027_U124 = ~R2027_U27; 
assign R2027_U138 = ~R2027_U108; 
assign R2027_U192 = ~(R2027_U27 & INSTADDRPOINTER_REG_15__SCAN_IN); 
assign R2027_U193 = ~(R2027_U108 & INSTADDRPOINTER_REG_14__SCAN_IN); 
assign R2358_U76 = ~(R2358_U441 & R2358_U440); 
assign R2358_U77 = ~(R2358_U454 & R2358_U453); 
assign R2358_U450 = ~(R2358_U449 & R2358_U448); 
assign R2358_U490 = ~(R2358_U489 & R2358_U488); 
assign R2358_U511 = ~(U2352 & R2358_U182); 
assign R2358_U513 = ~(U2352 & R2358_U182); 
assign R2358_U518 = ~(R2358_U517 & R2358_U516); 
assign R2358_U522 = ~(U2352 & R2358_U184); 
assign R2358_U529 = ~(U2352 & R2358_U184); 
assign R2337_U74 = ~(R2337_U181 & R2337_U180); 
assign R2337_U75 = ~(R2337_U183 & R2337_U182); 
assign R2337_U119 = ~R2337_U101; 
assign R2337_U120 = ~R2337_U29; 
assign R2337_U176 = ~(R2337_U29 & PHYADDRPOINTER_REG_18__SCAN_IN); 
assign R2337_U178 = ~(R2337_U101 & PHYADDRPOINTER_REG_17__SCAN_IN); 
assign R2144_U202 = ~(U2355 & R2144_U76); 
assign R2144_U205 = ~(U2355 & R2144_U77); 
assign R2144_U220 = ~(U2355 & R2144_U85); 
assign R2144_U223 = ~(U2355 & R2144_U86); 
assign R2144_U226 = ~(U2355 & R2144_U87); 
assign R2144_U229 = ~(U2355 & R2144_U88); 
assign R2144_U232 = ~(U2355 & R2144_U89); 
assign R2144_U235 = ~(U2355 & R2144_U90); 
assign R2099_U26 = ~(R2099_U210 & R2099_U209); 
assign R2099_U27 = ~(R2099_U183 & R2099_U182); 
assign R2099_U28 = ~(R2099_U204 & R2099_U203); 
assign R2099_U29 = ~(R2099_U207 & R2099_U206); 
assign R2099_U30 = ~(R2099_U198 & R2099_U197); 
assign R2099_U31 = ~(R2099_U201 & R2099_U200); 
assign R2099_U32 = ~(R2099_U186 & R2099_U185); 
assign R2099_U33 = ~(R2099_U189 & R2099_U188); 
assign R2099_U34 = ~(R2099_U195 & R2099_U194); 
assign R2099_U35 = ~(R2099_U192 & R2099_U191); 
assign R2099_U43 = ~(R2099_U284 & R2099_U283); 
assign R2099_U44 = ~(R2099_U287 & R2099_U286); 
assign R2099_U45 = ~(R2099_U227 & R2099_U226); 
assign R2099_U46 = ~(R2099_U230 & R2099_U229); 
assign R2099_U47 = ~(R2099_U233 & R2099_U232); 
assign R2099_U48 = ~(R2099_U236 & R2099_U235); 
assign R2099_U49 = ~(R2099_U239 & R2099_U238); 
assign R2099_U50 = ~(R2099_U242 & R2099_U241); 
assign R2099_U51 = ~(R2099_U245 & R2099_U244); 
assign R2099_U52 = ~(R2099_U248 & R2099_U247); 
assign R2099_U53 = ~(R2099_U251 & R2099_U250); 
assign R2099_U54 = ~(R2099_U254 & R2099_U253); 
assign R2099_U55 = ~(R2099_U257 & R2099_U256); 
assign R2099_U56 = ~(R2099_U278 & R2099_U277); 
assign R2099_U57 = ~(R2099_U281 & R2099_U280); 
assign R2099_U58 = ~(R2099_U272 & R2099_U271); 
assign R2099_U59 = ~(R2099_U275 & R2099_U274); 
assign R2099_U60 = ~(R2099_U266 & R2099_U265); 
assign R2099_U61 = ~(R2099_U269 & R2099_U268); 
assign R2099_U62 = ~(R2099_U260 & R2099_U259); 
assign R2099_U63 = ~(R2099_U263 & R2099_U262); 
assign R2099_U97 = ~(R2099_U290 & R2099_U289); 
assign R2167_U8 = ~U2720; 
assign R2167_U9 = ~U2719; 
assign R2167_U10 = ~U2713; 
assign R2167_U11 = ~U2712; 
assign R2167_U22 = ~U2721; 
assign R2167_U24 = ~(U2715 & R2167_U23); 
assign R2167_U26 = U2721 | U2722; 
assign R2167_U29 = ~(U2720 & R2167_U7); 
assign R2096_U63 = ~(R2096_U126 & R2096_U125); 
assign R2096_U100 = ~R2096_U19; 
assign R2096_U123 = ~(R2096_U19 & REIP_REG_9__SCAN_IN); 
assign ADD_371_U28 = ~ADD_371_U9; 
assign ADD_371_U39 = ~(U3218 & ADD_371_U9); 
assign ADD_371_U42 = ~(ADD_371_U27 & ADD_371_U8); 
assign ADD_405_U64 = ~(ADD_405_U130 & ADD_405_U129); 
assign ADD_405_U103 = ~ADD_405_U19; 
assign ADD_405_U127 = ~(ADD_405_U19 & INSTADDRPOINTER_REG_9__SCAN_IN); 
assign GTE_485_U7 = ~(R2238_U19 | R2238_U20 | R2238_U22 | R2238_U21); 
assign ADD_515_U63 = ~(ADD_515_U126 & ADD_515_U125); 
assign ADD_515_U100 = ~ADD_515_U19; 
assign ADD_515_U123 = ~(ADD_515_U19 & INSTADDRPOINTER_REG_9__SCAN_IN); 
assign U2711 = ~(U7365 & U7364); 
assign U2716 = ~(U7353 & U7352); 
assign U2717 = ~(U7355 & U7354); 
assign U2723 = U7224 & U7071; 
assign U2724 = U7241 & U7071; 
assign U2725 = U7258 & U7071; 
assign U2726 = U7608 & U7071; 
assign U2727 = U7290 & U7071; 
assign U2728 = U7307 & U7071; 
assign U2729 = U7324 & U7071; 
assign U2730 = U7341 & U7071; 
assign U2732 = U7071 & U7070; 
assign U2733 = U7102 & U7071; 
assign U2734 = U7119 & U7071; 
assign U2735 = U7606 & U7071; 
assign U2736 = U7151 & U7071; 
assign U2737 = U7168 & U7071; 
assign U2738 = U7185 & U7071; 
assign U2739 = U7202 & U7071; 
assign U2761 = ~(U6916 & U6915); 
assign U2762 = ~(U6918 & U6917); 
assign U2763 = ~(U6920 & U6919); 
assign U2764 = ~(U6922 & U6921); 
assign U3437 = ~(U4062 & U7081 & U4063 & U4065); 
assign U4102 = U7078 & U3421 & U4099 & U4101; 
assign U4104 = U7493 & U7477 & U7476 & U7475; 
assign U4144 = U4143 & U7347; 
assign U5487 = ~(U4482 & U7695); 
assign U6828 = ~(R2337_U74 & U2352); 
assign U6831 = ~(R2337_U75 & U2352); 
assign U7467 = ~(U4105 & U7081 & U4106 & U4108); 
assign U7780 = ~(U7695 & U4482); 
assign R2027_U31 = ~(R2027_U88 & R2027_U124); 
assign R2027_U107 = ~(R2027_U124 & INSTADDRPOINTER_REG_15__SCAN_IN); 
assign R2027_U191 = ~(R2027_U124 & R2027_U26); 
assign R2027_U194 = ~(R2027_U138 & R2027_U23); 
assign R2358_U183 = ~U2617; 
assign R2358_U185 = ~U2616; 
assign R2358_U442 = ~R2358_U76; 
assign R2358_U455 = ~R2358_U77; 
assign R2358_U515 = ~(R2358_U514 & R2358_U513); 
assign R2358_U520 = ~(U2617 & R2358_U22); 
assign R2358_U525 = ~(U2616 & R2358_U22); 
assign R2358_U531 = ~(R2358_U530 & R2358_U529); 
assign R2337_U32 = ~(R2337_U87 & R2337_U120); 
assign R2337_U100 = ~(R2337_U120 & PHYADDRPOINTER_REG_18__SCAN_IN); 
assign R2337_U177 = ~(R2337_U120 & R2337_U31); 
assign R2337_U179 = ~(R2337_U119 & R2337_U27); 
assign R2144_U14 = ~U2751; 
assign R2144_U27 = ~(R2144_U206 & R2144_U205); 
assign R2144_U29 = ~(R2144_U203 & R2144_U202); 
assign R2144_U31 = ~(R2144_U224 & R2144_U223); 
assign R2144_U32 = ~(R2144_U221 & R2144_U220); 
assign R2144_U33 = ~(R2144_U227 & R2144_U226); 
assign R2144_U34 = ~(R2144_U230 & R2144_U229); 
assign R2144_U35 = ~(R2144_U233 & R2144_U232); 
assign R2144_U36 = ~(R2144_U236 & R2144_U235); 
assign R2099_U88 = R2099_U34 & R2099_U35; 
assign R2099_U89 = R2099_U31 & R2099_U30; 
assign R2099_U90 = R2099_U29 & R2099_U28; 
assign R2099_U91 = R2099_U26 & R2099_U27; 
assign R2099_U92 = R2099_U63 & R2099_U62; 
assign R2099_U93 = R2099_U61 & R2099_U60; 
assign R2099_U94 = R2099_U59 & R2099_U58; 
assign R2099_U95 = R2099_U57 & R2099_U56; 
assign R2099_U96 = R2099_U44 & R2099_U43; 
assign R2099_U147 = ~(R2099_U32 & R2099_U146); 
assign R2099_U152 = ~(U2678 & R2099_U33); 
assign R2099_U184 = ~R2099_U27; 
assign R2099_U187 = ~R2099_U32; 
assign R2099_U190 = ~R2099_U33; 
assign R2099_U193 = ~R2099_U35; 
assign R2099_U196 = ~R2099_U34; 
assign R2099_U199 = ~R2099_U30; 
assign R2099_U202 = ~R2099_U31; 
assign R2099_U205 = ~R2099_U28; 
assign R2099_U208 = ~R2099_U29; 
assign R2099_U211 = ~R2099_U26; 
assign R2099_U228 = ~R2099_U45; 
assign R2099_U231 = ~R2099_U46; 
assign R2099_U234 = ~R2099_U47; 
assign R2099_U237 = ~R2099_U48; 
assign R2099_U240 = ~R2099_U49; 
assign R2099_U243 = ~R2099_U50; 
assign R2099_U246 = ~R2099_U51; 
assign R2099_U249 = ~R2099_U52; 
assign R2099_U252 = ~R2099_U53; 
assign R2099_U255 = ~R2099_U54; 
assign R2099_U258 = ~R2099_U55; 
assign R2099_U261 = ~R2099_U62; 
assign R2099_U264 = ~R2099_U63; 
assign R2099_U267 = ~R2099_U60; 
assign R2099_U270 = ~R2099_U61; 
assign R2099_U273 = ~R2099_U58; 
assign R2099_U276 = ~R2099_U59; 
assign R2099_U279 = ~R2099_U56; 
assign R2099_U282 = ~R2099_U57; 
assign R2099_U285 = ~R2099_U43; 
assign R2099_U288 = ~R2099_U44; 
assign R2099_U291 = ~R2099_U97; 
assign R2099_U319 = ~(R2099_U33 & R2099_U6); 
assign R2099_U321 = ~(R2099_U33 & R2099_U6); 
assign R2099_U348 = ~(R2099_U32 & R2099_U347); 
assign R2167_U12 = ~U2718; 
assign R2167_U15 = ~U2356; 
assign R2167_U25 = ~(U2715 & R2167_U22); 
assign R2167_U27 = ~(U2714 & R2167_U8); 
assign R2167_U30 = ~(U2719 & R2167_U10); 
assign R2167_U32 = ~(U2713 & R2167_U9); 
assign R2167_U35 = ~(U2718 & R2167_U11); 
assign R2096_U20 = ~(R2096_U100 & REIP_REG_9__SCAN_IN); 
assign R2096_U124 = ~(R2096_U100 & R2096_U18); 
assign ADD_371_U11 = ~(U3218 & ADD_371_U28); 
assign ADD_371_U25 = ADD_371_U42 & ADD_371_U41; 
assign ADD_371_U40 = ~(ADD_371_U28 & ADD_371_U10); 
assign ADD_405_U20 = ~(ADD_405_U103 & INSTADDRPOINTER_REG_9__SCAN_IN); 
assign ADD_405_U128 = ~(ADD_405_U103 & ADD_405_U18); 
assign GTE_485_U6 = ~(R2238_U6 | GTE_485_U7); 
assign ADD_515_U20 = ~(ADD_515_U100 & INSTADDRPOINTER_REG_9__SCAN_IN); 
assign ADD_515_U124 = ~(ADD_515_U100 & ADD_515_U18); 
assign U2519 = U3732 & U5487; 
assign U2618 = ~(U6829 & U6830 & U6831); 
assign U2744 = U7467 & U7466; 
assign U3233 = ~(U7780 & U7779 & U4146 & U4144); 
assign U3375 = ~GTE_485_U6; 
assign U4013 = U6826 & U6827 & U6828; 
assign U5458 = ~(U4203 & U3244 & GTE_485_U6); 
assign U6137 = ~(U4182 & U2447 & GTE_485_U6); 
assign U6348 = ~(U4192 & GTE_485_U6); 
assign U6796 = ~(U2724 & U6734); 
assign U6800 = ~(U2725 & U6734); 
assign U6804 = ~(U2726 & U6734); 
assign U6813 = ~(U2727 & U6734); 
assign U6817 = ~(U2728 & U6734); 
assign U6821 = ~(U2729 & U6734); 
assign U6825 = ~(U2730 & U6734); 
assign U6870 = ~(ADD_371_U25 & U4196); 
assign U7082 = ~U3437; 
assign U7084 = ~(U3437 & INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign U7494 = ~(U4104 & U4103 & U4102); 
assign R2027_U76 = ~(R2027_U192 & R2027_U191); 
assign R2027_U77 = ~(R2027_U194 & R2027_U193); 
assign R2027_U117 = ~R2027_U31; 
assign R2027_U137 = ~R2027_U107; 
assign R2027_U188 = ~(R2027_U31 & INSTADDRPOINTER_REG_17__SCAN_IN); 
assign R2027_U189 = ~(R2027_U107 & INSTADDRPOINTER_REG_16__SCAN_IN); 
assign R2358_U519 = ~(U2352 & R2358_U183); 
assign R2358_U524 = ~(U2352 & R2358_U185); 
assign R2337_U72 = ~(R2337_U177 & R2337_U176); 
assign R2337_U73 = ~(R2337_U179 & R2337_U178); 
assign R2337_U121 = ~R2337_U100; 
assign R2337_U122 = ~R2337_U32; 
assign R2337_U172 = ~(R2337_U32 & PHYADDRPOINTER_REG_20__SCAN_IN); 
assign R2337_U174 = ~(R2337_U100 & PHYADDRPOINTER_REG_19__SCAN_IN); 
assign R2182_U14 = ~U2737; 
assign R2182_U15 = ~U2738; 
assign R2182_U16 = ~(U2723 & U2739); 
assign R2182_U17 = ~U2736; 
assign R2182_U18 = ~U2735; 
assign R2182_U20 = ~U2734; 
assign R2182_U23 = ~U2733; 
assign R2182_U36 = U2738 & U2737; 
assign R2182_U37 = U2735 & U2736; 
assign R2182_U39 = ~U2732; 
assign R2182_U60 = U2739 | U2723; 
assign R2144_U6 = R2144_U36 & R2144_U35 & R2144_U27 & R2144_U29; 
assign R2144_U64 = R2144_U34 & R2144_U33 & R2144_U31 & R2144_U32; 
assign R2144_U65 = R2144_U34 & R2144_U33; 
assign R2144_U66 = R2144_U36 & R2144_U27 & R2144_U29; 
assign R2144_U67 = R2144_U29 & R2144_U27; 
assign R2144_U68 = ~U2762; 
assign R2144_U69 = ~U2761; 
assign R2144_U70 = ~U2763; 
assign R2144_U71 = ~U2764; 
assign R2144_U165 = ~(U2762 & R2144_U12); 
assign R2144_U167 = ~(U2761 & R2144_U12); 
assign R2144_U169 = ~(U2763 & R2144_U12); 
assign R2144_U172 = ~(U2762 & R2144_U12); 
assign R2144_U175 = ~(U2763 & R2144_U12); 
assign R2144_U177 = ~(U2764 & R2144_U12); 
assign R2144_U180 = ~(U2761 & R2144_U12); 
assign R2144_U201 = ~(U2764 & R2144_U12); 
assign R2144_U204 = ~R2144_U29; 
assign R2144_U207 = ~R2144_U27; 
assign R2144_U222 = ~R2144_U32; 
assign R2144_U225 = ~R2144_U31; 
assign R2144_U228 = ~R2144_U33; 
assign R2144_U231 = ~R2144_U34; 
assign R2144_U234 = ~R2144_U35; 
assign R2144_U237 = ~R2144_U36; 
assign R2099_U140 = ~(R2099_U148 & R2099_U147); 
assign R2099_U150 = ~(R2099_U190 & R2099_U6); 
assign R2099_U318 = ~(R2099_U190 & U2678); 
assign R2099_U320 = ~(R2099_U190 & U2678); 
assign R2099_U349 = ~(R2099_U98 & R2099_U187); 
assign R2167_U6 = ~U2716; 
assign R2167_U13 = ~U2717; 
assign R2167_U14 = ~U2711; 
assign R2167_U18 = R2167_U29 & R2167_U30; 
assign R2167_U28 = ~(R2167_U27 & R2167_U26 & R2167_U25 & R2167_U24); 
assign R2167_U33 = ~(U2712 & R2167_U12); 
assign R2167_U41 = ~(U2716 & R2167_U15); 
assign R2167_U43 = ~(U2716 & R2167_U16); 
assign R2096_U62 = ~(R2096_U124 & R2096_U123); 
assign R2096_U101 = ~R2096_U20; 
assign R2096_U181 = ~(R2096_U20 & REIP_REG_10__SCAN_IN); 
assign ADD_371_U20 = ~(ADD_371_U40 & ADD_371_U39); 
assign ADD_371_U29 = ~ADD_371_U11; 
assign ADD_371_U37 = ~(U3219 & ADD_371_U11); 
assign ADD_405_U63 = ~(ADD_405_U128 & ADD_405_U127); 
assign ADD_405_U104 = ~ADD_405_U20; 
assign ADD_405_U185 = ~(ADD_405_U20 & INSTADDRPOINTER_REG_10__SCAN_IN); 
assign ADD_515_U62 = ~(ADD_515_U124 & ADD_515_U123); 
assign ADD_515_U101 = ~ADD_515_U20; 
assign ADD_515_U181 = ~(ADD_515_U20 & INSTADDRPOINTER_REG_10__SCAN_IN); 
assign U2666 = ~(U6825 & U4013); 
assign U2741 = ~(U4066 & U7084); 
assign U2743 = U7494 & U7458; 
assign U3725 = U3724 & U5458; 
assign U4486 = ~(U4465 & U3375); 
assign U4495 = ~(U4203 & U3375); 
assign U5557 = ~(U3746 & U2519); 
assign U6820 = ~(R2337_U72 & U2352); 
assign U6824 = ~(R2337_U73 & U2352); 
assign U6868 = ~(ADD_371_U20 & U4196); 
assign U7480 = ~(U4097 & U7082); 
assign U7497 = ~(U3734 & U2519); 
assign U7728 = ~(U4465 & U3375); 
assign R2027_U34 = ~(R2027_U89 & R2027_U117); 
assign R2027_U106 = ~(R2027_U117 & INSTADDRPOINTER_REG_17__SCAN_IN); 
assign R2027_U187 = ~(R2027_U117 & R2027_U30); 
assign R2027_U190 = ~(R2027_U137 & R2027_U28); 
assign R2358_U79 = ~(R2358_U520 & R2358_U519); 
assign R2358_U80 = ~(R2358_U525 & R2358_U524); 
assign R2358_U186 = ~U2618; 
assign R2358_U528 = ~(U2618 & R2358_U22); 
assign R2358_U533 = ~(U2618 & R2358_U22); 
assign R2337_U35 = ~(R2337_U88 & R2337_U122); 
assign R2337_U99 = ~(R2337_U122 & PHYADDRPOINTER_REG_20__SCAN_IN); 
assign R2337_U173 = ~(R2337_U122 & R2337_U34); 
assign R2337_U175 = ~(R2337_U121 & R2337_U30); 
assign R2182_U6 = R2182_U60 & R2182_U16; 
assign R2182_U7 = ~U2744; 
assign R2182_U8 = ~U3233; 
assign R2182_U9 = ~(U3233 & U2744); 
assign R2182_U49 = ~R2182_U16; 
assign R2182_U82 = ~(U2738 & R2182_U16); 
assign R2144_U63 = R2144_U6 & R2144_U64; 
assign R2144_U164 = ~(U2355 & R2144_U68); 
assign R2144_U166 = ~(U2355 & R2144_U69); 
assign R2144_U168 = ~(U2355 & R2144_U70); 
assign R2144_U171 = ~(U2355 & R2144_U68); 
assign R2144_U174 = ~(U2355 & R2144_U70); 
assign R2144_U176 = ~(U2355 & R2144_U71); 
assign R2144_U179 = ~(U2355 & R2144_U69); 
assign R2144_U200 = ~(U2355 & R2144_U71); 
assign R2099_U86 = ~(R2099_U349 & R2099_U348); 
assign R2099_U139 = R2099_U319 & R2099_U318; 
assign R2099_U149 = ~R2099_U140; 
assign R2099_U151 = ~(R2099_U150 & R2099_U140); 
assign R2099_U322 = ~(R2099_U321 & R2099_U320); 
assign R2167_U19 = R2167_U32 & R2167_U33; 
assign R2167_U31 = ~(R2167_U18 & R2167_U28); 
assign R2167_U36 = ~(U2717 & R2167_U14); 
assign R2167_U38 = ~(U2711 & R2167_U13); 
assign R2167_U39 = ~(U2356 & R2167_U6); 
assign R2167_U46 = ~(R2167_U6 & STATE2_REG_0__SCAN_IN); 
assign R2096_U22 = ~(R2096_U101 & REIP_REG_10__SCAN_IN); 
assign R2096_U182 = ~(R2096_U101 & R2096_U21); 
assign ADD_371_U13 = ~(U3219 & ADD_371_U29); 
assign ADD_371_U38 = ~(ADD_371_U29 & ADD_371_U12); 
assign ADD_405_U22 = ~(ADD_405_U104 & INSTADDRPOINTER_REG_10__SCAN_IN); 
assign ADD_405_U186 = ~(ADD_405_U104 & ADD_405_U21); 
assign ADD_515_U22 = ~(ADD_515_U101 & INSTADDRPOINTER_REG_10__SCAN_IN); 
assign ADD_515_U182 = ~(ADD_515_U101 & ADD_515_U21); 
assign U2742 = U7480 & U7479; 
assign U3424 = ~(U2447 & U4486); 
assign U3726 = U3725 & U2518; 
assign U4011 = U6818 & U6819 & U6820; 
assign U4012 = U6822 & U6823 & U6824; 
assign U6792 = ~(R2182_U6 & U6734); 
assign R2027_U74 = ~(R2027_U188 & R2027_U187); 
assign R2027_U75 = ~(R2027_U190 & R2027_U189); 
assign R2027_U114 = ~R2027_U34; 
assign R2027_U136 = ~R2027_U106; 
assign R2027_U184 = ~(R2027_U34 & INSTADDRPOINTER_REG_19__SCAN_IN); 
assign R2027_U185 = ~(R2027_U106 & INSTADDRPOINTER_REG_18__SCAN_IN); 
assign R2358_U189 = ~U2666; 
assign R2358_U521 = ~R2358_U79; 
assign R2358_U526 = ~R2358_U80; 
assign R2358_U527 = ~(U2352 & R2358_U186); 
assign R2358_U532 = ~(U2352 & R2358_U186); 
assign R2358_U540 = ~(U2666 & R2358_U22); 
assign R2358_U600 = ~(U2666 & R2358_U22); 
assign R2337_U70 = ~(R2337_U173 & R2337_U172); 
assign R2337_U71 = ~(R2337_U175 & R2337_U174); 
assign R2337_U123 = ~R2337_U99; 
assign R2337_U124 = ~R2337_U35; 
assign R2337_U168 = ~(R2337_U35 & PHYADDRPOINTER_REG_22__SCAN_IN); 
assign R2337_U170 = ~(R2337_U99 & PHYADDRPOINTER_REG_21__SCAN_IN); 
assign R2182_U11 = ~U2741; 
assign R2182_U19 = ~(R2182_U36 & R2182_U49); 
assign R2182_U44 = ~(R2182_U49 & U2738); 
assign R2182_U50 = ~R2182_U9; 
assign R2182_U51 = U2743 | U2731; 
assign R2182_U52 = ~(U2731 & U2743); 
assign R2182_U62 = ~(U2731 & U2743); 
assign R2182_U81 = ~(R2182_U49 & R2182_U15); 
assign R2182_U85 = ~(U3233 & R2182_U7); 
assign R2182_U86 = ~(U2744 & R2182_U8); 
assign R2144_U81 = ~(R2144_U165 & R2144_U164 & R2144_U22); 
assign R2144_U104 = ~(R2144_U167 & R2144_U166 & R2144_U17); 
assign R2144_U105 = ~(R2144_U175 & R2144_U174 & R2144_U20); 
assign R2144_U106 = ~(R2144_U201 & R2144_U200 & R2144_U18); 
assign R2144_U170 = ~(R2144_U169 & R2144_U168); 
assign R2144_U173 = ~(R2144_U172 & R2144_U171); 
assign R2144_U178 = ~(R2144_U177 & R2144_U176); 
assign R2144_U181 = ~(R2144_U180 & R2144_U179); 
assign R2099_U137 = ~(R2099_U152 & R2099_U151); 
assign R2099_U323 = ~(R2099_U139 & R2099_U140); 
assign R2099_U324 = ~(R2099_U149 & R2099_U322); 
assign R2167_U20 = R2167_U35 & R2167_U36; 
assign R2167_U21 = R2167_U38 & R2167_U39; 
assign R2167_U34 = ~(R2167_U19 & R2167_U31); 
assign R2096_U91 = ~(R2096_U182 & R2096_U181); 
assign R2096_U102 = ~R2096_U22; 
assign R2096_U179 = ~(R2096_U22 & REIP_REG_11__SCAN_IN); 
assign ADD_371_U19 = ~(ADD_371_U38 & ADD_371_U37); 
assign ADD_371_U30 = ~ADD_371_U13; 
assign ADD_371_U35 = ~(U3220 & ADD_371_U13); 
assign ADD_405_U91 = ~(ADD_405_U186 & ADD_405_U185); 
assign ADD_405_U105 = ~ADD_405_U22; 
assign ADD_405_U183 = ~(ADD_405_U22 & INSTADDRPOINTER_REG_11__SCAN_IN); 
assign ADD_515_U91 = ~(ADD_515_U182 & ADD_515_U181); 
assign ADD_515_U102 = ~ADD_515_U22; 
assign ADD_515_U179 = ~(ADD_515_U22 & INSTADDRPOINTER_REG_11__SCAN_IN); 
assign U2664 = ~(U6817 & U4011); 
assign U2665 = ~(U6821 & U4012); 
assign U4487 = ~U3424; 
assign U6807 = ~(R2337_U70 & U2352); 
assign U6816 = ~(R2337_U71 & U2352); 
assign U6866 = ~(ADD_371_U19 & U4196); 
assign U7667 = ~(U4482 & U3424); 
assign R2027_U36 = ~(R2027_U90 & R2027_U114); 
assign R2027_U105 = ~(R2027_U114 & INSTADDRPOINTER_REG_19__SCAN_IN); 
assign R2027_U183 = ~(R2027_U114 & R2027_U33); 
assign R2027_U186 = ~(R2027_U136 & R2027_U29); 
assign R2358_U13 = R2358_U528 & R2358_U527; 
assign R2358_U81 = ~(R2358_U533 & R2358_U532); 
assign R2358_U539 = ~(U2352 & R2358_U189); 
assign R2358_U599 = ~(U2352 & R2358_U189); 
assign R2337_U38 = ~(R2337_U89 & R2337_U124); 
assign R2337_U98 = ~(R2337_U124 & PHYADDRPOINTER_REG_22__SCAN_IN); 
assign R2337_U169 = ~(R2337_U124 & R2337_U37); 
assign R2337_U171 = ~(R2337_U123 & R2337_U33); 
assign R2182_U10 = ~U2742; 
assign R2182_U32 = ~(R2182_U82 & R2182_U81); 
assign R2182_U34 = ~(R2182_U86 & R2182_U85); 
assign R2182_U35 = U2742 & U2741; 
assign R2182_U45 = ~(R2182_U51 & R2182_U62); 
assign R2182_U46 = ~R2182_U19; 
assign R2182_U53 = ~(R2182_U50 & R2182_U51); 
assign R2182_U59 = ~R2182_U44; 
assign R2182_U78 = ~(U2736 & R2182_U19); 
assign R2182_U79 = ~(U2737 & R2182_U44); 
assign R2144_U7 = R2144_U104 & R2144_U81; 
assign R2144_U19 = ~(U2748 & R2144_U178); 
assign R2144_U21 = ~(U2747 & R2144_U170); 
assign R2144_U23 = ~(U2746 & R2144_U173); 
assign R2144_U52 = R2144_U106 & R2144_U105; 
assign R2144_U102 = ~R2144_U81; 
assign R2144_U103 = ~(U2745 & R2144_U181); 
assign R2099_U7 = ~(R2099_U88 & R2099_U137); 
assign R2099_U87 = ~(R2099_U324 & R2099_U323); 
assign R2099_U112 = ~(R2099_U35 & R2099_U137); 
assign R2099_U153 = ~R2099_U137; 
assign R2099_U297 = ~(R2099_U35 & R2099_U137); 
assign R2167_U37 = ~(R2167_U20 & R2167_U34); 
assign R2096_U24 = ~(R2096_U102 & REIP_REG_11__SCAN_IN); 
assign R2096_U180 = ~(R2096_U102 & R2096_U23); 
assign ADD_371_U6 = ADD_371_U22 & ADD_371_U30; 
assign ADD_371_U23 = ~(U3220 & ADD_371_U30); 
assign ADD_371_U36 = ~(ADD_371_U30 & ADD_371_U15); 
assign ADD_405_U24 = ~(ADD_405_U105 & INSTADDRPOINTER_REG_11__SCAN_IN); 
assign ADD_405_U184 = ~(ADD_405_U105 & ADD_405_U23); 
assign ADD_515_U24 = ~(ADD_515_U102 & INSTADDRPOINTER_REG_11__SCAN_IN); 
assign ADD_515_U180 = ~(ADD_515_U102 & ADD_515_U23); 
assign U3305 = ~R2182_U34; 
assign U4008 = U6805 & U6806 & U6807; 
assign U4010 = U6814 & U6815 & U6816; 
assign U5518 = ~(R2182_U34 & U7497); 
assign U5543 = ~(R2182_U34 & U5526); 
assign U6788 = ~(R2182_U32 & U6734); 
assign U6852 = ~(R2182_U34 & U6734); 
assign U6860 = ~(ADD_371_U6 & U4196); 
assign U7034 = ~(R2182_U34 & U3281); 
assign R2027_U72 = ~(R2027_U184 & R2027_U183); 
assign R2027_U73 = ~(R2027_U186 & R2027_U185); 
assign R2027_U121 = ~R2027_U36; 
assign R2027_U135 = ~R2027_U105; 
assign R2027_U178 = ~(R2027_U36 & INSTADDRPOINTER_REG_21__SCAN_IN); 
assign R2027_U179 = ~(R2027_U105 & INSTADDRPOINTER_REG_20__SCAN_IN); 
assign R2358_U187 = ~U2664; 
assign R2358_U188 = ~U2665; 
assign R2358_U534 = ~R2358_U81; 
assign R2358_U536 = ~(U2664 & R2358_U22); 
assign R2358_U538 = ~(U2665 & R2358_U22); 
assign R2358_U601 = ~(R2358_U600 & R2358_U599); 
assign R2358_U603 = ~(U2664 & R2358_U22); 
assign R2358_U606 = ~(U2665 & R2358_U22); 
assign R2337_U68 = ~(R2337_U169 & R2337_U168); 
assign R2337_U69 = ~(R2337_U171 & R2337_U170); 
assign R2337_U125 = ~R2337_U98; 
assign R2337_U126 = ~R2337_U38; 
assign R2337_U164 = ~(R2337_U38 & PHYADDRPOINTER_REG_24__SCAN_IN); 
assign R2337_U166 = ~(R2337_U98 & PHYADDRPOINTER_REG_23__SCAN_IN); 
assign R2182_U21 = ~(R2182_U37 & R2182_U46); 
assign R2182_U41 = ~(R2182_U52 & R2182_U53); 
assign R2182_U43 = ~(R2182_U46 & U2736); 
assign R2182_U61 = ~R2182_U45; 
assign R2182_U77 = ~(R2182_U46 & R2182_U17); 
assign R2182_U80 = ~(R2182_U59 & R2182_U14); 
assign R2182_U83 = ~(R2182_U50 & R2182_U45); 
assign R2144_U5 = R2144_U104 & R2144_U103; 
assign R2144_U44 = R2144_U21 & R2144_U105; 
assign R2144_U46 = R2144_U19 & R2144_U106; 
assign R2144_U53 = R2144_U7 & R2144_U52; 
assign R2144_U61 = R2144_U23 & R2144_U81; 
assign R2144_U107 = ~R2144_U21; 
assign R2144_U108 = ~R2144_U23; 
assign R2144_U120 = ~R2144_U19; 
assign R2144_U126 = ~(R2144_U23 & R2144_U81); 
assign R2144_U149 = ~(R2144_U21 & R2144_U105); 
assign R2144_U150 = ~(R2144_U19 & R2144_U106); 
assign R2144_U156 = ~(R2144_U104 & R2144_U103); 
assign R2099_U154 = ~R2099_U112; 
assign R2099_U155 = ~R2099_U7; 
assign R2099_U223 = ~(R2099_U30 & R2099_U7); 
assign R2099_U225 = ~(R2099_U34 & R2099_U112); 
assign R2099_U296 = ~(R2099_U153 & R2099_U193); 
assign R2167_U40 = ~(R2167_U21 & R2167_U37); 
assign R2096_U90 = ~(R2096_U180 & R2096_U179); 
assign R2096_U103 = ~R2096_U24; 
assign R2096_U177 = ~(R2096_U24 & REIP_REG_12__SCAN_IN); 
assign ADD_371_U18 = ~(ADD_371_U36 & ADD_371_U35); 
assign ADD_371_U31 = ~ADD_371_U23; 
assign ADD_371_U33 = ~(U3221 & ADD_371_U23); 
assign ADD_405_U90 = ~(ADD_405_U184 & ADD_405_U183); 
assign ADD_405_U106 = ~ADD_405_U24; 
assign ADD_405_U181 = ~(ADD_405_U24 & INSTADDRPOINTER_REG_12__SCAN_IN); 
assign ADD_515_U90 = ~(ADD_515_U180 & ADD_515_U179); 
assign ADD_515_U103 = ~ADD_515_U24; 
assign ADD_515_U177 = ~(ADD_515_U24 & INSTADDRPOINTER_REG_12__SCAN_IN); 
assign U2662 = ~(U6804 & U4008); 
assign U2663 = ~(U6813 & U4010); 
assign U2672 = ~(U6854 & U6852 & U6853 & U6856 & U6855); 
assign U2768 = ~(U7034 & U7032 & U7033); 
assign U5519 = ~(U4163 & U5518); 
assign U6799 = ~(R2337_U68 & U2352); 
assign U6803 = ~(R2337_U69 & U2352); 
assign U6864 = ~(ADD_371_U18 & U4196); 
assign R2027_U40 = ~(R2027_U91 & R2027_U121); 
assign R2027_U104 = ~(R2027_U121 & INSTADDRPOINTER_REG_21__SCAN_IN); 
assign R2027_U177 = ~(R2027_U121 & R2027_U35); 
assign R2027_U180 = ~(R2027_U135 & R2027_U32); 
assign R2358_U535 = ~(U2352 & R2358_U187); 
assign R2358_U537 = ~(U2352 & R2358_U188); 
assign R2358_U602 = ~(U2352 & R2358_U187); 
assign R2358_U605 = ~(U2352 & R2358_U188); 
assign R2337_U41 = ~(R2337_U90 & R2337_U126); 
assign R2337_U97 = ~(R2337_U126 & PHYADDRPOINTER_REG_24__SCAN_IN); 
assign R2337_U165 = ~(R2337_U126 & R2337_U40); 
assign R2337_U167 = ~(R2337_U125 & R2337_U36); 
assign R2182_U13 = ~(R2182_U35 & R2182_U41); 
assign R2182_U30 = ~(R2182_U78 & R2182_U77); 
assign R2182_U31 = ~(R2182_U80 & R2182_U79); 
assign R2182_U38 = ~(U2742 & R2182_U41); 
assign R2182_U48 = ~R2182_U21; 
assign R2182_U54 = ~R2182_U41; 
assign R2182_U58 = ~R2182_U43; 
assign R2182_U69 = ~(U2742 & R2182_U41); 
assign R2182_U74 = ~(U2734 & R2182_U21); 
assign R2182_U75 = ~(U2735 & R2182_U43); 
assign R2182_U84 = ~(R2182_U61 & R2182_U9); 
assign R2144_U57 = R2144_U156 & R2144_U21; 
assign R2144_U59 = R2144_U5 & R2144_U105; 
assign R2144_U60 = R2144_U126 & R2144_U21; 
assign R2144_U151 = ~(R2144_U120 & R2144_U105 & R2144_U7); 
assign R2144_U152 = ~(R2144_U107 & R2144_U7); 
assign R2144_U153 = ~(R2144_U108 & R2144_U7); 
assign R2144_U213 = ~(R2144_U5 & R2144_U108); 
assign R2144_U214 = ~(R2144_U102 & R2144_U156); 
assign R2099_U8 = ~(R2099_U89 & R2099_U155); 
assign R2099_U111 = ~(R2099_U155 & R2099_U30); 
assign R2099_U138 = R2099_U297 & R2099_U296; 
assign R2099_U222 = ~(R2099_U199 & R2099_U155); 
assign R2099_U224 = ~(R2099_U154 & R2099_U196); 
assign R2167_U42 = ~(R2167_U40 & R2167_U41); 
assign R2096_U26 = ~(R2096_U103 & REIP_REG_12__SCAN_IN); 
assign R2096_U178 = ~(R2096_U103 & R2096_U25); 
assign ADD_371_U34 = ~(ADD_371_U31 & ADD_371_U14); 
assign ADD_405_U26 = ~(ADD_405_U106 & INSTADDRPOINTER_REG_12__SCAN_IN); 
assign ADD_405_U182 = ~(ADD_405_U106 & ADD_405_U25); 
assign ADD_515_U26 = ~(ADD_515_U103 & INSTADDRPOINTER_REG_12__SCAN_IN); 
assign ADD_515_U178 = ~(ADD_515_U103 & ADD_515_U25); 
assign U4006 = U6797 & U6798 & U6799; 
assign U4007 = U6801 & U6802 & U6803; 
assign U5521 = ~(U2427 & U5519); 
assign U6780 = ~(R2182_U30 & U6734); 
assign U6784 = ~(R2182_U31 & U6734); 
assign R2027_U69 = ~(R2027_U178 & R2027_U177); 
assign R2027_U70 = ~(R2027_U180 & R2027_U179); 
assign R2027_U115 = ~R2027_U40; 
assign R2027_U134 = ~R2027_U104; 
assign R2027_U174 = ~(R2027_U40 & INSTADDRPOINTER_REG_23__SCAN_IN); 
assign R2027_U175 = ~(R2027_U104 & INSTADDRPOINTER_REG_22__SCAN_IN); 
assign R2358_U172 = ~U2672; 
assign R2358_U190 = ~U2663; 
assign R2358_U195 = ~U2662; 
assign R2358_U473 = ~(U2672 & R2358_U22); 
assign R2358_U478 = ~(U2672 & R2358_U22); 
assign R2358_U542 = ~(U2663 & R2358_U22); 
assign R2358_U552 = ~(U2662 & R2358_U22); 
assign R2358_U597 = ~(U2663 & R2358_U22); 
assign R2358_U604 = ~(R2358_U603 & R2358_U602); 
assign R2358_U607 = ~(R2358_U606 & R2358_U605); 
assign R2337_U66 = ~(R2337_U165 & R2337_U164); 
assign R2337_U67 = ~(R2337_U167 & R2337_U166); 
assign R2337_U127 = ~R2337_U97; 
assign R2337_U128 = ~R2337_U41; 
assign R2337_U160 = ~(R2337_U41 & PHYADDRPOINTER_REG_26__SCAN_IN); 
assign R2337_U162 = ~(R2337_U97 & PHYADDRPOINTER_REG_25__SCAN_IN); 
assign R2182_U22 = ~(R2182_U48 & U2734); 
assign R2182_U33 = ~(R2182_U84 & R2182_U83); 
assign R2182_U47 = ~R2182_U13; 
assign R2182_U55 = ~R2182_U38; 
assign R2182_U64 = ~(U2740 & R2182_U13); 
assign R2182_U65 = ~(U2741 & R2182_U38); 
assign R2182_U70 = ~(R2182_U54 & R2182_U10); 
assign R2182_U73 = ~(R2182_U48 & R2182_U20); 
assign R2182_U76 = ~(R2182_U58 & R2182_U18); 
assign R2144_U54 = R2144_U103 & R2144_U151 & R2144_U153 & R2144_U152; 
assign R2144_U74 = ~U2768; 
assign R2144_U189 = ~(U2768 & R2144_U12); 
assign R2144_U191 = ~(U2768 & R2144_U12); 
assign R2099_U41 = ~(R2099_U223 & R2099_U222); 
assign R2099_U42 = ~(R2099_U225 & R2099_U224); 
assign R2099_U156 = ~R2099_U111; 
assign R2099_U157 = ~R2099_U8; 
assign R2099_U219 = ~(R2099_U28 & R2099_U8); 
assign R2099_U221 = ~(R2099_U31 & R2099_U111); 
assign R2167_U44 = ~(R2167_U42 & R2167_U6); 
assign R2167_U47 = ~(U2716 & R2167_U42); 
assign R2096_U89 = ~(R2096_U178 & R2096_U177); 
assign R2096_U104 = ~R2096_U26; 
assign R2096_U175 = ~(R2096_U26 & REIP_REG_13__SCAN_IN); 
assign ADD_371_U17 = ~(ADD_371_U34 & ADD_371_U33); 
assign ADD_405_U89 = ~(ADD_405_U182 & ADD_405_U181); 
assign ADD_405_U107 = ~ADD_405_U26; 
assign ADD_405_U179 = ~(ADD_405_U26 & INSTADDRPOINTER_REG_13__SCAN_IN); 
assign ADD_515_U89 = ~(ADD_515_U178 & ADD_515_U177); 
assign ADD_515_U104 = ~ADD_515_U26; 
assign ADD_515_U175 = ~(ADD_515_U26 & INSTADDRPOINTER_REG_13__SCAN_IN); 
assign U2442 = R2182_U33 & R2182_U34; 
assign U2443 = R2182_U33 & U3305; 
assign U2445 = ~(R2182_U33 | R2182_U34); 
assign U2660 = ~(U6796 & U4006); 
assign U2661 = ~(U6800 & U4007); 
assign U3306 = ~R2182_U33; 
assign U5511 = ~(R2182_U33 & U7497); 
assign U5540 = ~(R2182_U33 & U5526); 
assign U6791 = ~(R2337_U66 & U2352); 
assign U6795 = ~(R2337_U67 & U2352); 
assign U6847 = ~(R2182_U33 & U6734); 
assign U6862 = ~(ADD_371_U17 & U4196); 
assign U7031 = ~(R2182_U33 & U3281); 
assign R2027_U43 = ~(R2027_U92 & R2027_U115); 
assign R2027_U103 = ~(R2027_U115 & INSTADDRPOINTER_REG_23__SCAN_IN); 
assign R2027_U173 = ~(R2027_U115 & R2027_U39); 
assign R2027_U176 = ~(R2027_U134 & R2027_U37); 
assign R2358_U472 = ~(U2352 & R2358_U172); 
assign R2358_U477 = ~(U2352 & R2358_U172); 
assign R2358_U541 = ~(U2352 & R2358_U190); 
assign R2358_U551 = ~(U2352 & R2358_U195); 
assign R2358_U596 = ~(U2352 & R2358_U190); 
assign R2337_U43 = ~(R2337_U128 & PHYADDRPOINTER_REG_26__SCAN_IN); 
assign R2337_U161 = ~(R2337_U128 & R2337_U42); 
assign R2337_U163 = ~(R2337_U127 & R2337_U39); 
assign R2182_U5 = R2182_U47 & U2740; 
assign R2182_U28 = ~(R2182_U74 & R2182_U73); 
assign R2182_U29 = ~(R2182_U76 & R2182_U75); 
assign R2182_U42 = R2182_U70 & R2182_U69; 
assign R2182_U56 = ~R2182_U22; 
assign R2182_U63 = ~(R2182_U47 & R2182_U12); 
assign R2182_U66 = ~(R2182_U55 & R2182_U11); 
assign R2182_U71 = ~(U2733 & R2182_U22); 
assign R2144_U188 = ~(U2355 & R2144_U74); 
assign R2144_U190 = ~(U2355 & R2144_U74); 
assign R2099_U9 = ~(R2099_U90 & R2099_U157); 
assign R2099_U110 = ~(R2099_U157 & R2099_U28); 
assign R2099_U218 = ~(R2099_U205 & R2099_U157); 
assign R2099_U220 = ~(R2099_U156 & R2099_U202); 
assign R2167_U45 = ~(R2167_U44 & R2167_U43); 
assign R2167_U48 = ~(R2167_U47 & R2167_U46); 
assign R2096_U28 = ~(R2096_U104 & REIP_REG_13__SCAN_IN); 
assign R2096_U176 = ~(R2096_U104 & R2096_U27); 
assign ADD_405_U28 = ~(ADD_405_U107 & INSTADDRPOINTER_REG_13__SCAN_IN); 
assign ADD_405_U180 = ~(ADD_405_U107 & ADD_405_U27); 
assign ADD_515_U28 = ~(ADD_515_U104 & INSTADDRPOINTER_REG_13__SCAN_IN); 
assign ADD_515_U176 = ~(ADD_515_U104 & ADD_515_U27); 
assign U2444 = R2182_U34 & U3306; 
assign U2671 = ~(U6851 & U6850 & U4015 & U6847); 
assign U2767 = ~(U7031 & U7029 & U7030); 
assign U3304 = ~R2182_U42; 
assign U4004 = U6789 & U6790 & U6791; 
assign U4005 = U6793 & U6794 & U6795; 
assign U5500 = ~(R2182_U42 & U7497); 
assign U5513 = ~(U3738 & U5511); 
assign U5535 = ~(R2182_U42 & U5526); 
assign U6747 = ~(R2182_U5 & U6734); 
assign U6772 = ~(R2182_U28 & U6734); 
assign U6776 = ~(R2182_U29 & U6734); 
assign U6808 = ~(R2182_U42 & U6734); 
assign U6928 = ~(R2182_U42 & U3281); 
assign R2027_U67 = ~(R2027_U174 & R2027_U173); 
assign R2027_U68 = ~(R2027_U176 & R2027_U175); 
assign R2027_U116 = ~R2027_U43; 
assign R2027_U133 = ~R2027_U103; 
assign R2027_U170 = ~(R2027_U43 & INSTADDRPOINTER_REG_25__SCAN_IN); 
assign R2027_U171 = ~(R2027_U103 & INSTADDRPOINTER_REG_24__SCAN_IN); 
assign R2358_U78 = ~(R2358_U552 & R2358_U551); 
assign R2358_U193 = ~U2660; 
assign R2358_U194 = ~U2661; 
assign R2358_U474 = ~(R2358_U473 & R2358_U472); 
assign R2358_U548 = ~(U2660 & R2358_U22); 
assign R2358_U550 = ~(U2661 & R2358_U22); 
assign R2358_U573 = ~(U2660 & R2358_U22); 
assign R2358_U576 = ~(U2661 & R2358_U22); 
assign R2358_U598 = ~(R2358_U597 & R2358_U596); 
assign R2337_U64 = ~(R2337_U161 & R2337_U160); 
assign R2337_U65 = ~(R2337_U163 & R2337_U162); 
assign R2337_U129 = ~R2337_U43; 
assign R2337_U158 = ~(R2337_U43 & PHYADDRPOINTER_REG_27__SCAN_IN); 
assign R2182_U24 = ~(R2182_U64 & R2182_U63); 
assign R2182_U25 = ~(R2182_U66 & R2182_U65); 
assign R2182_U40 = ~(U2733 & R2182_U56); 
assign R2182_U72 = ~(R2182_U56 & R2182_U23); 
assign R2144_U112 = ~(R2144_U189 & R2144_U188 & R2144_U15); 
assign R2144_U192 = ~(R2144_U191 & R2144_U190); 
assign R2099_U39 = ~(R2099_U219 & R2099_U218); 
assign R2099_U40 = ~(R2099_U221 & R2099_U220); 
assign R2099_U158 = ~R2099_U110; 
assign R2099_U159 = ~R2099_U9; 
assign R2099_U215 = ~(R2099_U27 & R2099_U9); 
assign R2099_U217 = ~(R2099_U29 & R2099_U110); 
assign R2167_U49 = ~(R2167_U45 & R2167_U15); 
assign R2167_U50 = ~(U2356 & R2167_U48); 
assign R2096_U88 = ~(R2096_U176 & R2096_U175); 
assign R2096_U105 = ~R2096_U28; 
assign R2096_U173 = ~(R2096_U28 & REIP_REG_14__SCAN_IN); 
assign ADD_405_U88 = ~(ADD_405_U180 & ADD_405_U179); 
assign ADD_405_U108 = ~ADD_405_U28; 
assign ADD_405_U177 = ~(ADD_405_U28 & INSTADDRPOINTER_REG_14__SCAN_IN); 
assign ADD_515_U88 = ~(ADD_515_U176 & ADD_515_U175); 
assign ADD_515_U105 = ~ADD_515_U28; 
assign ADD_515_U173 = ~(ADD_515_U28 & INSTADDRPOINTER_REG_14__SCAN_IN); 
assign U2438 = R2182_U42 & R2182_U25; 
assign U2440 = R2182_U25 & U3304; 
assign U2441 = ~(R2182_U42 | R2182_U25); 
assign U2658 = ~(U6788 & U4004); 
assign U2659 = ~(U6792 & U4005); 
assign U2667 = ~(U6747 & U3994); 
assign U2670 = ~(U6812 & U6811 & U4009 & U6808); 
assign U2766 = ~(U6927 & U6926 & U6928); 
assign U3303 = ~R2182_U25; 
assign U3454 = U2427 & U4203 & R2182_U24; 
assign U3475 = R2182_U24 & U4203; 
assign U5491 = ~(R2182_U25 & U7497); 
assign U5502 = ~(U3737 & U5500); 
assign U5516 = ~(U2427 & U5513); 
assign U5531 = ~(R2182_U25 & U5526); 
assign U6751 = ~(R2182_U24 & U6734); 
assign U6763 = ~(R2182_U25 & U6734); 
assign U6783 = ~(R2337_U64 & U2352); 
assign U6787 = ~(R2337_U65 & U2352); 
assign U6925 = ~(R2182_U25 & U3281); 
assign R2027_U46 = ~(R2027_U93 & R2027_U116); 
assign R2027_U102 = ~(R2027_U116 & INSTADDRPOINTER_REG_25__SCAN_IN); 
assign R2027_U169 = ~(R2027_U116 & R2027_U42); 
assign R2027_U172 = ~(R2027_U133 & R2027_U38); 
assign R2358_U171 = ~U2671; 
assign R2358_U470 = ~(U2671 & R2358_U22); 
assign R2358_U476 = ~(U2671 & R2358_U22); 
assign R2358_U547 = ~(U2352 & R2358_U193); 
assign R2358_U549 = ~(U2352 & R2358_U194); 
assign R2358_U553 = ~R2358_U78; 
assign R2358_U572 = ~(U2352 & R2358_U193); 
assign R2358_U575 = ~(U2352 & R2358_U194); 
assign R2337_U45 = ~(R2337_U129 & PHYADDRPOINTER_REG_27__SCAN_IN); 
assign R2337_U159 = ~(R2337_U129 & R2337_U44); 
assign R2182_U27 = ~(R2182_U72 & R2182_U71); 
assign R2182_U57 = ~R2182_U40; 
assign R2182_U67 = ~(U2732 & R2182_U40); 
assign R2144_U73 = ~U2767; 
assign R2144_U113 = ~(U2752 & R2144_U192); 
assign R2144_U115 = ~(U2355 & R2144_U112); 
assign R2144_U129 = ~(U2355 & R2144_U112); 
assign R2144_U186 = ~(U2767 & R2144_U12); 
assign R2099_U10 = ~(R2099_U91 & R2099_U159); 
assign R2099_U109 = ~(R2099_U159 & R2099_U27); 
assign R2099_U214 = ~(R2099_U184 & R2099_U159); 
assign R2099_U216 = ~(R2099_U158 & R2099_U208); 
assign R2167_U17 = ~(R2167_U50 & R2167_U49); 
assign R2096_U30 = ~(R2096_U105 & REIP_REG_14__SCAN_IN); 
assign R2096_U174 = ~(R2096_U105 & R2096_U29); 
assign ADD_405_U30 = ~(ADD_405_U108 & INSTADDRPOINTER_REG_14__SCAN_IN); 
assign ADD_405_U178 = ~(ADD_405_U108 & ADD_405_U29); 
assign ADD_515_U30 = ~(ADD_515_U105 & INSTADDRPOINTER_REG_14__SCAN_IN); 
assign ADD_515_U174 = ~(ADD_515_U105 & ADD_515_U29); 
assign U2357 = U5947 & U3853 & R2167_U17; 
assign U2439 = R2182_U42 & U3303; 
assign U2448 = R2167_U17 & U3271; 
assign U2668 = ~(U6755 & U6754 & U3996 & U6751); 
assign U2669 = ~(U6767 & U6766 & U3998 & U6763); 
assign U2765 = ~(U6924 & U6923 & U6925); 
assign U3260 = ~R2167_U17; 
assign U3268 = ~(R2167_U17 & U4485); 
assign U3286 = ~(R2167_U17 & STATE2_REG_3__SCAN_IN); 
assign U4002 = U6781 & U6782 & U6783; 
assign U4003 = U6785 & U6786 & U6787; 
assign U4523 = ~(U2438 & U2442); 
assign U4591 = ~(U2443 & U2438); 
assign U4649 = ~(U2444 & U2438); 
assign U4707 = ~(U2445 & U2438); 
assign U4764 = ~(U2440 & U2442); 
assign U4822 = ~(U2440 & U2443); 
assign U4879 = ~(U2440 & U2444); 
assign U4937 = ~(U2440 & U2445); 
assign U5222 = ~(U2441 & U2442); 
assign U5280 = ~(U2441 & U2443); 
assign U5337 = ~(U2441 & U2444); 
assign U5395 = ~(U2441 & U2445); 
assign U5494 = ~(U5491 & U3735); 
assign U5505 = ~(U2427 & U5502); 
assign U6139 = ~(U4188 & U3270 & R2167_U17); 
assign U6349 = ~(U4190 & R2167_U17); 
assign U6768 = ~(R2182_U27 & U6734); 
assign U7489 = ~(U7481 & R2167_U17); 
assign U7490 = ~(U7481 & U4189 & R2167_U17); 
assign U7669 = ~(U4204 & R2167_U17); 
assign U7686 = ~(R2167_U17 & U7485); 
assign U7731 = ~(R2167_U17 & U7599 & U4420); 
assign R2027_U65 = ~(R2027_U170 & R2027_U169); 
assign R2027_U66 = ~(R2027_U172 & R2027_U171); 
assign R2027_U122 = ~R2027_U46; 
assign R2027_U132 = ~R2027_U102; 
assign R2027_U166 = ~(R2027_U46 & INSTADDRPOINTER_REG_27__SCAN_IN); 
assign R2027_U167 = ~(R2027_U102 & INSTADDRPOINTER_REG_26__SCAN_IN); 
assign R2358_U168 = ~U2667; 
assign R2358_U170 = ~U2670; 
assign R2358_U191 = ~U2658; 
assign R2358_U192 = ~U2659; 
assign R2358_U457 = ~(U2667 & R2358_U22); 
assign R2358_U463 = ~(U2667 & R2358_U22); 
assign R2358_U467 = ~(U2670 & R2358_U22); 
assign R2358_U469 = ~(U2352 & R2358_U171); 
assign R2358_U475 = ~(U2352 & R2358_U171); 
assign R2358_U480 = ~(U2670 & R2358_U22); 
assign R2358_U544 = ~(U2658 & R2358_U22); 
assign R2358_U546 = ~(U2659 & R2358_U22); 
assign R2358_U567 = ~(U2658 & R2358_U22); 
assign R2358_U570 = ~(U2659 & R2358_U22); 
assign R2358_U574 = ~(R2358_U573 & R2358_U572); 
assign R2358_U577 = ~(R2358_U576 & R2358_U575); 
assign R2337_U63 = ~(R2337_U159 & R2337_U158); 
assign R2337_U130 = ~R2337_U45; 
assign R2337_U156 = ~(R2337_U45 & PHYADDRPOINTER_REG_28__SCAN_IN); 
assign R2182_U68 = ~(R2182_U57 & R2182_U39); 
assign R2144_U72 = ~U2766; 
assign R2144_U93 = ~(R2144_U129 & R2144_U113); 
assign R2144_U98 = ~(R2144_U113 & R2144_U112); 
assign R2144_U183 = ~(U2766 & R2144_U12); 
assign R2144_U185 = ~(U2355 & R2144_U73); 
assign R2144_U194 = ~(U2766 & R2144_U12); 
assign R2099_U37 = ~(R2099_U215 & R2099_U214); 
assign R2099_U38 = ~(R2099_U217 & R2099_U216); 
assign R2099_U160 = ~R2099_U109; 
assign R2099_U161 = ~R2099_U10; 
assign R2099_U213 = ~(R2099_U26 & R2099_U109); 
assign R2099_U344 = ~(R2099_U62 & R2099_U10); 
assign R2096_U87 = ~(R2096_U174 & R2096_U173); 
assign R2096_U106 = ~R2096_U30; 
assign R2096_U171 = ~(R2096_U30 & REIP_REG_15__SCAN_IN); 
assign ADD_405_U87 = ~(ADD_405_U178 & ADD_405_U177); 
assign ADD_405_U109 = ~ADD_405_U30; 
assign ADD_405_U175 = ~(ADD_405_U30 & INSTADDRPOINTER_REG_15__SCAN_IN); 
assign ADD_515_U87 = ~(ADD_515_U174 & ADD_515_U173); 
assign ADD_515_U106 = ~ADD_515_U30; 
assign ADD_515_U171 = ~(ADD_515_U30 & INSTADDRPOINTER_REG_15__SCAN_IN); 
assign U2381 = U2357 & U3258; 
assign U2382 = U2357 & U4465; 
assign U2425 = U2368 & U2448; 
assign U2656 = ~(U6780 & U4002); 
assign U2657 = ~(U6784 & U4003); 
assign U3308 = ~(U3293 & U4523); 
assign U3315 = ~(U3311 & U4591); 
assign U3322 = ~(U3317 & U4649); 
assign U3326 = ~(U3324 & U4707); 
assign U3331 = ~(U3328 & U4764); 
assign U3335 = ~(U3333 & U4822); 
assign U3338 = ~(U3336 & U4879); 
assign U3342 = ~(U3340 & U4937); 
assign U3362 = ~(U3360 & U5222); 
assign U3366 = ~(U3364 & U5280); 
assign U3369 = ~(U3367 & U5337); 
assign U3373 = ~(U3371 & U5395); 
assign U3393 = ~(U3258 & U3260); 
assign U3871 = U6139 & U6138; 
assign U4236 = ~(U2451 & U2353 & U3850 & U2448); 
assign U4240 = ~U3286; 
assign U4247 = ~U3268; 
assign U4497 = ~(U2448 & U4250); 
assign U4535 = ~(U4534 & U3284 & U3286); 
assign U4993 = ~(U2439 & U2442); 
assign U5050 = ~(U2439 & U2443); 
assign U5107 = ~(U2439 & U2444); 
assign U5165 = ~(U2439 & U2445); 
assign U5496 = ~(U2427 & U5494); 
assign U6251 = ~(U4186 & U3260); 
assign U6779 = ~(R2337_U63 & U2352); 
assign U7491 = ~(U7490 & U6137); 
assign U7529 = ~(U2357 & U7481); 
assign U7531 = ~(U2357 & U7481); 
assign U7533 = ~(U2357 & U7481); 
assign U7535 = ~(U2357 & U7481); 
assign U7537 = ~(U2357 & U7481); 
assign U7539 = ~(U2357 & U7481); 
assign U7541 = ~(U2357 & U7481); 
assign U7543 = ~(U2357 & U7481); 
assign U7545 = ~(U2357 & U7481); 
assign U7547 = ~(U2357 & U7481); 
assign U7549 = ~(U2357 & U7481); 
assign U7551 = ~(U2357 & U7481); 
assign U7553 = ~(U2357 & U7481); 
assign U7555 = ~(U2357 & U7481); 
assign U7557 = ~(U2357 & U7481); 
assign U7559 = ~(U2357 & U7481); 
assign U7561 = ~(U2357 & U7481); 
assign U7563 = ~(U2357 & U7481); 
assign U7565 = ~(U2357 & U7481); 
assign U7567 = ~(U2357 & U7481); 
assign U7569 = ~(U2357 & U7481); 
assign U7571 = ~(U2357 & U7481); 
assign U7573 = ~(U2357 & U7481); 
assign U7575 = ~(U2357 & U7481); 
assign U7577 = ~(U2357 & U7481); 
assign U7579 = ~(U2357 & U7481); 
assign U7581 = ~(U2357 & U7481); 
assign U7583 = ~(U2357 & U7481); 
assign U7585 = ~(U2357 & U7481); 
assign U7587 = ~(U2357 & U7481); 
assign U7589 = ~(U2357 & U7481); 
assign U7668 = ~(U7489 & U3271); 
assign U7670 = ~(U4494 & U3260); 
assign U7685 = ~(U4204 & U3260); 
assign U7729 = ~(U3258 & U3268); 
assign R2027_U48 = ~(R2027_U94 & R2027_U122); 
assign R2027_U101 = ~(R2027_U122 & INSTADDRPOINTER_REG_27__SCAN_IN); 
assign R2027_U165 = ~(R2027_U122 & R2027_U44); 
assign R2027_U168 = ~(R2027_U132 & R2027_U41); 
assign R2358_U169 = ~U2668; 
assign R2358_U173 = ~U2669; 
assign R2358_U456 = ~(U2352 & R2358_U168); 
assign R2358_U460 = ~(U2668 & R2358_U22); 
assign R2358_U462 = ~(U2352 & R2358_U168); 
assign R2358_U465 = ~(U2668 & R2358_U22); 
assign R2358_U466 = ~(U2352 & R2358_U170); 
assign R2358_U471 = ~(R2358_U470 & R2358_U469); 
assign R2358_U479 = ~(U2352 & R2358_U170); 
assign R2358_U482 = ~(U2669 & R2358_U22); 
assign R2358_U484 = ~(U2669 & R2358_U22); 
assign R2358_U543 = ~(U2352 & R2358_U191); 
assign R2358_U545 = ~(U2352 & R2358_U192); 
assign R2358_U566 = ~(U2352 & R2358_U191); 
assign R2358_U569 = ~(U2352 & R2358_U192); 
assign R2337_U47 = ~(R2337_U130 & PHYADDRPOINTER_REG_28__SCAN_IN); 
assign R2337_U157 = ~(R2337_U130 & R2337_U46); 
assign R2182_U26 = ~(R2182_U68 & R2182_U67); 
assign R2144_U28 = ~(R2144_U186 & R2144_U185); 
assign R2144_U75 = ~U2765; 
assign R2144_U130 = ~R2144_U93; 
assign R2144_U148 = ~R2144_U98; 
assign R2144_U182 = ~(U2355 & R2144_U72); 
assign R2144_U193 = ~(U2355 & R2144_U72); 
assign R2144_U196 = ~(U2765 & R2144_U12); 
assign R2144_U198 = ~(U2765 & R2144_U12); 
assign R2144_U259 = ~(U2355 & R2144_U98); 
assign R2099_U11 = ~(R2099_U92 & R2099_U161); 
assign R2099_U144 = ~(R2099_U161 & R2099_U62); 
assign R2099_U212 = ~(R2099_U160 & R2099_U211); 
assign R2099_U343 = ~(R2099_U261 & R2099_U161); 
assign R2096_U32 = ~(R2096_U106 & REIP_REG_15__SCAN_IN); 
assign R2096_U172 = ~(R2096_U106 & R2096_U31); 
assign ADD_405_U32 = ~(ADD_405_U109 & INSTADDRPOINTER_REG_15__SCAN_IN); 
assign ADD_405_U176 = ~(ADD_405_U109 & ADD_405_U31); 
assign ADD_515_U32 = ~(ADD_515_U106 & INSTADDRPOINTER_REG_15__SCAN_IN); 
assign ADD_515_U172 = ~(ADD_515_U106 & ADD_515_U31); 
assign U2473 = U7668 & U7667 & U3393; 
assign U3287 = ~(U4535 & U3281); 
assign U3348 = ~(U3343 & U4993); 
assign U3352 = ~(U3350 & U5050); 
assign U3355 = ~(U3353 & U5107); 
assign U3359 = ~(U3357 & U5165); 
assign U3403 = ~(U3851 & U4236); 
assign U4001 = U6777 & U6778 & U6779; 
assign U4170 = ~(U7686 & U7685 & U3726); 
assign U4248 = ~U3393; 
assign U4496 = ~(U7670 & U7669 & U4495); 
assign U4509 = ~(U4240 & U4249); 
assign U4524 = ~U3308; 
assign U4592 = ~U3315; 
assign U4650 = ~U3322; 
assign U4708 = ~U3326; 
assign U4765 = ~U3331; 
assign U4823 = ~U3335; 
assign U4880 = ~U3338; 
assign U4938 = ~U3342; 
assign U5223 = ~U3362; 
assign U5281 = ~U3366; 
assign U5338 = ~U3369; 
assign U5396 = ~U3373; 
assign U5495 = ~(U4240 & U3425); 
assign U5504 = ~(U4240 & U3388); 
assign U5515 = ~(U5507 & U4240); 
assign U5520 = ~(U4240 & U3253); 
assign U5948 = ~(U2382 & EAX_REG_15__SCAN_IN); 
assign U5949 = ~(DATAI_15_ & U2381); 
assign U5951 = ~(U2382 & EAX_REG_14__SCAN_IN); 
assign U5952 = ~(DATAI_14_ & U2381); 
assign U5954 = ~(U2382 & EAX_REG_13__SCAN_IN); 
assign U5955 = ~(DATAI_13_ & U2381); 
assign U5957 = ~(U2382 & EAX_REG_12__SCAN_IN); 
assign U5958 = ~(DATAI_12_ & U2381); 
assign U5960 = ~(U2382 & EAX_REG_11__SCAN_IN); 
assign U5961 = ~(DATAI_11_ & U2381); 
assign U5963 = ~(U2382 & EAX_REG_10__SCAN_IN); 
assign U5964 = ~(DATAI_10_ & U2381); 
assign U5966 = ~(U2382 & EAX_REG_9__SCAN_IN); 
assign U5967 = ~(DATAI_9_ & U2381); 
assign U5969 = ~(U2382 & EAX_REG_8__SCAN_IN); 
assign U5970 = ~(DATAI_8_ & U2381); 
assign U5972 = ~(U2382 & EAX_REG_7__SCAN_IN); 
assign U5973 = ~(U2381 & DATAI_7_); 
assign U5975 = ~(U2382 & EAX_REG_6__SCAN_IN); 
assign U5976 = ~(U2381 & DATAI_6_); 
assign U5978 = ~(U2382 & EAX_REG_5__SCAN_IN); 
assign U5979 = ~(U2381 & DATAI_5_); 
assign U5981 = ~(U2382 & EAX_REG_4__SCAN_IN); 
assign U5982 = ~(U2381 & DATAI_4_); 
assign U5984 = ~(U2382 & EAX_REG_3__SCAN_IN); 
assign U5985 = ~(U2381 & DATAI_3_); 
assign U5987 = ~(U2382 & EAX_REG_2__SCAN_IN); 
assign U5988 = ~(U2381 & DATAI_2_); 
assign U5990 = ~(U2382 & EAX_REG_1__SCAN_IN); 
assign U5991 = ~(U2381 & DATAI_1_); 
assign U5993 = ~(U2382 & EAX_REG_0__SCAN_IN); 
assign U5994 = ~(U2381 & DATAI_0_); 
assign U5996 = ~(U2382 & EAX_REG_30__SCAN_IN); 
assign U5997 = ~(DATAI_14_ & U2381); 
assign U5999 = ~(U2382 & EAX_REG_29__SCAN_IN); 
assign U6000 = ~(DATAI_13_ & U2381); 
assign U6002 = ~(U2382 & EAX_REG_28__SCAN_IN); 
assign U6003 = ~(DATAI_12_ & U2381); 
assign U6005 = ~(U2382 & EAX_REG_27__SCAN_IN); 
assign U6006 = ~(DATAI_11_ & U2381); 
assign U6008 = ~(U2382 & EAX_REG_26__SCAN_IN); 
assign U6009 = ~(DATAI_10_ & U2381); 
assign U6011 = ~(U2382 & EAX_REG_25__SCAN_IN); 
assign U6012 = ~(DATAI_9_ & U2381); 
assign U6014 = ~(U2382 & EAX_REG_24__SCAN_IN); 
assign U6015 = ~(DATAI_8_ & U2381); 
assign U6017 = ~(U2382 & EAX_REG_23__SCAN_IN); 
assign U6018 = ~(U2381 & DATAI_7_); 
assign U6020 = ~(U2382 & EAX_REG_22__SCAN_IN); 
assign U6021 = ~(U2381 & DATAI_6_); 
assign U6023 = ~(U2382 & EAX_REG_21__SCAN_IN); 
assign U6024 = ~(U2381 & DATAI_5_); 
assign U6026 = ~(U2382 & EAX_REG_20__SCAN_IN); 
assign U6027 = ~(U2381 & DATAI_4_); 
assign U6029 = ~(U2382 & EAX_REG_19__SCAN_IN); 
assign U6030 = ~(U2381 & DATAI_3_); 
assign U6032 = ~(U2382 & EAX_REG_18__SCAN_IN); 
assign U6033 = ~(U2381 & DATAI_2_); 
assign U6035 = ~(U2382 & EAX_REG_17__SCAN_IN); 
assign U6036 = ~(U2381 & DATAI_1_); 
assign U6038 = ~(U2382 & EAX_REG_16__SCAN_IN); 
assign U6039 = ~(U2381 & DATAI_0_); 
assign U6041 = ~(U4223 & U7594 & U4247); 
assign U6140 = ~(U7491 & U3244); 
assign U6252 = ~(U4193 & U6251); 
assign U6604 = ~(U4487 & U3957 & U3393); 
assign U6759 = ~(R2182_U26 & U6734); 
assign U7486 = ~(U2425 & U7481); 
assign U7487 = ~(U2425 & U7481); 
assign U7530 = ~(U7529 & UWORD_REG_0__SCAN_IN); 
assign U7532 = ~(U7531 & UWORD_REG_1__SCAN_IN); 
assign U7534 = ~(U7533 & UWORD_REG_2__SCAN_IN); 
assign U7536 = ~(U7535 & UWORD_REG_3__SCAN_IN); 
assign U7538 = ~(U7537 & UWORD_REG_4__SCAN_IN); 
assign U7540 = ~(U7539 & UWORD_REG_5__SCAN_IN); 
assign U7542 = ~(U7541 & UWORD_REG_6__SCAN_IN); 
assign U7544 = ~(U7543 & UWORD_REG_7__SCAN_IN); 
assign U7546 = ~(U7545 & UWORD_REG_8__SCAN_IN); 
assign U7548 = ~(U7547 & UWORD_REG_9__SCAN_IN); 
assign U7550 = ~(U7549 & UWORD_REG_10__SCAN_IN); 
assign U7552 = ~(U7551 & UWORD_REG_11__SCAN_IN); 
assign U7554 = ~(U7553 & UWORD_REG_12__SCAN_IN); 
assign U7556 = ~(U7555 & UWORD_REG_13__SCAN_IN); 
assign U7558 = ~(U7557 & UWORD_REG_14__SCAN_IN); 
assign U7560 = ~(U7559 & LWORD_REG_0__SCAN_IN); 
assign U7562 = ~(U7561 & LWORD_REG_1__SCAN_IN); 
assign U7564 = ~(U7563 & LWORD_REG_2__SCAN_IN); 
assign U7566 = ~(U7565 & LWORD_REG_3__SCAN_IN); 
assign U7568 = ~(U7567 & LWORD_REG_4__SCAN_IN); 
assign U7570 = ~(U7569 & LWORD_REG_5__SCAN_IN); 
assign U7572 = ~(U7571 & LWORD_REG_6__SCAN_IN); 
assign U7574 = ~(U7573 & LWORD_REG_7__SCAN_IN); 
assign U7576 = ~(U7575 & LWORD_REG_8__SCAN_IN); 
assign U7578 = ~(U7577 & LWORD_REG_9__SCAN_IN); 
assign U7580 = ~(U7579 & LWORD_REG_10__SCAN_IN); 
assign U7582 = ~(U7581 & LWORD_REG_11__SCAN_IN); 
assign U7584 = ~(U7583 & LWORD_REG_12__SCAN_IN); 
assign U7586 = ~(U7585 & LWORD_REG_13__SCAN_IN); 
assign U7588 = ~(U7587 & LWORD_REG_14__SCAN_IN); 
assign U7590 = ~(U7589 & LWORD_REG_15__SCAN_IN); 
assign U7591 = ~(U7481 & U3556 & U4247); 
assign U7730 = ~(U7729 & U7728 & U3244 & U4159); 
assign R2027_U63 = ~(R2027_U166 & R2027_U165); 
assign R2027_U64 = ~(R2027_U168 & R2027_U167); 
assign R2027_U123 = ~R2027_U48; 
assign R2027_U131 = ~R2027_U101; 
assign R2027_U162 = ~(R2027_U48 & INSTADDRPOINTER_REG_29__SCAN_IN); 
assign R2027_U163 = ~(R2027_U101 & INSTADDRPOINTER_REG_28__SCAN_IN); 
assign R2358_U198 = ~U2656; 
assign R2358_U199 = ~U2657; 
assign R2358_U458 = ~(R2358_U457 & R2358_U456); 
assign R2358_U459 = ~(U2352 & R2358_U169); 
assign R2358_U464 = ~(U2352 & R2358_U169); 
assign R2358_U468 = ~(R2358_U467 & R2358_U466); 
assign R2358_U481 = ~(U2352 & R2358_U173); 
assign R2358_U483 = ~(U2352 & R2358_U173); 
assign R2358_U559 = ~(U2656 & R2358_U22); 
assign R2358_U561 = ~(U2657 & R2358_U22); 
assign R2358_U568 = ~(R2358_U567 & R2358_U566); 
assign R2358_U571 = ~(R2358_U570 & R2358_U569); 
assign R2358_U582 = ~(U2657 & R2358_U22); 
assign R2358_U585 = ~(U2656 & R2358_U22); 
assign R2337_U62 = ~(R2337_U157 & R2337_U156); 
assign R2337_U131 = ~R2337_U47; 
assign R2337_U154 = ~(R2337_U47 & PHYADDRPOINTER_REG_29__SCAN_IN); 
assign R2144_U100 = ~(U2751 & R2144_U28); 
assign R2144_U109 = ~(R2144_U194 & R2144_U193 & R2144_U13); 
assign R2144_U184 = ~(R2144_U183 & R2144_U182); 
assign R2144_U187 = ~R2144_U28; 
assign R2144_U195 = ~(U2355 & R2144_U75); 
assign R2144_U197 = ~(U2355 & R2144_U75); 
assign R2144_U241 = ~(R2144_U28 & R2144_U14); 
assign R2144_U243 = ~(R2144_U28 & R2144_U14); 
assign R2144_U260 = ~(R2144_U148 & R2144_U12); 
assign R2099_U36 = ~(R2099_U213 & R2099_U212); 
assign R2099_U85 = ~(R2099_U344 & R2099_U343); 
assign R2099_U162 = ~R2099_U144; 
assign R2099_U163 = ~R2099_U11; 
assign R2099_U340 = ~(R2099_U60 & R2099_U11); 
assign R2099_U342 = ~(R2099_U63 & R2099_U144); 
assign R2096_U86 = ~(R2096_U172 & R2096_U171); 
assign R2096_U107 = ~R2096_U32; 
assign R2096_U169 = ~(R2096_U32 & REIP_REG_16__SCAN_IN); 
assign ADD_405_U86 = ~(ADD_405_U176 & ADD_405_U175); 
assign ADD_405_U110 = ~ADD_405_U32; 
assign ADD_405_U173 = ~(ADD_405_U32 & INSTADDRPOINTER_REG_16__SCAN_IN); 
assign ADD_515_U86 = ~(ADD_515_U172 & ADD_515_U171); 
assign ADD_515_U107 = ~ADD_515_U32; 
assign ADD_515_U169 = ~(ADD_515_U32 & INSTADDRPOINTER_REG_16__SCAN_IN); 
assign U2364 = U3852 & U3403; 
assign U2365 = U4249 & U3403; 
assign U2372 = U3403 & STATE2_REG_0__SCAN_IN; 
assign U2376 = U5786 & U3403; 
assign U2655 = ~(U6776 & U4001); 
assign U3272 = ~(U2473 & U4489); 
assign U3404 = ~(U6042 & U6041); 
assign U3413 = ~(U4223 & U6252); 
assign U3569 = U7591 & STATE2_REG_2__SCAN_IN; 
assign U4166 = ~(U4496 & U3378); 
assign U4212 = ~U3287; 
assign U4994 = ~U3348; 
assign U5051 = ~U3352; 
assign U5108 = ~U3355; 
assign U5166 = ~U3359; 
assign U5461 = ~U4170; 
assign U5462 = ~(U2368 & U4170); 
assign U5497 = ~(U5496 & U5495); 
assign U5506 = ~(U5505 & U5503 & U5504); 
assign U5517 = ~(U5516 & U5514 & U5515); 
assign U5523 = ~(U5521 & U5522 & U5520); 
assign U5547 = ~(U4248 & U2431); 
assign U5783 = ~U3403; 
assign U5950 = ~(U5949 & U5948); 
assign U5953 = ~(U5952 & U5951); 
assign U5956 = ~(U5955 & U5954); 
assign U5959 = ~(U5958 & U5957); 
assign U5962 = ~(U5961 & U5960); 
assign U5965 = ~(U5964 & U5963); 
assign U5968 = ~(U5967 & U5966); 
assign U5971 = ~(U5970 & U5969); 
assign U5974 = ~(U5973 & U5972); 
assign U5977 = ~(U5976 & U5975); 
assign U5980 = ~(U5979 & U5978); 
assign U5983 = ~(U5982 & U5981); 
assign U5986 = ~(U5985 & U5984); 
assign U5989 = ~(U5988 & U5987); 
assign U5992 = ~(U5991 & U5990); 
assign U5995 = ~(U5994 & U5993); 
assign U5998 = ~(U5997 & U5996); 
assign U6001 = ~(U6000 & U5999); 
assign U6004 = ~(U6003 & U6002); 
assign U6007 = ~(U6006 & U6005); 
assign U6010 = ~(U6009 & U6008); 
assign U6013 = ~(U6012 & U6011); 
assign U6016 = ~(U6015 & U6014); 
assign U6019 = ~(U6018 & U6017); 
assign U6022 = ~(U6021 & U6020); 
assign U6025 = ~(U6024 & U6023); 
assign U6028 = ~(U6027 & U6026); 
assign U6031 = ~(U6030 & U6029); 
assign U6034 = ~(U6033 & U6032); 
assign U6037 = ~(U6036 & U6035); 
assign U6040 = ~(U6039 & U6038); 
assign U6141 = ~(U3871 & U6140); 
assign U6598 = ~(U2368 & U2473); 
assign U6605 = ~(U6604 & MEMORYFETCH_REG_SCAN_IN); 
assign U6775 = ~(R2337_U62 & U2352); 
assign U7488 = ~(U6349 & U6348 & U7487); 
assign U7762 = ~(U3475 & U4170); 
assign U7765 = ~(U5494 & U4170); 
assign U7767 = ~(U5502 & U4170); 
assign U7769 = ~(U5513 & U4170); 
assign U7771 = ~(U5519 & U4170); 
assign R2027_U49 = ~(R2027_U123 & INSTADDRPOINTER_REG_29__SCAN_IN); 
assign R2027_U161 = ~(R2027_U123 & R2027_U47); 
assign R2027_U164 = ~(R2027_U131 & R2027_U45); 
assign R2358_U461 = ~(R2358_U460 & R2358_U459); 
assign R2358_U485 = ~(R2358_U484 & R2358_U483); 
assign R2358_U558 = ~(U2352 & R2358_U198); 
assign R2358_U560 = ~(U2352 & R2358_U199); 
assign R2358_U581 = ~(U2352 & R2358_U199); 
assign R2358_U584 = ~(U2352 & R2358_U198); 
assign R2337_U49 = ~(R2337_U131 & PHYADDRPOINTER_REG_29__SCAN_IN); 
assign R2337_U155 = ~(R2337_U131 & R2337_U48); 
assign R2144_U43 = ~(R2144_U260 & R2144_U259); 
assign R2144_U55 = R2144_U109 & R2144_U106; 
assign R2144_U110 = ~(R2144_U196 & R2144_U195 & R2144_U16); 
assign R2144_U114 = ~(R2144_U187 & R2144_U14); 
assign R2144_U116 = ~(U2750 & R2144_U184); 
assign R2144_U131 = ~(R2144_U187 & R2144_U14); 
assign R2144_U154 = ~(R2144_U113 & R2144_U115 & R2144_U100); 
assign R2144_U157 = ~(U2750 & R2144_U184); 
assign R2144_U162 = ~(U2750 & R2144_U184); 
assign R2144_U199 = ~(R2144_U198 & R2144_U197); 
assign R2144_U240 = ~(R2144_U187 & U2751); 
assign R2144_U242 = ~(R2144_U187 & U2751); 
assign R2099_U12 = ~(R2099_U93 & R2099_U163); 
assign R2099_U143 = ~(R2099_U163 & R2099_U60); 
assign R2099_U339 = ~(R2099_U267 & R2099_U163); 
assign R2099_U341 = ~(R2099_U162 & R2099_U264); 
assign R2096_U34 = ~(R2096_U107 & REIP_REG_16__SCAN_IN); 
assign R2096_U170 = ~(R2096_U107 & R2096_U33); 
assign ADD_405_U34 = ~(ADD_405_U110 & INSTADDRPOINTER_REG_16__SCAN_IN); 
assign ADD_405_U174 = ~(ADD_405_U110 & ADD_405_U33); 
assign ADD_515_U34 = ~(ADD_515_U107 & INSTADDRPOINTER_REG_16__SCAN_IN); 
assign ADD_515_U170 = ~(ADD_515_U107 & ADD_515_U33); 
assign U2358 = U2388 & U4212; 
assign U2361 = U4212 & STATE2_REG_3__SCAN_IN; 
assign U2384 = U3404 & STATE2_REG_0__SCAN_IN; 
assign U2385 = U3404 & U3281; 
assign U2390 = DATAI_0_ & U4212; 
assign U2391 = DATAI_1_ & U4212; 
assign U2392 = DATAI_2_ & U4212; 
assign U2393 = DATAI_3_ & U4212; 
assign U2394 = DATAI_4_ & U4212; 
assign U2395 = DATAI_5_ & U4212; 
assign U2396 = DATAI_6_ & U4212; 
assign U2397 = DATAI_7_ & U4212; 
assign U2788 = ~(U6605 & U3419 & U7486); 
assign U3296 = ~R2144_U43; 
assign U3411 = ~(U4223 & U6141); 
assign U3575 = U4540 & U4541 & U4212; 
assign U3584 = U4598 & U4599 & U4212; 
assign U3593 = U4657 & U4658 & U4212; 
assign U3602 = U4714 & U4715 & U4212; 
assign U3611 = U4772 & U4773 & U4212; 
assign U3620 = U4829 & U4830 & U4212; 
assign U3629 = U4887 & U4888 & U4212; 
assign U3638 = U4944 & U4945 & U4212; 
assign U3647 = U5000 & U5001 & U4212; 
assign U3656 = U5057 & U5058 & U4212; 
assign U3665 = U5115 & U5116 & U4212; 
assign U3674 = U5172 & U5173 & U4212; 
assign U3683 = U5230 & U5231 & U4212; 
assign U3692 = U5287 & U5288 & U4212; 
assign U3701 = U5345 & U5346 & U4212; 
assign U3710 = U5402 & U5403 & U4212; 
assign U4000 = U6773 & U6774 & U6775; 
assign U4160 = ~(U3727 & U5462); 
assign U4165 = ~(U2368 & U3272); 
assign U4210 = ~U3413; 
assign U4216 = ~(U4223 & U7488); 
assign U4225 = ~U4166; 
assign U4490 = ~U3272; 
assign U5544 = ~(R2144_U43 & U4197); 
assign U5548 = ~(U2518 & U5547 & U7731 & U7730); 
assign U5787 = ~(U2376 & PHYADDRPOINTER_REG_0__SCAN_IN); 
assign U5789 = ~(U2365 & REIP_REG_0__SCAN_IN); 
assign U5791 = ~(U5783 & PHYADDRPOINTER_REG_0__SCAN_IN); 
assign U5792 = ~(R2337_U5 & U2376); 
assign U5794 = ~(U2365 & REIP_REG_1__SCAN_IN); 
assign U5796 = ~(U5783 & PHYADDRPOINTER_REG_1__SCAN_IN); 
assign U5797 = ~(R2337_U60 & U2376); 
assign U5799 = ~(U2365 & REIP_REG_2__SCAN_IN); 
assign U5801 = ~(U5783 & PHYADDRPOINTER_REG_2__SCAN_IN); 
assign U5802 = ~(R2337_U57 & U2376); 
assign U5804 = ~(U2365 & REIP_REG_3__SCAN_IN); 
assign U5806 = ~(U5783 & PHYADDRPOINTER_REG_3__SCAN_IN); 
assign U5807 = ~(R2337_U56 & U2376); 
assign U5809 = ~(U2365 & REIP_REG_4__SCAN_IN); 
assign U5811 = ~(U5783 & PHYADDRPOINTER_REG_4__SCAN_IN); 
assign U5812 = ~(R2337_U55 & U2376); 
assign U5814 = ~(U2365 & REIP_REG_5__SCAN_IN); 
assign U5816 = ~(U5783 & PHYADDRPOINTER_REG_5__SCAN_IN); 
assign U5817 = ~(R2337_U54 & U2376); 
assign U5819 = ~(U2365 & REIP_REG_6__SCAN_IN); 
assign U5821 = ~(U5783 & PHYADDRPOINTER_REG_6__SCAN_IN); 
assign U5822 = ~(R2337_U53 & U2376); 
assign U5824 = ~(U2365 & REIP_REG_7__SCAN_IN); 
assign U5826 = ~(U5783 & PHYADDRPOINTER_REG_7__SCAN_IN); 
assign U5827 = ~(R2337_U52 & U2376); 
assign U5829 = ~(U2365 & REIP_REG_8__SCAN_IN); 
assign U5831 = ~(U5783 & PHYADDRPOINTER_REG_8__SCAN_IN); 
assign U5832 = ~(R2337_U51 & U2376); 
assign U5834 = ~(U2365 & REIP_REG_9__SCAN_IN); 
assign U5836 = ~(U5783 & PHYADDRPOINTER_REG_9__SCAN_IN); 
assign U5837 = ~(R2337_U80 & U2376); 
assign U5839 = ~(U2365 & REIP_REG_10__SCAN_IN); 
assign U5841 = ~(U5783 & PHYADDRPOINTER_REG_10__SCAN_IN); 
assign U5842 = ~(R2337_U79 & U2376); 
assign U5844 = ~(U2365 & REIP_REG_11__SCAN_IN); 
assign U5846 = ~(U5783 & PHYADDRPOINTER_REG_11__SCAN_IN); 
assign U5847 = ~(R2337_U78 & U2376); 
assign U5849 = ~(U2365 & REIP_REG_12__SCAN_IN); 
assign U5851 = ~(U5783 & PHYADDRPOINTER_REG_12__SCAN_IN); 
assign U5852 = ~(R2337_U77 & U2376); 
assign U5854 = ~(U2365 & REIP_REG_13__SCAN_IN); 
assign U5856 = ~(U5783 & PHYADDRPOINTER_REG_13__SCAN_IN); 
assign U5857 = ~(R2337_U76 & U2376); 
assign U5859 = ~(U2365 & REIP_REG_14__SCAN_IN); 
assign U5861 = ~(U5783 & PHYADDRPOINTER_REG_14__SCAN_IN); 
assign U5862 = ~(R2337_U75 & U2376); 
assign U5864 = ~(U2365 & REIP_REG_15__SCAN_IN); 
assign U5866 = ~(U5783 & PHYADDRPOINTER_REG_15__SCAN_IN); 
assign U5867 = ~(R2337_U74 & U2376); 
assign U5869 = ~(U2365 & REIP_REG_16__SCAN_IN); 
assign U5871 = ~(U5783 & PHYADDRPOINTER_REG_16__SCAN_IN); 
assign U5872 = ~(R2337_U73 & U2376); 
assign U5874 = ~(U2365 & REIP_REG_17__SCAN_IN); 
assign U5876 = ~(U5783 & PHYADDRPOINTER_REG_17__SCAN_IN); 
assign U5877 = ~(R2337_U72 & U2376); 
assign U5879 = ~(U2365 & REIP_REG_18__SCAN_IN); 
assign U5881 = ~(U5783 & PHYADDRPOINTER_REG_18__SCAN_IN); 
assign U5882 = ~(R2337_U71 & U2376); 
assign U5884 = ~(U2365 & REIP_REG_19__SCAN_IN); 
assign U5886 = ~(U5783 & PHYADDRPOINTER_REG_19__SCAN_IN); 
assign U5887 = ~(R2337_U70 & U2376); 
assign U5889 = ~(U2365 & REIP_REG_20__SCAN_IN); 
assign U5891 = ~(U5783 & PHYADDRPOINTER_REG_20__SCAN_IN); 
assign U5892 = ~(R2337_U69 & U2376); 
assign U5894 = ~(U2365 & REIP_REG_21__SCAN_IN); 
assign U5896 = ~(U5783 & PHYADDRPOINTER_REG_21__SCAN_IN); 
assign U5897 = ~(R2337_U68 & U2376); 
assign U5899 = ~(U2365 & REIP_REG_22__SCAN_IN); 
assign U5901 = ~(U5783 & PHYADDRPOINTER_REG_22__SCAN_IN); 
assign U5902 = ~(R2337_U67 & U2376); 
assign U5904 = ~(U2365 & REIP_REG_23__SCAN_IN); 
assign U5906 = ~(U5783 & PHYADDRPOINTER_REG_23__SCAN_IN); 
assign U5907 = ~(R2337_U66 & U2376); 
assign U5909 = ~(U2365 & REIP_REG_24__SCAN_IN); 
assign U5911 = ~(U5783 & PHYADDRPOINTER_REG_24__SCAN_IN); 
assign U5912 = ~(R2337_U65 & U2376); 
assign U5914 = ~(U2365 & REIP_REG_25__SCAN_IN); 
assign U5916 = ~(U5783 & PHYADDRPOINTER_REG_25__SCAN_IN); 
assign U5917 = ~(R2337_U64 & U2376); 
assign U5919 = ~(U2365 & REIP_REG_26__SCAN_IN); 
assign U5921 = ~(U5783 & PHYADDRPOINTER_REG_26__SCAN_IN); 
assign U5922 = ~(R2337_U63 & U2376); 
assign U5924 = ~(U2365 & REIP_REG_27__SCAN_IN); 
assign U5926 = ~(U5783 & PHYADDRPOINTER_REG_27__SCAN_IN); 
assign U5927 = ~(R2337_U62 & U2376); 
assign U5929 = ~(U2365 & REIP_REG_28__SCAN_IN); 
assign U5931 = ~(U5783 & PHYADDRPOINTER_REG_28__SCAN_IN); 
assign U5934 = ~(U2365 & REIP_REG_29__SCAN_IN); 
assign U5936 = ~(U5783 & PHYADDRPOINTER_REG_29__SCAN_IN); 
assign U5939 = ~(U2365 & REIP_REG_30__SCAN_IN); 
assign U5941 = ~(U5783 & PHYADDRPOINTER_REG_30__SCAN_IN); 
assign U5944 = ~(U2365 & REIP_REG_31__SCAN_IN); 
assign U5946 = ~(U5783 & PHYADDRPOINTER_REG_31__SCAN_IN); 
assign U6043 = ~U3404; 
assign U6255 = ~(U3413 & EBX_REG_0__SCAN_IN); 
assign U6258 = ~(U3413 & EBX_REG_1__SCAN_IN); 
assign U6261 = ~(U3413 & EBX_REG_2__SCAN_IN); 
assign U6264 = ~(U3413 & EBX_REG_3__SCAN_IN); 
assign U6267 = ~(U3413 & EBX_REG_4__SCAN_IN); 
assign U6270 = ~(U3413 & EBX_REG_5__SCAN_IN); 
assign U6273 = ~(U3413 & EBX_REG_6__SCAN_IN); 
assign U6276 = ~(U3413 & EBX_REG_7__SCAN_IN); 
assign U6279 = ~(U3413 & EBX_REG_8__SCAN_IN); 
assign U6282 = ~(U3413 & EBX_REG_9__SCAN_IN); 
assign U6285 = ~(U3413 & EBX_REG_10__SCAN_IN); 
assign U6288 = ~(U3413 & EBX_REG_11__SCAN_IN); 
assign U6291 = ~(U3413 & EBX_REG_12__SCAN_IN); 
assign U6294 = ~(U3413 & EBX_REG_13__SCAN_IN); 
assign U6297 = ~(U3413 & EBX_REG_14__SCAN_IN); 
assign U6300 = ~(U3413 & EBX_REG_15__SCAN_IN); 
assign U6303 = ~(U3413 & EBX_REG_16__SCAN_IN); 
assign U6306 = ~(U3413 & EBX_REG_17__SCAN_IN); 
assign U6309 = ~(U3413 & EBX_REG_18__SCAN_IN); 
assign U6312 = ~(U3413 & EBX_REG_19__SCAN_IN); 
assign U6315 = ~(U3413 & EBX_REG_20__SCAN_IN); 
assign U6318 = ~(U3413 & EBX_REG_21__SCAN_IN); 
assign U6321 = ~(U3413 & EBX_REG_22__SCAN_IN); 
assign U6324 = ~(U3413 & EBX_REG_23__SCAN_IN); 
assign U6327 = ~(U3413 & EBX_REG_24__SCAN_IN); 
assign U6330 = ~(U3413 & EBX_REG_25__SCAN_IN); 
assign U6333 = ~(U3413 & EBX_REG_26__SCAN_IN); 
assign U6336 = ~(U3413 & EBX_REG_27__SCAN_IN); 
assign U6339 = ~(U3413 & EBX_REG_28__SCAN_IN); 
assign U6342 = ~(U3413 & EBX_REG_29__SCAN_IN); 
assign U6345 = ~(U3413 & EBX_REG_30__SCAN_IN); 
assign U6347 = ~(U3413 & EBX_REG_31__SCAN_IN); 
assign U6599 = ~(U6598 & CODEFETCH_REG_SCAN_IN); 
assign U6877 = ~(U4147 & R2144_U43); 
assign U7498 = ~(U7481 & U5950); 
assign U7499 = ~(U7481 & U5953); 
assign U7500 = ~(U7481 & U5956); 
assign U7501 = ~(U7481 & U5959); 
assign U7502 = ~(U7481 & U5962); 
assign U7503 = ~(U7481 & U5965); 
assign U7504 = ~(U7481 & U5968); 
assign U7505 = ~(U7481 & U5971); 
assign U7506 = ~(U7481 & U5974); 
assign U7507 = ~(U7481 & U5977); 
assign U7508 = ~(U7481 & U5980); 
assign U7509 = ~(U7481 & U5983); 
assign U7510 = ~(U7481 & U5986); 
assign U7511 = ~(U7481 & U5989); 
assign U7512 = ~(U7481 & U5992); 
assign U7513 = ~(U7481 & U5995); 
assign U7514 = ~(U7481 & U5998); 
assign U7515 = ~(U7481 & U6001); 
assign U7516 = ~(U7481 & U6004); 
assign U7517 = ~(U7481 & U6007); 
assign U7518 = ~(U7481 & U6010); 
assign U7519 = ~(U7481 & U6013); 
assign U7520 = ~(U7481 & U6016); 
assign U7521 = ~(U7481 & U6019); 
assign U7522 = ~(U7481 & U6022); 
assign U7523 = ~(U7481 & U6025); 
assign U7524 = ~(U7481 & U6028); 
assign U7525 = ~(U7481 & U6031); 
assign U7526 = ~(U7481 & U6034); 
assign U7527 = ~(U7481 & U6037); 
assign U7528 = ~(U7481 & U6040); 
assign U7763 = ~(U5461 & INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign U7764 = ~(U5461 & INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign U7766 = ~(U5461 & INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign U7768 = ~(U5461 & INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U7770 = ~(U5461 & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign R2027_U61 = ~(R2027_U162 & R2027_U161); 
assign R2027_U62 = ~(R2027_U164 & R2027_U163); 
assign R2027_U128 = ~R2027_U49; 
assign R2027_U157 = ~(R2027_U49 & INSTADDRPOINTER_REG_30__SCAN_IN); 
assign R2358_U197 = ~U2655; 
assign R2358_U557 = ~(U2655 & R2358_U22); 
assign R2358_U583 = ~(R2358_U582 & R2358_U581); 
assign R2358_U586 = ~(R2358_U585 & R2358_U584); 
assign R2358_U588 = ~(U2655 & R2358_U22); 
assign R2337_U61 = ~(R2337_U155 & R2337_U154); 
assign R2337_U132 = ~R2337_U49; 
assign R2337_U150 = ~(R2337_U49 & PHYADDRPOINTER_REG_30__SCAN_IN); 
assign R2144_U48 = R2144_U162 & R2144_U109; 
assign R2144_U51 = R2144_U110 & R2144_U109; 
assign R2144_U92 = R2144_U241 & R2144_U240; 
assign R2144_U111 = ~(U2749 & R2144_U199); 
assign R2144_U132 = ~(R2144_U131 & R2144_U93); 
assign R2144_U155 = ~(R2144_U154 & R2144_U114); 
assign R2144_U159 = ~(U2749 & R2144_U106 & R2144_U199); 
assign R2144_U161 = ~(U2749 & R2144_U199); 
assign R2144_U163 = ~(R2144_U116 & R2144_U109); 
assign R2144_U244 = ~(R2144_U243 & R2144_U242); 
assign R2099_U83 = ~(R2099_U340 & R2099_U339); 
assign R2099_U84 = ~(R2099_U342 & R2099_U341); 
assign R2099_U164 = ~R2099_U143; 
assign R2099_U165 = ~R2099_U12; 
assign R2099_U336 = ~(R2099_U58 & R2099_U12); 
assign R2099_U338 = ~(R2099_U61 & R2099_U143); 
assign R2096_U85 = ~(R2096_U170 & R2096_U169); 
assign R2096_U108 = ~R2096_U34; 
assign R2096_U167 = ~(R2096_U34 & REIP_REG_17__SCAN_IN); 
assign ADD_405_U85 = ~(ADD_405_U174 & ADD_405_U173); 
assign ADD_405_U111 = ~ADD_405_U34; 
assign ADD_405_U171 = ~(ADD_405_U34 & INSTADDRPOINTER_REG_17__SCAN_IN); 
assign ADD_515_U85 = ~(ADD_515_U170 & ADD_515_U169); 
assign ADD_515_U108 = ~ADD_515_U34; 
assign ADD_515_U167 = ~(ADD_515_U34 & INSTADDRPOINTER_REG_17__SCAN_IN); 
assign U2371 = U4210 & U4437; 
assign U2383 = U4210 & U3378; 
assign U2398 = DATAI_24_ & U2358; 
assign U2399 = DATAI_16_ & U2358; 
assign U2400 = DATAI_25_ & U2358; 
assign U2401 = DATAI_17_ & U2358; 
assign U2402 = DATAI_26_ & U2358; 
assign U2403 = DATAI_18_ & U2358; 
assign U2404 = DATAI_27_ & U2358; 
assign U2405 = DATAI_19_ & U2358; 
assign U2406 = DATAI_28_ & U2358; 
assign U2407 = DATAI_20_ & U2358; 
assign U2408 = DATAI_29_ & U2358; 
assign U2409 = DATAI_21_ & U2358; 
assign U2410 = DATAI_30_ & U2358; 
assign U2411 = DATAI_22_ & U2358; 
assign U2412 = DATAI_31_ & U2358; 
assign U2413 = DATAI_23_ & U2358; 
assign U2414 = U2361 & U3258; 
assign U2415 = U2361 & U3378; 
assign U2416 = U2361 & U3264; 
assign U2417 = U2361 & U3271; 
assign U2418 = U2361 & U3270; 
assign U2419 = U2361 & U3265; 
assign U2420 = U2361 & U4161; 
assign U2421 = U2361 & U4159; 
assign U2424 = U2384 & U3271; 
assign U2654 = ~(U6772 & U4000); 
assign U2787 = ~(U6878 & U6879 & U6877); 
assign U2790 = ~(U6600 & U6599); 
assign U2892 = U6043 & DATAO_REG_31__SCAN_IN; 
assign U2924 = ~(U7528 & U7530); 
assign U2925 = ~(U7527 & U7532); 
assign U2926 = ~(U7526 & U7534); 
assign U2927 = ~(U7525 & U7536); 
assign U2928 = ~(U7524 & U7538); 
assign U2929 = ~(U7523 & U7540); 
assign U2930 = ~(U7522 & U7542); 
assign U2931 = ~(U7521 & U7544); 
assign U2932 = ~(U7520 & U7546); 
assign U2933 = ~(U7519 & U7548); 
assign U2934 = ~(U7518 & U7550); 
assign U2935 = ~(U7517 & U7552); 
assign U2936 = ~(U7516 & U7554); 
assign U2937 = ~(U7515 & U7556); 
assign U2938 = ~(U7514 & U7558); 
assign U2939 = ~(U7513 & U7560); 
assign U2940 = ~(U7512 & U7562); 
assign U2941 = ~(U7511 & U7564); 
assign U2942 = ~(U7510 & U7566); 
assign U2943 = ~(U7509 & U7568); 
assign U2944 = ~(U7508 & U7570); 
assign U2945 = ~(U7507 & U7572); 
assign U2946 = ~(U7506 & U7574); 
assign U2947 = ~(U7505 & U7576); 
assign U2948 = ~(U7504 & U7578); 
assign U2949 = ~(U7503 & U7580); 
assign U2950 = ~(U7502 & U7582); 
assign U2951 = ~(U7501 & U7584); 
assign U2952 = ~(U7500 & U7586); 
assign U2953 = ~(U7499 & U7588); 
assign U2954 = ~(U7498 & U7590); 
assign U3418 = ~(U4216 & U3875); 
assign U3476 = ~(U7763 & U7762); 
assign U3477 = ~(U7765 & U7764); 
assign U3478 = ~(U7767 & U7766); 
assign U3479 = ~(U7769 & U7768); 
assign U3480 = ~(U7771 & U7770); 
assign U4168 = ~(U3955 & U4216); 
assign U4169 = ~(U4216 & U3419); 
assign U4211 = ~U3411; 
assign U5464 = ~U4160; 
assign U5550 = ~(U2368 & U5548); 
assign U5932 = ~(R2337_U61 & U2376); 
assign U6044 = ~(U2385 & LWORD_REG_0__SCAN_IN); 
assign U6045 = ~(U2384 & EAX_REG_0__SCAN_IN); 
assign U6046 = ~(U6043 & DATAO_REG_0__SCAN_IN); 
assign U6047 = ~(U2385 & LWORD_REG_1__SCAN_IN); 
assign U6048 = ~(U2384 & EAX_REG_1__SCAN_IN); 
assign U6049 = ~(U6043 & DATAO_REG_1__SCAN_IN); 
assign U6050 = ~(U2385 & LWORD_REG_2__SCAN_IN); 
assign U6051 = ~(U2384 & EAX_REG_2__SCAN_IN); 
assign U6052 = ~(U6043 & DATAO_REG_2__SCAN_IN); 
assign U6053 = ~(U2385 & LWORD_REG_3__SCAN_IN); 
assign U6054 = ~(U2384 & EAX_REG_3__SCAN_IN); 
assign U6055 = ~(U6043 & DATAO_REG_3__SCAN_IN); 
assign U6056 = ~(U2385 & LWORD_REG_4__SCAN_IN); 
assign U6057 = ~(U2384 & EAX_REG_4__SCAN_IN); 
assign U6058 = ~(U6043 & DATAO_REG_4__SCAN_IN); 
assign U6059 = ~(U2385 & LWORD_REG_5__SCAN_IN); 
assign U6060 = ~(U2384 & EAX_REG_5__SCAN_IN); 
assign U6061 = ~(U6043 & DATAO_REG_5__SCAN_IN); 
assign U6062 = ~(U2385 & LWORD_REG_6__SCAN_IN); 
assign U6063 = ~(U2384 & EAX_REG_6__SCAN_IN); 
assign U6064 = ~(U6043 & DATAO_REG_6__SCAN_IN); 
assign U6065 = ~(U2385 & LWORD_REG_7__SCAN_IN); 
assign U6066 = ~(U2384 & EAX_REG_7__SCAN_IN); 
assign U6067 = ~(U6043 & DATAO_REG_7__SCAN_IN); 
assign U6068 = ~(U2385 & LWORD_REG_8__SCAN_IN); 
assign U6069 = ~(U2384 & EAX_REG_8__SCAN_IN); 
assign U6070 = ~(U6043 & DATAO_REG_8__SCAN_IN); 
assign U6071 = ~(U2385 & LWORD_REG_9__SCAN_IN); 
assign U6072 = ~(U2384 & EAX_REG_9__SCAN_IN); 
assign U6073 = ~(U6043 & DATAO_REG_9__SCAN_IN); 
assign U6074 = ~(U2385 & LWORD_REG_10__SCAN_IN); 
assign U6075 = ~(U2384 & EAX_REG_10__SCAN_IN); 
assign U6076 = ~(U6043 & DATAO_REG_10__SCAN_IN); 
assign U6077 = ~(U2385 & LWORD_REG_11__SCAN_IN); 
assign U6078 = ~(U2384 & EAX_REG_11__SCAN_IN); 
assign U6079 = ~(U6043 & DATAO_REG_11__SCAN_IN); 
assign U6080 = ~(U2385 & LWORD_REG_12__SCAN_IN); 
assign U6081 = ~(U2384 & EAX_REG_12__SCAN_IN); 
assign U6082 = ~(U6043 & DATAO_REG_12__SCAN_IN); 
assign U6083 = ~(U2385 & LWORD_REG_13__SCAN_IN); 
assign U6084 = ~(U2384 & EAX_REG_13__SCAN_IN); 
assign U6085 = ~(U6043 & DATAO_REG_13__SCAN_IN); 
assign U6086 = ~(U2385 & LWORD_REG_14__SCAN_IN); 
assign U6087 = ~(U2384 & EAX_REG_14__SCAN_IN); 
assign U6088 = ~(U6043 & DATAO_REG_14__SCAN_IN); 
assign U6089 = ~(U2385 & LWORD_REG_15__SCAN_IN); 
assign U6090 = ~(U2384 & EAX_REG_15__SCAN_IN); 
assign U6091 = ~(U6043 & DATAO_REG_15__SCAN_IN); 
assign U6093 = ~(U2385 & UWORD_REG_0__SCAN_IN); 
assign U6094 = ~(U6043 & DATAO_REG_16__SCAN_IN); 
assign U6096 = ~(U2385 & UWORD_REG_1__SCAN_IN); 
assign U6097 = ~(U6043 & DATAO_REG_17__SCAN_IN); 
assign U6099 = ~(U2385 & UWORD_REG_2__SCAN_IN); 
assign U6100 = ~(U6043 & DATAO_REG_18__SCAN_IN); 
assign U6102 = ~(U2385 & UWORD_REG_3__SCAN_IN); 
assign U6103 = ~(U6043 & DATAO_REG_19__SCAN_IN); 
assign U6105 = ~(U2385 & UWORD_REG_4__SCAN_IN); 
assign U6106 = ~(U6043 & DATAO_REG_20__SCAN_IN); 
assign U6108 = ~(U2385 & UWORD_REG_5__SCAN_IN); 
assign U6109 = ~(U6043 & DATAO_REG_21__SCAN_IN); 
assign U6111 = ~(U2385 & UWORD_REG_6__SCAN_IN); 
assign U6112 = ~(U6043 & DATAO_REG_22__SCAN_IN); 
assign U6114 = ~(U2385 & UWORD_REG_7__SCAN_IN); 
assign U6115 = ~(U6043 & DATAO_REG_23__SCAN_IN); 
assign U6117 = ~(U2385 & UWORD_REG_8__SCAN_IN); 
assign U6118 = ~(U6043 & DATAO_REG_24__SCAN_IN); 
assign U6120 = ~(U2385 & UWORD_REG_9__SCAN_IN); 
assign U6121 = ~(U6043 & DATAO_REG_25__SCAN_IN); 
assign U6123 = ~(U2385 & UWORD_REG_10__SCAN_IN); 
assign U6124 = ~(U6043 & DATAO_REG_26__SCAN_IN); 
assign U6126 = ~(U2385 & UWORD_REG_11__SCAN_IN); 
assign U6127 = ~(U6043 & DATAO_REG_27__SCAN_IN); 
assign U6129 = ~(U2385 & UWORD_REG_12__SCAN_IN); 
assign U6130 = ~(U6043 & DATAO_REG_28__SCAN_IN); 
assign U6132 = ~(U2385 & UWORD_REG_13__SCAN_IN); 
assign U6133 = ~(U6043 & DATAO_REG_29__SCAN_IN); 
assign U6135 = ~(U2385 & UWORD_REG_14__SCAN_IN); 
assign U6136 = ~(U6043 & DATAO_REG_30__SCAN_IN); 
assign U6144 = ~(U3411 & EAX_REG_0__SCAN_IN); 
assign U6147 = ~(U3411 & EAX_REG_1__SCAN_IN); 
assign U6150 = ~(U3411 & EAX_REG_2__SCAN_IN); 
assign U6153 = ~(U3411 & EAX_REG_3__SCAN_IN); 
assign U6156 = ~(U3411 & EAX_REG_4__SCAN_IN); 
assign U6159 = ~(U3411 & EAX_REG_5__SCAN_IN); 
assign U6162 = ~(U3411 & EAX_REG_6__SCAN_IN); 
assign U6165 = ~(U3411 & EAX_REG_7__SCAN_IN); 
assign U6168 = ~(U3411 & EAX_REG_8__SCAN_IN); 
assign U6171 = ~(U3411 & EAX_REG_9__SCAN_IN); 
assign U6174 = ~(U3411 & EAX_REG_10__SCAN_IN); 
assign U6177 = ~(U3411 & EAX_REG_11__SCAN_IN); 
assign U6180 = ~(U3411 & EAX_REG_12__SCAN_IN); 
assign U6183 = ~(U3411 & EAX_REG_13__SCAN_IN); 
assign U6186 = ~(U3411 & EAX_REG_14__SCAN_IN); 
assign U6189 = ~(U3411 & EAX_REG_15__SCAN_IN); 
assign U6193 = ~(U3411 & EAX_REG_16__SCAN_IN); 
assign U6197 = ~(U3411 & EAX_REG_17__SCAN_IN); 
assign U6201 = ~(U3411 & EAX_REG_18__SCAN_IN); 
assign U6205 = ~(U3411 & EAX_REG_19__SCAN_IN); 
assign U6209 = ~(U3411 & EAX_REG_20__SCAN_IN); 
assign U6213 = ~(U3411 & EAX_REG_21__SCAN_IN); 
assign U6217 = ~(U3411 & EAX_REG_22__SCAN_IN); 
assign U6221 = ~(U3411 & EAX_REG_23__SCAN_IN); 
assign U6225 = ~(U3411 & EAX_REG_24__SCAN_IN); 
assign U6229 = ~(U3411 & EAX_REG_25__SCAN_IN); 
assign U6233 = ~(U3411 & EAX_REG_26__SCAN_IN); 
assign U6237 = ~(U3411 & EAX_REG_27__SCAN_IN); 
assign U6241 = ~(U3411 & EAX_REG_28__SCAN_IN); 
assign U6245 = ~(U3411 & EAX_REG_29__SCAN_IN); 
assign U6249 = ~(U3411 & EAX_REG_30__SCAN_IN); 
assign U6588 = ~U4165; 
assign U6589 = ~(U4165 & FLUSH_REG_SCAN_IN); 
assign U6771 = ~(R2337_U61 & U2352); 
assign U6858 = ~(U3426 & U4448 & U3296); 
assign U7614 = ~(U4490 & U4498); 
assign U7689 = ~(U3454 & U4160); 
assign U7697 = ~(U5497 & U4160); 
assign U7710 = ~(U5506 & U4160); 
assign U7712 = ~(U5517 & U4160); 
assign U7716 = ~(U5523 & U4160); 
assign U7732 = ~(U3411 & EAX_REG_31__SCAN_IN); 
assign U7750 = ~(U4165 & MORE_REG_SCAN_IN); 
assign R2027_U99 = ~(R2027_U128 & INSTADDRPOINTER_REG_30__SCAN_IN); 
assign R2027_U158 = ~(R2027_U128 & R2027_U50); 
assign R2358_U556 = ~(U2352 & R2358_U197); 
assign R2358_U587 = ~(U2352 & R2358_U197); 
assign R2337_U96 = ~(R2337_U132 & PHYADDRPOINTER_REG_30__SCAN_IN); 
assign R2337_U151 = ~(R2337_U132 & R2337_U50); 
assign R2144_U56 = R2144_U159 & R2144_U19; 
assign R2144_U58 = R2144_U19 & R2144_U21 & R2144_U159; 
assign R2144_U62 = R2144_U111 & R2144_U110; 
assign R2144_U91 = ~(R2144_U100 & R2144_U132); 
assign R2144_U117 = ~(R2144_U155 & R2144_U157); 
assign R2144_U137 = ~(R2144_U161 & R2144_U110); 
assign R2144_U245 = ~(R2144_U92 & R2144_U93); 
assign R2144_U246 = ~(R2144_U130 & R2144_U244); 
assign R2099_U13 = ~(R2099_U94 & R2099_U165); 
assign R2099_U142 = ~(R2099_U165 & R2099_U58); 
assign R2099_U335 = ~(R2099_U273 & R2099_U165); 
assign R2099_U337 = ~(R2099_U164 & R2099_U270); 
assign R2096_U36 = ~(R2096_U108 & REIP_REG_17__SCAN_IN); 
assign R2096_U168 = ~(R2096_U108 & R2096_U35); 
assign ADD_405_U36 = ~(ADD_405_U111 & INSTADDRPOINTER_REG_17__SCAN_IN); 
assign ADD_405_U172 = ~(ADD_405_U111 & ADD_405_U35); 
assign ADD_515_U36 = ~(ADD_515_U108 & INSTADDRPOINTER_REG_17__SCAN_IN); 
assign ADD_515_U168 = ~(ADD_515_U108 & ADD_515_U35); 
assign U2359 = U3418 & STATE2_REG_2__SCAN_IN; 
assign U2373 = U3418 & STATE2_REG_3__SCAN_IN; 
assign U2386 = U4211 & U3410; 
assign U2387 = U3872 & U4211; 
assign U2422 = U4211 & U5449; 
assign U2423 = U4211 & U4219; 
assign U2426 = U3877 & U3418; 
assign U2650 = U6858 & STATE2_REG_2__SCAN_IN; 
assign U2793 = ~(U6589 & U4236); 
assign U2908 = ~(U6090 & U6089 & U6091); 
assign U2909 = ~(U6087 & U6086 & U6088); 
assign U2910 = ~(U6084 & U6083 & U6085); 
assign U2911 = ~(U6081 & U6080 & U6082); 
assign U2912 = ~(U6078 & U6077 & U6079); 
assign U2913 = ~(U6075 & U6074 & U6076); 
assign U2914 = ~(U6072 & U6071 & U6073); 
assign U2915 = ~(U6069 & U6068 & U6070); 
assign U2916 = ~(U6066 & U6065 & U6067); 
assign U2917 = ~(U6063 & U6062 & U6064); 
assign U2918 = ~(U6060 & U6059 & U6061); 
assign U2919 = ~(U6057 & U6056 & U6058); 
assign U2920 = ~(U6054 & U6053 & U6055); 
assign U2921 = ~(U6051 & U6050 & U6052); 
assign U2922 = ~(U6048 & U6047 & U6049); 
assign U2923 = ~(U6045 & U6044 & U6046); 
assign U3401 = ~(U3744 & U5550); 
assign U3856 = U6093 & U6094; 
assign U3857 = U6096 & U6097; 
assign U3858 = U6099 & U6100; 
assign U3859 = U6102 & U6103; 
assign U3860 = U6105 & U6106; 
assign U3861 = U6108 & U6109; 
assign U3862 = U6111 & U6112; 
assign U3863 = U6114 & U6115; 
assign U3864 = U6117 & U6118; 
assign U3865 = U6120 & U6121; 
assign U3866 = U6123 & U6124; 
assign U3867 = U6126 & U6127; 
assign U3868 = U6129 & U6130; 
assign U3869 = U6132 & U6133; 
assign U3870 = U6135 & U6136; 
assign U3999 = U6769 & U6770 & U6771; 
assign U4215 = ~(U4243 & U3418); 
assign U4548 = ~(U2415 & U4522); 
assign U4553 = ~(U2416 & U4522); 
assign U4558 = ~(U2420 & U4522); 
assign U4563 = ~(U2419 & U4522); 
assign U4568 = ~(U2418 & U4522); 
assign U4573 = ~(U2421 & U4522); 
assign U4578 = ~(U2414 & U4522); 
assign U4583 = ~(U2417 & U4522); 
assign U4606 = ~(U4590 & U2415); 
assign U4611 = ~(U4590 & U2416); 
assign U4616 = ~(U4590 & U2420); 
assign U4621 = ~(U4590 & U2419); 
assign U4626 = ~(U4590 & U2418); 
assign U4631 = ~(U4590 & U2421); 
assign U4636 = ~(U4590 & U2414); 
assign U4641 = ~(U4590 & U2417); 
assign U4665 = ~(U4648 & U2415); 
assign U4670 = ~(U4648 & U2416); 
assign U4675 = ~(U4648 & U2420); 
assign U4680 = ~(U4648 & U2419); 
assign U4685 = ~(U4648 & U2418); 
assign U4690 = ~(U4648 & U2421); 
assign U4695 = ~(U4648 & U2414); 
assign U4700 = ~(U4648 & U2417); 
assign U4722 = ~(U4706 & U2415); 
assign U4727 = ~(U4706 & U2416); 
assign U4732 = ~(U4706 & U2420); 
assign U4737 = ~(U4706 & U2419); 
assign U4742 = ~(U4706 & U2418); 
assign U4747 = ~(U4706 & U2421); 
assign U4752 = ~(U4706 & U2414); 
assign U4757 = ~(U4706 & U2417); 
assign U4780 = ~(U4763 & U2415); 
assign U4785 = ~(U4763 & U2416); 
assign U4790 = ~(U4763 & U2420); 
assign U4795 = ~(U4763 & U2419); 
assign U4800 = ~(U4763 & U2418); 
assign U4805 = ~(U4763 & U2421); 
assign U4810 = ~(U4763 & U2414); 
assign U4815 = ~(U4763 & U2417); 
assign U4837 = ~(U4821 & U2415); 
assign U4842 = ~(U4821 & U2416); 
assign U4847 = ~(U4821 & U2420); 
assign U4852 = ~(U4821 & U2419); 
assign U4857 = ~(U4821 & U2418); 
assign U4862 = ~(U4821 & U2421); 
assign U4867 = ~(U4821 & U2414); 
assign U4872 = ~(U4821 & U2417); 
assign U4895 = ~(U4878 & U2415); 
assign U4900 = ~(U4878 & U2416); 
assign U4905 = ~(U4878 & U2420); 
assign U4910 = ~(U4878 & U2419); 
assign U4915 = ~(U4878 & U2418); 
assign U4920 = ~(U4878 & U2421); 
assign U4925 = ~(U4878 & U2414); 
assign U4930 = ~(U4878 & U2417); 
assign U4952 = ~(U4936 & U2415); 
assign U4957 = ~(U4936 & U2416); 
assign U4962 = ~(U4936 & U2420); 
assign U4967 = ~(U4936 & U2419); 
assign U4972 = ~(U4936 & U2418); 
assign U4977 = ~(U4936 & U2421); 
assign U4982 = ~(U4936 & U2414); 
assign U4987 = ~(U4936 & U2417); 
assign U5008 = ~(U4525 & U2415); 
assign U5013 = ~(U4525 & U2416); 
assign U5018 = ~(U4525 & U2420); 
assign U5023 = ~(U4525 & U2419); 
assign U5028 = ~(U4525 & U2418); 
assign U5033 = ~(U4525 & U2421); 
assign U5038 = ~(U4525 & U2414); 
assign U5043 = ~(U4525 & U2417); 
assign U5065 = ~(U5049 & U2415); 
assign U5070 = ~(U5049 & U2416); 
assign U5075 = ~(U5049 & U2420); 
assign U5080 = ~(U5049 & U2419); 
assign U5085 = ~(U5049 & U2418); 
assign U5090 = ~(U5049 & U2421); 
assign U5095 = ~(U5049 & U2414); 
assign U5100 = ~(U5049 & U2417); 
assign U5123 = ~(U5106 & U2415); 
assign U5128 = ~(U5106 & U2416); 
assign U5133 = ~(U5106 & U2420); 
assign U5138 = ~(U5106 & U2419); 
assign U5143 = ~(U5106 & U2418); 
assign U5148 = ~(U5106 & U2421); 
assign U5153 = ~(U5106 & U2414); 
assign U5158 = ~(U5106 & U2417); 
assign U5180 = ~(U5164 & U2415); 
assign U5185 = ~(U5164 & U2416); 
assign U5190 = ~(U5164 & U2420); 
assign U5195 = ~(U5164 & U2419); 
assign U5200 = ~(U5164 & U2418); 
assign U5205 = ~(U5164 & U2421); 
assign U5210 = ~(U5164 & U2414); 
assign U5215 = ~(U5164 & U2417); 
assign U5238 = ~(U5221 & U2415); 
assign U5243 = ~(U5221 & U2416); 
assign U5248 = ~(U5221 & U2420); 
assign U5253 = ~(U5221 & U2419); 
assign U5258 = ~(U5221 & U2418); 
assign U5263 = ~(U5221 & U2421); 
assign U5268 = ~(U5221 & U2414); 
assign U5273 = ~(U5221 & U2417); 
assign U5295 = ~(U5279 & U2415); 
assign U5300 = ~(U5279 & U2416); 
assign U5305 = ~(U5279 & U2420); 
assign U5310 = ~(U5279 & U2419); 
assign U5315 = ~(U5279 & U2418); 
assign U5320 = ~(U5279 & U2421); 
assign U5325 = ~(U5279 & U2414); 
assign U5330 = ~(U5279 & U2417); 
assign U5353 = ~(U5336 & U2415); 
assign U5358 = ~(U5336 & U2416); 
assign U5363 = ~(U5336 & U2420); 
assign U5368 = ~(U5336 & U2419); 
assign U5373 = ~(U5336 & U2418); 
assign U5378 = ~(U5336 & U2421); 
assign U5383 = ~(U5336 & U2414); 
assign U5388 = ~(U5336 & U2417); 
assign U5410 = ~(U5394 & U2415); 
assign U5415 = ~(U5394 & U2416); 
assign U5420 = ~(U5394 & U2420); 
assign U5425 = ~(U5394 & U2419); 
assign U5429 = ~(U5394 & U2418); 
assign U5434 = ~(U5394 & U2421); 
assign U5439 = ~(U5394 & U2414); 
assign U5444 = ~(U5394 & U2417); 
assign U6092 = ~(U2424 & EAX_REG_16__SCAN_IN); 
assign U6095 = ~(U2424 & EAX_REG_17__SCAN_IN); 
assign U6098 = ~(U2424 & EAX_REG_18__SCAN_IN); 
assign U6101 = ~(U2424 & EAX_REG_19__SCAN_IN); 
assign U6104 = ~(U2424 & EAX_REG_20__SCAN_IN); 
assign U6107 = ~(U2424 & EAX_REG_21__SCAN_IN); 
assign U6110 = ~(U2424 & EAX_REG_22__SCAN_IN); 
assign U6113 = ~(U2424 & EAX_REG_23__SCAN_IN); 
assign U6116 = ~(U2424 & EAX_REG_24__SCAN_IN); 
assign U6119 = ~(U2424 & EAX_REG_25__SCAN_IN); 
assign U6122 = ~(U2424 & EAX_REG_26__SCAN_IN); 
assign U6125 = ~(U2424 & EAX_REG_27__SCAN_IN); 
assign U6128 = ~(U2424 & EAX_REG_28__SCAN_IN); 
assign U6131 = ~(U2424 & EAX_REG_29__SCAN_IN); 
assign U6134 = ~(U2424 & EAX_REG_30__SCAN_IN); 
assign U6254 = ~(U2371 & R2099_U86); 
assign U6257 = ~(U2371 & R2099_U87); 
assign U6260 = ~(U2371 & R2099_U138); 
assign U6263 = ~(U2371 & R2099_U42); 
assign U6266 = ~(U2371 & R2099_U41); 
assign U6269 = ~(U2371 & R2099_U40); 
assign U6272 = ~(U2371 & R2099_U39); 
assign U6275 = ~(U2371 & R2099_U38); 
assign U6278 = ~(U2371 & R2099_U37); 
assign U6281 = ~(U2371 & R2099_U36); 
assign U6284 = ~(U2371 & R2099_U85); 
assign U6287 = ~(U2371 & R2099_U84); 
assign U6290 = ~(U2371 & R2099_U83); 
assign U6351 = ~U3418; 
assign U6591 = ~U4168; 
assign U6602 = ~U4169; 
assign U7446 = ~(U3476 & U3249); 
assign U7448 = ~(U3477 & U3249); 
assign U7451 = ~(U3478 & U3249); 
assign U7454 = ~(U3479 & U3249); 
assign U7690 = ~(U5464 & INSTQUEUERD_ADDR_REG_4__SCAN_IN); 
assign U7696 = ~(U5464 & INSTQUEUERD_ADDR_REG_3__SCAN_IN); 
assign U7709 = ~(U5464 & INSTQUEUERD_ADDR_REG_2__SCAN_IN); 
assign U7711 = ~(U5464 & INSTQUEUERD_ADDR_REG_1__SCAN_IN); 
assign U7715 = ~(U5464 & INSTQUEUERD_ADDR_REG_0__SCAN_IN); 
assign U7751 = ~(U4225 & U6588); 
assign U7755 = ~(U6597 & U4168); 
assign U7761 = ~(U6603 & U4169); 
assign U7781 = ~(U3480 & U3249); 
assign R2027_U59 = ~(R2027_U158 & R2027_U157); 
assign R2027_U129 = ~R2027_U99; 
assign R2027_U155 = ~(R2027_U99 & INSTADDRPOINTER_REG_31__SCAN_IN); 
assign R2278_U19 = ~(U2787 & INSTADDRPOINTER_REG_0__SCAN_IN); 
assign R2278_U292 = U2787 | INSTADDRPOINTER_REG_0__SCAN_IN; 
assign R2358_U196 = ~U2654; 
assign R2358_U555 = ~(U2654 & R2358_U22); 
assign R2358_U589 = ~(R2358_U588 & R2358_U587); 
assign R2358_U591 = ~(U2654 & R2358_U22); 
assign R2337_U59 = ~(R2337_U151 & R2337_U150); 
assign R2337_U133 = ~R2337_U96; 
assign R2337_U148 = ~(R2337_U96 & PHYADDRPOINTER_REG_31__SCAN_IN); 
assign R2144_U50 = ~(R2144_U246 & R2144_U245); 
assign R2144_U118 = ~(R2144_U51 & R2144_U117); 
assign R2144_U133 = ~R2144_U91; 
assign R2144_U134 = ~(R2144_U91 & R2144_U109); 
assign R2144_U158 = ~(R2144_U117 & R2144_U110 & R2144_U55); 
assign R2144_U238 = ~(R2144_U163 & R2144_U91); 
assign R2099_U81 = ~(R2099_U336 & R2099_U335); 
assign R2099_U82 = ~(R2099_U338 & R2099_U337); 
assign R2099_U166 = ~R2099_U142; 
assign R2099_U167 = ~R2099_U13; 
assign R2099_U332 = ~(R2099_U56 & R2099_U13); 
assign R2099_U334 = ~(R2099_U59 & R2099_U142); 
assign R2096_U84 = ~(R2096_U168 & R2096_U167); 
assign R2096_U109 = ~R2096_U36; 
assign R2096_U165 = ~(R2096_U36 & REIP_REG_18__SCAN_IN); 
assign LT_563_U8 = ~U3478; 
assign LT_563_U9 = ~U3477; 
assign LT_563_U12 = ~U3476; 
assign LT_563_U15 = ~U3479; 
assign LT_563_U16 = ~U3480; 
assign LT_563_U21 = ~(U3478 & LT_563_U7); 
assign LT_563_U22 = ~(U3477 & LT_563_U10); 
assign LT_563_U27 = ~(U3476 & LT_563_U11); 
assign ADD_405_U84 = ~(ADD_405_U172 & ADD_405_U171); 
assign ADD_405_U112 = ~ADD_405_U36; 
assign ADD_405_U169 = ~(ADD_405_U36 & INSTADDRPOINTER_REG_18__SCAN_IN); 
assign ADD_515_U84 = ~(ADD_515_U168 & ADD_515_U167); 
assign ADD_515_U109 = ~ADD_515_U36; 
assign ADD_515_U165 = ~(ADD_515_U36 & INSTADDRPOINTER_REG_18__SCAN_IN); 
assign U2360 = U3401 & STATE2_REG_2__SCAN_IN; 
assign U2362 = U2359 & U4196; 
assign U2363 = U2359 & U4198; 
assign U2370 = U3401 & U3250; 
assign U2377 = U3750 & U3401; 
assign U2486 = ~(R2144_U43 | R2144_U50); 
assign U2649 = R2144_U50 & U6734; 
assign U2653 = ~(U6768 & U3999); 
assign U2673 = ~(U7446 & U7445); 
assign U2674 = ~(U7448 & U7447); 
assign U2675 = ~(U4156 & U7451); 
assign U2676 = ~(U4157 & U7454); 
assign U2677 = ~(U7782 & U7781 & U7455); 
assign U2893 = ~(U3870 & U6134); 
assign U2894 = ~(U3869 & U6131); 
assign U2895 = ~(U3868 & U6128); 
assign U2896 = ~(U3867 & U6125); 
assign U2897 = ~(U3866 & U6122); 
assign U2898 = ~(U3865 & U6119); 
assign U2899 = ~(U3864 & U6116); 
assign U2900 = ~(U3863 & U6113); 
assign U2901 = ~(U3862 & U6110); 
assign U2902 = ~(U3861 & U6107); 
assign U2903 = ~(U3860 & U6104); 
assign U2904 = ~(U3859 & U6101); 
assign U2905 = ~(U3858 & U6098); 
assign U2906 = ~(U3857 & U6095); 
assign U2907 = ~(U3856 & U6092); 
assign U3297 = ~R2144_U50; 
assign U3300 = ~(R2144_U50 & R2144_U43); 
assign U3312 = ~(R2144_U50 & U3296); 
assign U3455 = ~(U7690 & U7689); 
assign U3456 = ~(U7697 & U7696); 
assign U3459 = ~(U7710 & U7709); 
assign U3460 = ~(U7712 & U7711); 
assign U3461 = ~(U7716 & U7715); 
assign U3471 = ~(U7751 & U7750); 
assign U5541 = ~(U4214 & R2144_U50); 
assign U5552 = ~U3401; 
assign U5937 = ~(R2337_U59 & U2376); 
assign U6142 = ~(U2422 & DATAI_0_); 
assign U6145 = ~(U2422 & DATAI_1_); 
assign U6148 = ~(U2422 & DATAI_2_); 
assign U6151 = ~(U2422 & DATAI_3_); 
assign U6154 = ~(U2422 & DATAI_4_); 
assign U6157 = ~(U2422 & DATAI_5_); 
assign U6160 = ~(U2422 & DATAI_6_); 
assign U6163 = ~(U2422 & DATAI_7_); 
assign U6166 = ~(U2422 & DATAI_8_); 
assign U6169 = ~(U2422 & DATAI_9_); 
assign U6172 = ~(U2422 & DATAI_10_); 
assign U6175 = ~(U2422 & DATAI_11_); 
assign U6178 = ~(U2422 & DATAI_12_); 
assign U6181 = ~(U2422 & DATAI_13_); 
assign U6184 = ~(U2422 & DATAI_14_); 
assign U6187 = ~(U2422 & DATAI_15_); 
assign U6190 = ~(U2423 & DATAI_16_); 
assign U6191 = ~(U2387 & DATAI_0_); 
assign U6194 = ~(U2423 & DATAI_17_); 
assign U6195 = ~(U2387 & DATAI_1_); 
assign U6198 = ~(U2423 & DATAI_18_); 
assign U6199 = ~(U2387 & DATAI_2_); 
assign U6202 = ~(U2423 & DATAI_19_); 
assign U6203 = ~(U2387 & DATAI_3_); 
assign U6206 = ~(U2423 & DATAI_20_); 
assign U6207 = ~(U2387 & DATAI_4_); 
assign U6210 = ~(U2423 & DATAI_21_); 
assign U6211 = ~(U2387 & DATAI_5_); 
assign U6214 = ~(U2423 & DATAI_22_); 
assign U6215 = ~(U2387 & DATAI_6_); 
assign U6218 = ~(U2423 & DATAI_23_); 
assign U6219 = ~(U2387 & DATAI_7_); 
assign U6222 = ~(U2423 & DATAI_24_); 
assign U6223 = ~(U2387 & DATAI_8_); 
assign U6226 = ~(U2423 & DATAI_25_); 
assign U6227 = ~(U2387 & DATAI_9_); 
assign U6230 = ~(U2423 & DATAI_26_); 
assign U6231 = ~(U2387 & DATAI_10_); 
assign U6234 = ~(U2423 & DATAI_27_); 
assign U6235 = ~(U2387 & DATAI_11_); 
assign U6238 = ~(U2423 & DATAI_28_); 
assign U6239 = ~(U2387 & DATAI_12_); 
assign U6242 = ~(U2423 & DATAI_29_); 
assign U6243 = ~(U2387 & DATAI_13_); 
assign U6246 = ~(U2423 & DATAI_30_); 
assign U6247 = ~(U2387 & DATAI_14_); 
assign U6250 = ~(U2423 & DATAI_31_); 
assign U6293 = ~(U2371 & R2099_U82); 
assign U6296 = ~(U2371 & R2099_U81); 
assign U6360 = ~(U2426 & R2182_U34); 
assign U6361 = ~(U2373 & PHYADDRPOINTER_REG_0__SCAN_IN); 
assign U6363 = ~(U6351 & REIP_REG_0__SCAN_IN); 
assign U6368 = ~(U2426 & R2182_U33); 
assign U6369 = ~(U2373 & PHYADDRPOINTER_REG_1__SCAN_IN); 
assign U6371 = ~(U6351 & REIP_REG_1__SCAN_IN); 
assign U6376 = ~(U2426 & R2182_U42); 
assign U6377 = ~(U2373 & PHYADDRPOINTER_REG_2__SCAN_IN); 
assign U6379 = ~(U6351 & REIP_REG_2__SCAN_IN); 
assign U6384 = ~(U2426 & R2182_U25); 
assign U6385 = ~(U2373 & PHYADDRPOINTER_REG_3__SCAN_IN); 
assign U6387 = ~(U6351 & REIP_REG_3__SCAN_IN); 
assign U6392 = ~(U2426 & R2182_U24); 
assign U6393 = ~(U2373 & PHYADDRPOINTER_REG_4__SCAN_IN); 
assign U6395 = ~(U6351 & REIP_REG_4__SCAN_IN); 
assign U6400 = ~(R2182_U5 & U2426); 
assign U6401 = ~(U2373 & PHYADDRPOINTER_REG_5__SCAN_IN); 
assign U6403 = ~(U6351 & REIP_REG_5__SCAN_IN); 
assign U6407 = ~(U2373 & PHYADDRPOINTER_REG_6__SCAN_IN); 
assign U6410 = ~(U6351 & REIP_REG_6__SCAN_IN); 
assign U6414 = ~(U2373 & PHYADDRPOINTER_REG_7__SCAN_IN); 
assign U6417 = ~(U6351 & REIP_REG_7__SCAN_IN); 
assign U6421 = ~(U2373 & PHYADDRPOINTER_REG_8__SCAN_IN); 
assign U6424 = ~(U6351 & REIP_REG_8__SCAN_IN); 
assign U6428 = ~(U2373 & PHYADDRPOINTER_REG_9__SCAN_IN); 
assign U6431 = ~(U6351 & REIP_REG_9__SCAN_IN); 
assign U6435 = ~(U2373 & PHYADDRPOINTER_REG_10__SCAN_IN); 
assign U6438 = ~(U6351 & REIP_REG_10__SCAN_IN); 
assign U6442 = ~(U2373 & PHYADDRPOINTER_REG_11__SCAN_IN); 
assign U6445 = ~(U6351 & REIP_REG_11__SCAN_IN); 
assign U6449 = ~(U2373 & PHYADDRPOINTER_REG_12__SCAN_IN); 
assign U6452 = ~(U6351 & REIP_REG_12__SCAN_IN); 
assign U6456 = ~(U2373 & PHYADDRPOINTER_REG_13__SCAN_IN); 
assign U6459 = ~(U6351 & REIP_REG_13__SCAN_IN); 
assign U6463 = ~(U2373 & PHYADDRPOINTER_REG_14__SCAN_IN); 
assign U6466 = ~(U6351 & REIP_REG_14__SCAN_IN); 
assign U6470 = ~(U2373 & PHYADDRPOINTER_REG_15__SCAN_IN); 
assign U6473 = ~(U6351 & REIP_REG_15__SCAN_IN); 
assign U6477 = ~(U2373 & PHYADDRPOINTER_REG_16__SCAN_IN); 
assign U6480 = ~(U6351 & REIP_REG_16__SCAN_IN); 
assign U6484 = ~(U2373 & PHYADDRPOINTER_REG_17__SCAN_IN); 
assign U6487 = ~(U6351 & REIP_REG_17__SCAN_IN); 
assign U6491 = ~(U2373 & PHYADDRPOINTER_REG_18__SCAN_IN); 
assign U6494 = ~(U6351 & REIP_REG_18__SCAN_IN); 
assign U6498 = ~(U2373 & PHYADDRPOINTER_REG_19__SCAN_IN); 
assign U6501 = ~(U6351 & REIP_REG_19__SCAN_IN); 
assign U6505 = ~(U2373 & PHYADDRPOINTER_REG_20__SCAN_IN); 
assign U6508 = ~(U6351 & REIP_REG_20__SCAN_IN); 
assign U6512 = ~(U2373 & PHYADDRPOINTER_REG_21__SCAN_IN); 
assign U6515 = ~(U6351 & REIP_REG_21__SCAN_IN); 
assign U6519 = ~(U2373 & PHYADDRPOINTER_REG_22__SCAN_IN); 
assign U6522 = ~(U6351 & REIP_REG_22__SCAN_IN); 
assign U6526 = ~(U2373 & PHYADDRPOINTER_REG_23__SCAN_IN); 
assign U6529 = ~(U6351 & REIP_REG_23__SCAN_IN); 
assign U6533 = ~(U2373 & PHYADDRPOINTER_REG_24__SCAN_IN); 
assign U6536 = ~(U6351 & REIP_REG_24__SCAN_IN); 
assign U6540 = ~(U2373 & PHYADDRPOINTER_REG_25__SCAN_IN); 
assign U6543 = ~(U6351 & REIP_REG_25__SCAN_IN); 
assign U6547 = ~(U2373 & PHYADDRPOINTER_REG_26__SCAN_IN); 
assign U6550 = ~(U6351 & REIP_REG_26__SCAN_IN); 
assign U6554 = ~(U2373 & PHYADDRPOINTER_REG_27__SCAN_IN); 
assign U6557 = ~(U6351 & REIP_REG_27__SCAN_IN); 
assign U6561 = ~(U2373 & PHYADDRPOINTER_REG_28__SCAN_IN); 
assign U6564 = ~(U6351 & REIP_REG_28__SCAN_IN); 
assign U6568 = ~(U2373 & PHYADDRPOINTER_REG_29__SCAN_IN); 
assign U6571 = ~(U6351 & REIP_REG_29__SCAN_IN); 
assign U6575 = ~(U2373 & PHYADDRPOINTER_REG_30__SCAN_IN); 
assign U6578 = ~(U6351 & REIP_REG_30__SCAN_IN); 
assign U6582 = ~(U2373 & PHYADDRPOINTER_REG_31__SCAN_IN); 
assign U6585 = ~(U6351 & REIP_REG_31__SCAN_IN); 
assign U6762 = ~(R2337_U59 & U2352); 
assign U6874 = ~(U4147 & R2144_U50); 
assign U7754 = ~(U6591 & REQUESTPENDING_REG_SCAN_IN); 
assign U7760 = ~(U6602 & READREQUEST_REG_SCAN_IN); 
assign R2027_U156 = ~(R2027_U129 & R2027_U98); 
assign R2278_U17 = R2278_U292 & R2278_U19; 
assign R2278_U161 = ~R2278_U19; 
assign R2358_U29 = ~U2650; 
assign R2358_U236 = ~(U2650 & R2358_U474); 
assign R2358_U554 = ~(U2352 & R2358_U196); 
assign R2358_U590 = ~(U2352 & R2358_U196); 
assign R2337_U149 = ~(R2337_U133 & R2337_U95); 
assign R2144_U83 = ~(R2144_U56 & R2144_U158); 
assign R2144_U84 = ~(R2144_U111 & R2144_U118); 
assign R2144_U135 = ~(R2144_U134 & R2144_U116); 
assign R2144_U138 = ~(R2144_U134 & R2144_U116 & R2144_U137); 
assign R2144_U160 = ~(R2144_U58 & R2144_U158); 
assign R2144_U239 = ~(R2144_U48 & R2144_U133); 
assign R2099_U14 = ~(R2099_U95 & R2099_U167); 
assign R2099_U141 = ~(R2099_U167 & R2099_U56); 
assign R2099_U331 = ~(R2099_U279 & R2099_U167); 
assign R2099_U333 = ~(R2099_U166 & R2099_U276); 
assign R2096_U38 = ~(R2096_U109 & REIP_REG_18__SCAN_IN); 
assign R2096_U166 = ~(R2096_U109 & R2096_U37); 
assign LT_563_U13 = LT_563_U21 & LT_563_U22; 
assign LT_563_U17 = ~(LT_563_U16 & LT_563_U15 & INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign LT_563_U18 = ~(LT_563_U15 & INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign LT_563_U19 = ~(LT_563_U8 & INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign LT_563_U24 = ~(LT_563_U9 & INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign LT_563_U25 = ~(LT_563_U12 & INSTQUEUEWR_ADDR_REG_4__SCAN_IN); 
assign LT_563_U28 = ~(LT_563_U16 & INSTQUEUEWR_ADDR_REG_1__SCAN_IN & INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign ADD_405_U38 = ~(ADD_405_U112 & INSTADDRPOINTER_REG_18__SCAN_IN); 
assign ADD_405_U170 = ~(ADD_405_U112 & ADD_405_U37); 
assign ADD_515_U38 = ~(ADD_515_U109 & INSTADDRPOINTER_REG_18__SCAN_IN); 
assign ADD_515_U166 = ~(ADD_515_U109 & ADD_515_U37); 
assign U2369 = U2362 & U4485; 
assign U2374 = U2360 & U4202; 
assign U2375 = U2360 & U4204; 
assign U2378 = U2360 & U5557; 
assign U2379 = U2363 & U3267; 
assign U2380 = U2360 & U7596; 
assign U2786 = ~(U4016 & U6875 & U6874); 
assign U3318 = ~(R2144_U43 & U3297); 
assign U3472 = ~(U7755 & U7754); 
assign U3474 = ~(U7761 & U7760); 
assign U3741 = U5540 & U5541; 
assign U3997 = U6760 & U6761 & U6762; 
assign U4217 = ~(U2362 & U3259); 
assign U4218 = ~(U2363 & U4365); 
assign U4512 = ~U3312; 
assign U4516 = ~U3300; 
assign U5560 = ~(R2278_U17 & U2377); 
assign U5563 = ~(U2370 & REIP_REG_0__SCAN_IN); 
assign U5564 = ~(U5552 & INSTADDRPOINTER_REG_0__SCAN_IN); 
assign U5570 = ~(U2370 & REIP_REG_1__SCAN_IN); 
assign U5571 = ~(U5552 & INSTADDRPOINTER_REG_1__SCAN_IN); 
assign U5577 = ~(U2370 & REIP_REG_2__SCAN_IN); 
assign U5578 = ~(U5552 & INSTADDRPOINTER_REG_2__SCAN_IN); 
assign U5584 = ~(U2370 & REIP_REG_3__SCAN_IN); 
assign U5585 = ~(U5552 & INSTADDRPOINTER_REG_3__SCAN_IN); 
assign U5591 = ~(U2370 & REIP_REG_4__SCAN_IN); 
assign U5592 = ~(U5552 & INSTADDRPOINTER_REG_4__SCAN_IN); 
assign U5598 = ~(U2370 & REIP_REG_5__SCAN_IN); 
assign U5599 = ~(U5552 & INSTADDRPOINTER_REG_5__SCAN_IN); 
assign U5605 = ~(U2370 & REIP_REG_6__SCAN_IN); 
assign U5606 = ~(U5552 & INSTADDRPOINTER_REG_6__SCAN_IN); 
assign U5612 = ~(U2370 & REIP_REG_7__SCAN_IN); 
assign U5613 = ~(U5552 & INSTADDRPOINTER_REG_7__SCAN_IN); 
assign U5619 = ~(U2370 & REIP_REG_8__SCAN_IN); 
assign U5620 = ~(U5552 & INSTADDRPOINTER_REG_8__SCAN_IN); 
assign U5626 = ~(U2370 & REIP_REG_9__SCAN_IN); 
assign U5627 = ~(U5552 & INSTADDRPOINTER_REG_9__SCAN_IN); 
assign U5633 = ~(U2370 & REIP_REG_10__SCAN_IN); 
assign U5634 = ~(U5552 & INSTADDRPOINTER_REG_10__SCAN_IN); 
assign U5640 = ~(U2370 & REIP_REG_11__SCAN_IN); 
assign U5641 = ~(U5552 & INSTADDRPOINTER_REG_11__SCAN_IN); 
assign U5647 = ~(U2370 & REIP_REG_12__SCAN_IN); 
assign U5648 = ~(U5552 & INSTADDRPOINTER_REG_12__SCAN_IN); 
assign U5654 = ~(U2370 & REIP_REG_13__SCAN_IN); 
assign U5655 = ~(U5552 & INSTADDRPOINTER_REG_13__SCAN_IN); 
assign U5661 = ~(U2370 & REIP_REG_14__SCAN_IN); 
assign U5662 = ~(U5552 & INSTADDRPOINTER_REG_14__SCAN_IN); 
assign U5668 = ~(U2370 & REIP_REG_15__SCAN_IN); 
assign U5669 = ~(U5552 & INSTADDRPOINTER_REG_15__SCAN_IN); 
assign U5675 = ~(U2370 & REIP_REG_16__SCAN_IN); 
assign U5676 = ~(U5552 & INSTADDRPOINTER_REG_16__SCAN_IN); 
assign U5682 = ~(U2370 & REIP_REG_17__SCAN_IN); 
assign U5683 = ~(U5552 & INSTADDRPOINTER_REG_17__SCAN_IN); 
assign U5689 = ~(U2370 & REIP_REG_18__SCAN_IN); 
assign U5690 = ~(U5552 & INSTADDRPOINTER_REG_18__SCAN_IN); 
assign U5696 = ~(U2370 & REIP_REG_19__SCAN_IN); 
assign U5697 = ~(U5552 & INSTADDRPOINTER_REG_19__SCAN_IN); 
assign U5703 = ~(U2370 & REIP_REG_20__SCAN_IN); 
assign U5704 = ~(U5552 & INSTADDRPOINTER_REG_20__SCAN_IN); 
assign U5710 = ~(U2370 & REIP_REG_21__SCAN_IN); 
assign U5711 = ~(U5552 & INSTADDRPOINTER_REG_21__SCAN_IN); 
assign U5717 = ~(U2370 & REIP_REG_22__SCAN_IN); 
assign U5718 = ~(U5552 & INSTADDRPOINTER_REG_22__SCAN_IN); 
assign U5724 = ~(U2370 & REIP_REG_23__SCAN_IN); 
assign U5725 = ~(U5552 & INSTADDRPOINTER_REG_23__SCAN_IN); 
assign U5731 = ~(U2370 & REIP_REG_24__SCAN_IN); 
assign U5732 = ~(U5552 & INSTADDRPOINTER_REG_24__SCAN_IN); 
assign U5738 = ~(U2370 & REIP_REG_25__SCAN_IN); 
assign U5739 = ~(U5552 & INSTADDRPOINTER_REG_25__SCAN_IN); 
assign U5745 = ~(U2370 & REIP_REG_26__SCAN_IN); 
assign U5746 = ~(U5552 & INSTADDRPOINTER_REG_26__SCAN_IN); 
assign U5752 = ~(U2370 & REIP_REG_27__SCAN_IN); 
assign U5753 = ~(U5552 & INSTADDRPOINTER_REG_27__SCAN_IN); 
assign U5759 = ~(U2370 & REIP_REG_28__SCAN_IN); 
assign U5760 = ~(U5552 & INSTADDRPOINTER_REG_28__SCAN_IN); 
assign U5766 = ~(U2370 & REIP_REG_29__SCAN_IN); 
assign U5767 = ~(U5552 & INSTADDRPOINTER_REG_29__SCAN_IN); 
assign U5773 = ~(U2370 & REIP_REG_30__SCAN_IN); 
assign U5774 = ~(U5552 & INSTADDRPOINTER_REG_30__SCAN_IN); 
assign U5780 = ~(U2370 & REIP_REG_31__SCAN_IN); 
assign U5781 = ~(U5552 & INSTADDRPOINTER_REG_31__SCAN_IN); 
assign U5788 = ~(U2372 & R2278_U17); 
assign R2027_U58 = ~(R2027_U156 & R2027_U155); 
assign R2358_U27 = ~U2649; 
assign R2358_U201 = ~U2653; 
assign R2358_U233 = ~(U2649 & R2358_U471); 
assign R2358_U235 = ~(R2358_U478 & R2358_U477 & R2358_U29); 
assign R2358_U237 = ~(R2358_U236 & R2358_U22); 
assign R2358_U565 = ~(U2653 & R2358_U22); 
assign R2358_U592 = ~(R2358_U591 & R2358_U590); 
assign R2358_U594 = ~(U2653 & R2358_U22); 
assign R2337_U58 = ~(R2337_U149 & R2337_U148); 
assign R2144_U49 = ~(R2144_U239 & R2144_U238); 
assign R2144_U99 = ~(R2144_U53 & R2144_U84); 
assign R2144_U119 = ~R2144_U84; 
assign R2144_U123 = ~R2144_U83; 
assign R2144_U124 = ~(R2144_U83 & R2144_U105); 
assign R2144_U136 = ~(R2144_U62 & R2144_U135); 
assign R2144_U215 = ~(R2144_U59 & R2144_U160 & R2144_U81); 
assign R2144_U216 = ~(R2144_U149 & R2144_U83); 
assign R2144_U218 = ~(R2144_U150 & R2144_U84); 
assign R584_U6 = ~U2676; 
assign R584_U7 = ~U2677; 
assign R584_U8 = ~U2674; 
assign R584_U9 = ~U2675; 
assign R2099_U79 = ~(R2099_U332 & R2099_U331); 
assign R2099_U80 = ~(R2099_U334 & R2099_U333); 
assign R2099_U168 = ~R2099_U141; 
assign R2099_U169 = ~R2099_U14; 
assign R2099_U328 = ~(R2099_U55 & R2099_U14); 
assign R2099_U330 = ~(R2099_U57 & R2099_U141); 
assign LT_563_1260_U7 = ~U2673; 
assign R2096_U83 = ~(R2096_U166 & R2096_U165); 
assign R2096_U110 = ~R2096_U38; 
assign R2096_U163 = ~(R2096_U38 & REIP_REG_19__SCAN_IN); 
assign LT_563_U14 = LT_563_U24 & LT_563_U25; 
assign LT_563_U20 = ~(LT_563_U28 & LT_563_U19 & LT_563_U18 & LT_563_U17); 
assign ADD_405_U83 = ~(ADD_405_U170 & ADD_405_U169); 
assign ADD_405_U113 = ~ADD_405_U38; 
assign ADD_405_U167 = ~(ADD_405_U38 & INSTADDRPOINTER_REG_19__SCAN_IN); 
assign ADD_515_U83 = ~(ADD_515_U166 & ADD_515_U165); 
assign ADD_515_U110 = ~ADD_515_U38; 
assign ADD_515_U163 = ~(ADD_515_U38 & INSTADDRPOINTER_REG_19__SCAN_IN); 
assign U2367 = U3418 & R2337_U58 & STATE2_REG_1__SCAN_IN; 
assign U2604 = U2379 & EBX_REG_31__SCAN_IN; 
assign U2652 = ~(U6759 & U3997); 
assign U3298 = ~R2144_U49; 
assign U3319 = ~(U3312 & U3318); 
assign U3417 = ~R2337_U58; 
assign U3753 = U5563 & U5564; 
assign U3757 = U5570 & U5571; 
assign U3761 = U5577 & U5578; 
assign U3765 = U5584 & U5585; 
assign U3767 = U5591 & U5592; 
assign U3770 = U5598 & U5599; 
assign U3773 = U5605 & U5606; 
assign U3776 = U5612 & U5613; 
assign U3779 = U5619 & U5620; 
assign U3782 = U5626 & U5627; 
assign U3785 = U5633 & U5634; 
assign U3788 = U5640 & U5641; 
assign U3791 = U5647 & U5648; 
assign U3794 = U5654 & U5655; 
assign U3797 = U5661 & U5662; 
assign U3800 = U5668 & U5669; 
assign U3803 = U5675 & U5676; 
assign U3806 = U5682 & U5683; 
assign U3809 = U5689 & U5690; 
assign U3812 = U5696 & U5697; 
assign U3815 = U5703 & U5704; 
assign U3818 = U5710 & U5711; 
assign U3821 = U5717 & U5718; 
assign U3824 = U5724 & U5725; 
assign U3827 = U5731 & U5732; 
assign U3830 = U5738 & U5739; 
assign U3833 = U5745 & U5746; 
assign U3836 = U5752 & U5753; 
assign U3839 = U5759 & U5760; 
assign U3842 = U5766 & U5767; 
assign U3845 = U5773 & U5774; 
assign U3848 = U5780 & U5781; 
assign U4513 = ~U3318; 
assign U5536 = ~(U4214 & R2144_U49); 
assign U5558 = ~(R2099_U86 & U2380); 
assign U5559 = ~(R2027_U5 & U2378); 
assign U5561 = ~(ADD_405_U4 & U2375); 
assign U5562 = ~(U2374 & INSTADDRPOINTER_REG_0__SCAN_IN); 
assign U5565 = ~(R2099_U87 & U2380); 
assign U5566 = ~(R2027_U71 & U2378); 
assign U5568 = ~(ADD_405_U81 & U2375); 
assign U5569 = ~(ADD_515_U4 & U2374); 
assign U5572 = ~(R2099_U138 & U2380); 
assign U5573 = ~(R2027_U60 & U2378); 
assign U5575 = ~(ADD_405_U5 & U2375); 
assign U5576 = ~(ADD_515_U71 & U2374); 
assign U5579 = ~(R2099_U42 & U2380); 
assign U5580 = ~(R2027_U57 & U2378); 
assign U5582 = ~(ADD_405_U93 & U2375); 
assign U5583 = ~(ADD_515_U68 & U2374); 
assign U5586 = ~(R2099_U41 & U2380); 
assign U5587 = ~(R2027_U56 & U2378); 
assign U5589 = ~(ADD_405_U68 & U2375); 
assign U5590 = ~(ADD_515_U67 & U2374); 
assign U5593 = ~(R2099_U40 & U2380); 
assign U5594 = ~(R2027_U55 & U2378); 
assign U5596 = ~(ADD_405_U67 & U2375); 
assign U5597 = ~(ADD_515_U66 & U2374); 
assign U5600 = ~(R2099_U39 & U2380); 
assign U5601 = ~(R2027_U54 & U2378); 
assign U5603 = ~(ADD_405_U66 & U2375); 
assign U5604 = ~(ADD_515_U65 & U2374); 
assign U5607 = ~(R2099_U38 & U2380); 
assign U5608 = ~(R2027_U53 & U2378); 
assign U5610 = ~(ADD_405_U65 & U2375); 
assign U5611 = ~(ADD_515_U64 & U2374); 
assign U5614 = ~(R2099_U37 & U2380); 
assign U5615 = ~(R2027_U52 & U2378); 
assign U5617 = ~(ADD_405_U64 & U2375); 
assign U5618 = ~(ADD_515_U63 & U2374); 
assign U5621 = ~(R2099_U36 & U2380); 
assign U5622 = ~(R2027_U51 & U2378); 
assign U5624 = ~(ADD_405_U63 & U2375); 
assign U5625 = ~(ADD_515_U62 & U2374); 
assign U5628 = ~(R2099_U85 & U2380); 
assign U5629 = ~(R2027_U81 & U2378); 
assign U5631 = ~(ADD_405_U91 & U2375); 
assign U5632 = ~(ADD_515_U91 & U2374); 
assign U5635 = ~(R2099_U84 & U2380); 
assign U5636 = ~(R2027_U80 & U2378); 
assign U5638 = ~(ADD_405_U90 & U2375); 
assign U5639 = ~(ADD_515_U90 & U2374); 
assign U5642 = ~(R2099_U83 & U2380); 
assign U5643 = ~(R2027_U79 & U2378); 
assign U5645 = ~(ADD_405_U89 & U2375); 
assign U5646 = ~(ADD_515_U89 & U2374); 
assign U5649 = ~(R2099_U82 & U2380); 
assign U5650 = ~(R2027_U78 & U2378); 
assign U5652 = ~(ADD_405_U88 & U2375); 
assign U5653 = ~(ADD_515_U88 & U2374); 
assign U5656 = ~(R2099_U81 & U2380); 
assign U5657 = ~(R2027_U77 & U2378); 
assign U5659 = ~(ADD_405_U87 & U2375); 
assign U5660 = ~(ADD_515_U87 & U2374); 
assign U5663 = ~(R2099_U80 & U2380); 
assign U5664 = ~(R2027_U76 & U2378); 
assign U5666 = ~(ADD_405_U86 & U2375); 
assign U5667 = ~(ADD_515_U86 & U2374); 
assign U5670 = ~(R2099_U79 & U2380); 
assign U5671 = ~(R2027_U75 & U2378); 
assign U5673 = ~(ADD_405_U85 & U2375); 
assign U5674 = ~(ADD_515_U85 & U2374); 
assign U5678 = ~(R2027_U74 & U2378); 
assign U5680 = ~(ADD_405_U84 & U2375); 
assign U5681 = ~(ADD_515_U84 & U2374); 
assign U5685 = ~(R2027_U73 & U2378); 
assign U5687 = ~(ADD_405_U83 & U2375); 
assign U5688 = ~(ADD_515_U83 & U2374); 
assign U5692 = ~(R2027_U72 & U2378); 
assign U5699 = ~(R2027_U70 & U2378); 
assign U5706 = ~(R2027_U69 & U2378); 
assign U5713 = ~(R2027_U68 & U2378); 
assign U5720 = ~(R2027_U67 & U2378); 
assign U5727 = ~(R2027_U66 & U2378); 
assign U5734 = ~(R2027_U65 & U2378); 
assign U5741 = ~(R2027_U64 & U2378); 
assign U5748 = ~(R2027_U63 & U2378); 
assign U5755 = ~(R2027_U62 & U2378); 
assign U5762 = ~(R2027_U61 & U2378); 
assign U5769 = ~(R2027_U59 & U2378); 
assign U5776 = ~(R2027_U58 & U2378); 
assign U5942 = ~(R2337_U58 & U2376); 
assign U6299 = ~(U2371 & R2099_U80); 
assign U6302 = ~(U2371 & R2099_U79); 
assign U6353 = ~(R2337_U58 & STATE2_REG_1__SCAN_IN); 
assign U6758 = ~(R2337_U58 & U2352); 
assign U6857 = ~(R2144_U49 & U6734); 
assign U6871 = ~(U4147 & R2144_U49); 
assign U7469 = ~(U2379 & U3416); 
assign U7470 = ~(U2369 & U6355); 
assign U7471 = ~(U3876 & U2369); 
assign U7679 = ~(R2144_U49 & U3300); 
assign R2278_U168 = U2786 | INSTADDRPOINTER_REG_1__SCAN_IN; 
assign R2278_U169 = ~(U2786 & INSTADDRPOINTER_REG_1__SCAN_IN); 
assign R2358_U218 = ~(R2358_U236 & R2358_U235); 
assign R2358_U232 = ~(R2358_U476 & R2358_U475 & R2358_U27); 
assign R2358_U268 = ~(U2352 & R2358_U235); 
assign R2358_U564 = ~(U2352 & R2358_U201); 
assign R2358_U593 = ~(U2352 & R2358_U201); 
assign R2144_U8 = R2144_U138 & R2144_U136; 
assign R2144_U79 = ~(R2144_U99 & R2144_U54); 
assign R2144_U82 = R2144_U215 & R2144_U214; 
assign R2144_U125 = ~(R2144_U21 & R2144_U124); 
assign R2144_U127 = ~(R2144_U60 & R2144_U124); 
assign R2144_U212 = ~(R2144_U57 & R2144_U124 & R2144_U23); 
assign R2144_U217 = ~(R2144_U44 & R2144_U123); 
assign R2144_U219 = ~(R2144_U46 & R2144_U119); 
assign LT_589_U7 = R584_U7 & R584_U6; 
assign R2099_U15 = ~(R2099_U169 & R2099_U55); 
assign R2099_U327 = ~(R2099_U258 & R2099_U169); 
assign R2099_U329 = ~(R2099_U168 & R2099_U282); 
assign LT_563_1260_U8 = ~(R584_U8 & LT_563_1260_U7); 
assign LT_563_1260_U9 = ~(R584_U9 & LT_563_1260_U7); 
assign R2096_U40 = ~(R2096_U110 & REIP_REG_19__SCAN_IN); 
assign R2096_U164 = ~(R2096_U110 & R2096_U39); 
assign LT_563_U23 = ~(LT_563_U13 & LT_563_U20); 
assign ADD_405_U40 = ~(ADD_405_U113 & INSTADDRPOINTER_REG_19__SCAN_IN); 
assign ADD_405_U168 = ~(ADD_405_U113 & ADD_405_U39); 
assign ADD_515_U40 = ~(ADD_515_U110 & INSTADDRPOINTER_REG_19__SCAN_IN); 
assign ADD_515_U164 = ~(ADD_515_U110 & ADD_515_U39); 
assign U2366 = U3418 & U3417 & STATE2_REG_1__SCAN_IN; 
assign U2476 = R2144_U8 & R2144_U49; 
assign U2508 = ~(R2144_U49 | R2144_U8); 
assign U2647 = R2144_U8 & U6734; 
assign U2648 = ~(U3427 & U6857); 
assign U2651 = ~(U6757 & U6756 & U6758); 
assign U2785 = ~(U6872 & U6873 & U6871); 
assign U3299 = ~R2144_U8; 
assign U3301 = ~(U3319 & U3296); 
assign U3313 = ~(R2144_U43 & U3319); 
assign U3329 = ~(R2144_U8 & U3298); 
assign U3740 = U5535 & U5536; 
assign U3751 = U5559 & U5558; 
assign U3752 = U5561 & U5560; 
assign U3754 = U3753 & U5562; 
assign U3755 = U5566 & U5565; 
assign U3758 = U3757 & U5569; 
assign U3759 = U5573 & U5572; 
assign U3762 = U3761 & U5576; 
assign U3763 = U5580 & U5579 & U5582; 
assign U3766 = U5587 & U5586 & U5589; 
assign U3768 = U3767 & U5590; 
assign U3769 = U5594 & U5593 & U5596; 
assign U3771 = U3770 & U5597; 
assign U3772 = U5601 & U5600 & U5603; 
assign U3774 = U3773 & U5604; 
assign U3775 = U5608 & U5607 & U5610; 
assign U3777 = U3776 & U5611; 
assign U3778 = U5615 & U5614 & U5617; 
assign U3780 = U3779 & U5618; 
assign U3781 = U5622 & U5621 & U5624; 
assign U3783 = U3782 & U5625; 
assign U3784 = U5629 & U5628 & U5631; 
assign U3786 = U3785 & U5632; 
assign U3787 = U5636 & U5635 & U5638; 
assign U3789 = U3788 & U5639; 
assign U3790 = U5643 & U5642 & U5645; 
assign U3792 = U3791 & U5646; 
assign U3793 = U5650 & U5652; 
assign U3795 = U3794 & U5653; 
assign U3796 = U5657 & U5659; 
assign U3798 = U3797 & U5660; 
assign U3799 = U5664 & U5666; 
assign U3801 = U3800 & U5667; 
assign U3802 = U5671 & U5673; 
assign U3804 = U3803 & U5674; 
assign U3805 = U5678 & U5680; 
assign U3807 = U3806 & U5681; 
assign U3808 = U5685 & U5687; 
assign U3810 = U3809 & U5688; 
assign U4514 = ~U3319; 
assign U4518 = ~(R2144_U8 & U3300); 
assign U5532 = ~(U4214 & R2144_U8); 
assign U6354 = ~(U6353 & U6352); 
assign U6356 = ~(U2604 & R2099_U86); 
assign U6364 = ~(U2604 & R2099_U87); 
assign U6372 = ~(U2604 & R2099_U138); 
assign U6380 = ~(U2604 & R2099_U42); 
assign U6388 = ~(U2604 & R2099_U41); 
assign U6396 = ~(U2604 & R2099_U40); 
assign U6404 = ~(U2604 & R2099_U39); 
assign U6411 = ~(U2604 & R2099_U38); 
assign U6418 = ~(U2604 & R2099_U37); 
assign U6425 = ~(U2604 & R2099_U36); 
assign U6432 = ~(U2604 & R2099_U85); 
assign U6439 = ~(U2604 & R2099_U84); 
assign U6446 = ~(U2604 & R2099_U83); 
assign U6453 = ~(U2604 & R2099_U82); 
assign U6460 = ~(U2604 & R2099_U81); 
assign U6467 = ~(U2604 & R2099_U80); 
assign U6474 = ~(U2604 & R2099_U79); 
assign U6869 = ~(U4147 & R2144_U8); 
assign U7472 = ~(U7469 & U4217 & U7470); 
assign U7473 = ~(U7471 & U4218); 
assign U7680 = ~(U4516 & U3298); 
assign R2278_U130 = ~(R2278_U168 & R2278_U169); 
assign R2278_U170 = ~(R2278_U161 & R2278_U168); 
assign R2358_U111 = R2358_U233 & R2358_U232; 
assign R2358_U123 = R2358_U235 & R2358_U232; 
assign R2358_U200 = ~U2652; 
assign R2358_U212 = ~(R2358_U236 & R2358_U268); 
assign R2358_U380 = ~R2358_U218; 
assign R2358_U395 = ~(R2358_U233 & R2358_U232); 
assign R2358_U563 = ~(U2652 & R2358_U22); 
assign R2358_U579 = ~(U2652 & R2358_U22); 
assign R2358_U595 = ~(R2358_U594 & R2358_U593); 
assign R2358_U653 = ~(U2352 & R2358_U218); 
assign R2144_U10 = R2144_U213 & R2144_U212 & R2144_U82; 
assign R2144_U24 = ~(R2144_U79 & R2144_U63); 
assign R2144_U25 = ~(R2144_U6 & R2144_U79); 
assign R2144_U45 = ~(R2144_U217 & R2144_U216); 
assign R2144_U47 = ~(R2144_U219 & R2144_U218); 
assign R2144_U78 = ~(R2144_U29 & R2144_U79); 
assign R2144_U96 = ~(R2144_U79 & R2144_U66); 
assign R2144_U97 = ~(R2144_U67 & R2144_U79); 
assign R2144_U121 = ~R2144_U79; 
assign R2144_U128 = ~(R2144_U61 & R2144_U125); 
assign R2144_U211 = ~(R2144_U29 & R2144_U79); 
assign LT_589_U8 = ~(LT_589_U7 | R584_U9 | R584_U8); 
assign R2099_U77 = ~(R2099_U328 & R2099_U327); 
assign R2099_U78 = ~(R2099_U330 & R2099_U329); 
assign R2099_U170 = ~R2099_U15; 
assign R2099_U326 = ~(R2099_U54 & R2099_U15); 
assign LT_563_1260_U6 = LT_563_1260_U9 & LT_563_1260_U8; 
assign R2096_U82 = ~(R2096_U164 & R2096_U163); 
assign R2096_U111 = ~R2096_U40; 
assign R2096_U161 = ~(R2096_U40 & REIP_REG_20__SCAN_IN); 
assign LT_563_U26 = ~(LT_563_U14 & LT_563_U23); 
assign ADD_405_U82 = ~(ADD_405_U168 & ADD_405_U167); 
assign ADD_405_U114 = ~ADD_405_U40; 
assign ADD_405_U163 = ~(ADD_405_U40 & INSTADDRPOINTER_REG_20__SCAN_IN); 
assign ADD_515_U82 = ~(ADD_515_U164 & ADD_515_U163); 
assign ADD_515_U111 = ~ADD_515_U40; 
assign ADD_515_U161 = ~(ADD_515_U40 & INSTADDRPOINTER_REG_20__SCAN_IN); 
assign U2429 = U6354 & U3418; 
assign U2474 = R2144_U49 & U3299; 
assign U2477 = U4516 & U2476; 
assign U2481 = U4512 & U2476; 
assign U2483 = U4513 & U2476; 
assign U2485 = U4514 & R2144_U43; 
assign U2487 = U2486 & U2476; 
assign U2509 = U2508 & U4516; 
assign U2512 = U2508 & U4512; 
assign U2514 = U2508 & U4513; 
assign U2516 = U2508 & U2486; 
assign U2643 = R2144_U10 & U6734; 
assign U2645 = R2144_U45 & U6734; 
assign U2646 = R2144_U47 & U6734; 
assign U2784 = ~(U6870 & U6869); 
assign U3018 = ~(U3752 & U3751 & U3754); 
assign U3320 = ~(U4514 & U3296); 
assign U3441 = ~(U7680 & U7679); 
assign U3739 = U5531 & U5532; 
assign U3882 = U6388 & U4215; 
assign U3884 = U6396 & U4215; 
assign U3886 = U6404 & U4215; 
assign U3888 = U6411 & U4215; 
assign U3890 = U6418 & U4215; 
assign U3892 = U6425 & U4215; 
assign U3894 = U6432 & U4215; 
assign U3896 = U6439 & U4215; 
assign U3898 = U6446 & U4215; 
assign U3900 = U6453 & U4215; 
assign U3902 = U6460 & U4215; 
assign U3904 = U6467 & U4215; 
assign U3906 = U6474 & U4215; 
assign U4213 = ~LT_563_1260_U6; 
assign U4515 = ~U3301; 
assign U4517 = ~U3329; 
assign U4536 = ~(U4516 & U2476); 
assign U4588 = ~U3313; 
assign U4594 = ~(U4512 & U2476); 
assign U4653 = ~(U4513 & U2476); 
assign U4710 = ~(U2486 & U2476); 
assign U5226 = ~(U2508 & U4516); 
assign U5283 = ~(U2508 & U4512); 
assign U5341 = ~(U2508 & U4513); 
assign U5398 = ~(U2508 & U2486); 
assign U5677 = ~(R2099_U78 & U2380); 
assign U5684 = ~(R2099_U77 & U2380); 
assign U5694 = ~(ADD_405_U82 & U2375); 
assign U5695 = ~(ADD_515_U82 & U2374); 
assign U6305 = ~(U2371 & R2099_U78); 
assign U6308 = ~(U2371 & R2099_U77); 
assign U6357 = ~(U7473 & REIP_REG_0__SCAN_IN); 
assign U6358 = ~(U7472 & EBX_REG_0__SCAN_IN); 
assign U6362 = ~(U2366 & PHYADDRPOINTER_REG_0__SCAN_IN); 
assign U6365 = ~(R2096_U4 & U7473); 
assign U6366 = ~(U7472 & EBX_REG_1__SCAN_IN); 
assign U6370 = ~(U2366 & R2337_U5); 
assign U6373 = ~(R2096_U71 & U7473); 
assign U6374 = ~(U7472 & EBX_REG_2__SCAN_IN); 
assign U6378 = ~(U2366 & R2337_U60); 
assign U6381 = ~(R2096_U68 & U7473); 
assign U6382 = ~(U7472 & EBX_REG_3__SCAN_IN); 
assign U6386 = ~(U2366 & R2337_U57); 
assign U6389 = ~(R2096_U67 & U7473); 
assign U6390 = ~(U7472 & EBX_REG_4__SCAN_IN); 
assign U6394 = ~(U2366 & R2337_U56); 
assign U6397 = ~(R2096_U66 & U7473); 
assign U6398 = ~(U7472 & EBX_REG_5__SCAN_IN); 
assign U6402 = ~(U2366 & R2337_U55); 
assign U6405 = ~(R2096_U65 & U7473); 
assign U6406 = ~(U7472 & EBX_REG_6__SCAN_IN); 
assign U6409 = ~(U2366 & R2337_U54); 
assign U6412 = ~(R2096_U64 & U7473); 
assign U6413 = ~(U7472 & EBX_REG_7__SCAN_IN); 
assign U6416 = ~(U2366 & R2337_U53); 
assign U6419 = ~(R2096_U63 & U7473); 
assign U6420 = ~(U7472 & EBX_REG_8__SCAN_IN); 
assign U6423 = ~(U2366 & R2337_U52); 
assign U6426 = ~(R2096_U62 & U7473); 
assign U6427 = ~(U7472 & EBX_REG_9__SCAN_IN); 
assign U6430 = ~(U2366 & R2337_U51); 
assign U6433 = ~(R2096_U91 & U7473); 
assign U6434 = ~(U7472 & EBX_REG_10__SCAN_IN); 
assign U6437 = ~(U2366 & R2337_U80); 
assign U6440 = ~(R2096_U90 & U7473); 
assign U6441 = ~(U7472 & EBX_REG_11__SCAN_IN); 
assign U6444 = ~(U2366 & R2337_U79); 
assign U6447 = ~(R2096_U89 & U7473); 
assign U6448 = ~(U7472 & EBX_REG_12__SCAN_IN); 
assign U6451 = ~(U2366 & R2337_U78); 
assign U6454 = ~(R2096_U88 & U7473); 
assign U6455 = ~(U7472 & EBX_REG_13__SCAN_IN); 
assign U6458 = ~(U2366 & R2337_U77); 
assign U6461 = ~(R2096_U87 & U7473); 
assign U6462 = ~(U7472 & EBX_REG_14__SCAN_IN); 
assign U6465 = ~(U2366 & R2337_U76); 
assign U6468 = ~(R2096_U86 & U7473); 
assign U6469 = ~(U7472 & EBX_REG_15__SCAN_IN); 
assign U6472 = ~(U2366 & R2337_U75); 
assign U6475 = ~(R2096_U85 & U7473); 
assign U6476 = ~(U7472 & EBX_REG_16__SCAN_IN); 
assign U6479 = ~(U2366 & R2337_U74); 
assign U6481 = ~(U2604 & R2099_U78); 
assign U6482 = ~(R2096_U84 & U7473); 
assign U6483 = ~(U7472 & EBX_REG_17__SCAN_IN); 
assign U6486 = ~(U2366 & R2337_U73); 
assign U6488 = ~(U2604 & R2099_U77); 
assign U6489 = ~(R2096_U83 & U7473); 
assign U6490 = ~(U7472 & EBX_REG_18__SCAN_IN); 
assign U6493 = ~(U2366 & R2337_U72); 
assign U6496 = ~(R2096_U82 & U7473); 
assign U6497 = ~(U7472 & EBX_REG_19__SCAN_IN); 
assign U6500 = ~(U2366 & R2337_U71); 
assign U6504 = ~(U7472 & EBX_REG_20__SCAN_IN); 
assign U6507 = ~(U2366 & R2337_U70); 
assign U6511 = ~(U7472 & EBX_REG_21__SCAN_IN); 
assign U6514 = ~(U2366 & R2337_U69); 
assign U6518 = ~(U7472 & EBX_REG_22__SCAN_IN); 
assign U6521 = ~(U2366 & R2337_U68); 
assign U6525 = ~(U7472 & EBX_REG_23__SCAN_IN); 
assign U6528 = ~(U2366 & R2337_U67); 
assign U6532 = ~(U7472 & EBX_REG_24__SCAN_IN); 
assign U6535 = ~(U2366 & R2337_U66); 
assign U6539 = ~(U7472 & EBX_REG_25__SCAN_IN); 
assign U6542 = ~(U2366 & R2337_U65); 
assign U6546 = ~(U7472 & EBX_REG_26__SCAN_IN); 
assign U6549 = ~(U2366 & R2337_U64); 
assign U6553 = ~(U7472 & EBX_REG_27__SCAN_IN); 
assign U6556 = ~(U2366 & R2337_U63); 
assign U6560 = ~(U7472 & EBX_REG_28__SCAN_IN); 
assign U6563 = ~(U2366 & R2337_U62); 
assign U6567 = ~(U7472 & EBX_REG_29__SCAN_IN); 
assign U6570 = ~(U2366 & R2337_U61); 
assign U6574 = ~(U7472 & EBX_REG_30__SCAN_IN); 
assign U6577 = ~(U2366 & R2337_U59); 
assign U6581 = ~(U7472 & EBX_REG_31__SCAN_IN); 
assign U6584 = ~(U2366 & R2337_U58); 
assign U6861 = ~(U4147 & R2144_U10); 
assign U6865 = ~(U4147 & R2144_U45); 
assign U6867 = ~(U4147 & R2144_U47); 
assign R2278_U99 = ~(R2278_U169 & R2278_U170); 
assign R2278_U167 = U2785 | INSTADDRPOINTER_REG_2__SCAN_IN; 
assign R2278_U172 = ~(U2785 & INSTADDRPOINTER_REG_2__SCAN_IN); 
assign R2278_U271 = ~R2278_U130; 
assign R2278_U299 = U2785 | INSTADDRPOINTER_REG_2__SCAN_IN; 
assign R2278_U401 = ~(R2278_U161 & R2278_U130); 
assign R2358_U28 = ~U2648; 
assign R2358_U30 = ~U2647; 
assign R2358_U179 = ~U2651; 
assign R2358_U230 = ~(U2647 & R2358_U485); 
assign R2358_U234 = ~(U2648 & R2358_U468); 
assign R2358_U238 = ~(R2358_U123 & R2358_U237); 
assign R2358_U269 = ~R2358_U212; 
assign R2358_U270 = ~(R2358_U212 & R2358_U232); 
assign R2358_U505 = ~(U2651 & R2358_U22); 
assign R2358_U507 = ~(U2651 & R2358_U22); 
assign R2358_U562 = ~(U2352 & R2358_U200); 
assign R2358_U578 = ~(U2352 & R2358_U200); 
assign R2358_U633 = ~(R2358_U395 & R2358_U212); 
assign R2358_U654 = ~(R2358_U380 & R2358_U22); 
assign R2144_U9 = R2144_U128 & R2144_U127; 
assign R2144_U101 = ~R2144_U24; 
assign R2144_U122 = ~R2144_U78; 
assign R2144_U139 = ~R2144_U97; 
assign R2144_U140 = ~R2144_U96; 
assign R2144_U141 = ~R2144_U25; 
assign R2144_U144 = ~(U2355 & R2144_U24); 
assign R2144_U209 = ~(R2144_U27 & R2144_U78); 
assign R2144_U210 = ~(R2144_U121 & R2144_U204); 
assign R2144_U254 = ~(R2144_U34 & R2144_U25); 
assign R2144_U256 = ~(R2144_U35 & R2144_U96); 
assign R2144_U258 = ~(R2144_U36 & R2144_U97); 
assign LT_589_U6 = LT_589_U8 | U2673; 
assign R2099_U16 = ~(R2099_U170 & R2099_U54); 
assign R2099_U325 = ~(R2099_U255 & R2099_U170); 
assign R2096_U42 = ~(R2096_U111 & REIP_REG_20__SCAN_IN); 
assign R2096_U162 = ~(R2096_U111 & R2096_U41); 
assign LT_563_U6 = LT_563_U27 & LT_563_U26; 
assign ADD_405_U42 = ~(ADD_405_U114 & INSTADDRPOINTER_REG_20__SCAN_IN); 
assign ADD_405_U164 = ~(ADD_405_U114 & ADD_405_U41); 
assign ADD_515_U42 = ~(ADD_515_U111 & INSTADDRPOINTER_REG_20__SCAN_IN); 
assign ADD_515_U162 = ~(ADD_515_U111 & ADD_515_U41); 
assign U2491 = U4517 & U4516; 
assign U2493 = U4517 & U4512; 
assign U2495 = U4517 & U4513; 
assign U2497 = U4517 & U2486; 
assign U2501 = U4512 & U2474; 
assign U2503 = U4513 & U2474; 
assign U2505 = U2486 & U2474; 
assign U2644 = R2144_U9 & U6734; 
assign U2780 = ~(U6862 & U6861); 
assign U2782 = ~(U6866 & U6865); 
assign U2783 = ~(U6868 & U6867); 
assign U3280 = ~(U4166 & U4497 & U7614 & U4213 & LT_563_U6); 
assign U3344 = ~(U2474 & U4516); 
assign U3390 = ~LT_589_U6; 
assign U3811 = U5692 & U5694; 
assign U3813 = U3812 & U5695; 
assign U3883 = U6393 & U6392 & U6395 & U6394; 
assign U3887 = U6410 & U6407 & U6409; 
assign U3889 = U6417 & U6414 & U6416; 
assign U3891 = U6424 & U6421 & U6423; 
assign U3893 = U6431 & U6428 & U6430; 
assign U3895 = U6438 & U6435 & U6437; 
assign U3897 = U6445 & U6442 & U6444; 
assign U3899 = U6452 & U6449 & U6451; 
assign U3901 = U6459 & U6456 & U6458; 
assign U3903 = U6466 & U6463 & U6465; 
assign U3905 = U6473 & U6470 & U6472; 
assign U3907 = U6480 & U6477 & U6479; 
assign U3908 = U4215 & U6482; 
assign U3909 = U6487 & U6484 & U6486; 
assign U3910 = U4215 & U6489; 
assign U3911 = U6494 & U6491 & U6493; 
assign U3912 = U4215 & U6496; 
assign U3913 = U6501 & U6498 & U6500; 
assign U3915 = U6507 & U6508; 
assign U3917 = U6514 & U6515; 
assign U3919 = U6521 & U6522; 
assign U3921 = U6528 & U6529; 
assign U3923 = U6535 & U6536; 
assign U3925 = U6542 & U6543; 
assign U3927 = U6549 & U6550; 
assign U3929 = U6556 & U6557; 
assign U3931 = U6563 & U6564; 
assign U3933 = U6570 & U6571; 
assign U3935 = U6577 & U6578; 
assign U3937 = U6584 & U6585; 
assign U4549 = ~(U2413 & U2477); 
assign U4554 = ~(U2411 & U2477); 
assign U4559 = ~(U2409 & U2477); 
assign U4564 = ~(U2407 & U2477); 
assign U4569 = ~(U2405 & U2477); 
assign U4574 = ~(U2403 & U2477); 
assign U4579 = ~(U2401 & U2477); 
assign U4584 = ~(U2399 & U2477); 
assign U4607 = ~(U2481 & U2413); 
assign U4612 = ~(U2481 & U2411); 
assign U4617 = ~(U2481 & U2409); 
assign U4622 = ~(U2481 & U2407); 
assign U4627 = ~(U2481 & U2405); 
assign U4632 = ~(U2481 & U2403); 
assign U4637 = ~(U2481 & U2401); 
assign U4642 = ~(U2481 & U2399); 
assign U4646 = ~U3320; 
assign U4666 = ~(U2483 & U2413); 
assign U4671 = ~(U2483 & U2411); 
assign U4676 = ~(U2483 & U2409); 
assign U4681 = ~(U2483 & U2407); 
assign U4686 = ~(U2483 & U2405); 
assign U4691 = ~(U2483 & U2403); 
assign U4696 = ~(U2483 & U2401); 
assign U4701 = ~(U2483 & U2399); 
assign U4723 = ~(U2487 & U2413); 
assign U4728 = ~(U2487 & U2411); 
assign U4733 = ~(U2487 & U2409); 
assign U4738 = ~(U2487 & U2407); 
assign U4743 = ~(U2487 & U2405); 
assign U4748 = ~(U2487 & U2403); 
assign U4753 = ~(U2487 & U2401); 
assign U4758 = ~(U2487 & U2399); 
assign U4768 = ~(U4517 & U4516); 
assign U4825 = ~(U4517 & U4512); 
assign U4883 = ~(U4517 & U4513); 
assign U4940 = ~(U4517 & U2486); 
assign U5053 = ~(U4512 & U2474); 
assign U5111 = ~(U4513 & U2474); 
assign U5168 = ~(U2486 & U2474); 
assign U5239 = ~(U2509 & U2413); 
assign U5244 = ~(U2509 & U2411); 
assign U5249 = ~(U2509 & U2409); 
assign U5254 = ~(U2509 & U2407); 
assign U5259 = ~(U2509 & U2405); 
assign U5264 = ~(U2509 & U2403); 
assign U5269 = ~(U2509 & U2401); 
assign U5274 = ~(U2509 & U2399); 
assign U5296 = ~(U2512 & U2413); 
assign U5301 = ~(U2512 & U2411); 
assign U5306 = ~(U2512 & U2409); 
assign U5311 = ~(U2512 & U2407); 
assign U5316 = ~(U2512 & U2405); 
assign U5321 = ~(U2512 & U2403); 
assign U5326 = ~(U2512 & U2401); 
assign U5331 = ~(U2512 & U2399); 
assign U5354 = ~(U2514 & U2413); 
assign U5359 = ~(U2514 & U2411); 
assign U5364 = ~(U2514 & U2409); 
assign U5369 = ~(U2514 & U2407); 
assign U5374 = ~(U2514 & U2405); 
assign U5379 = ~(U2514 & U2403); 
assign U5384 = ~(U2514 & U2401); 
assign U5389 = ~(U2514 & U2399); 
assign U5411 = ~(U2516 & U2413); 
assign U5416 = ~(U2516 & U2411); 
assign U5421 = ~(U2516 & U2409); 
assign U5426 = ~(U2516 & U2407); 
assign U5430 = ~(U2516 & U2405); 
assign U5435 = ~(U2516 & U2403); 
assign U5440 = ~(U2516 & U2401); 
assign U5445 = ~(U2516 & U2399); 
assign U5524 = ~(U2428 & LT_589_U6 & STATE2_REG_0__SCAN_IN); 
assign U5527 = ~(U4515 & U3441); 
assign U5538 = ~(U3313 & U3320); 
assign U6863 = ~(U4147 & R2144_U9); 
assign U7681 = ~U3441; 
assign U7720 = ~(U3441 & U3301); 
assign R2278_U100 = ~(R2278_U167 & R2278_U172); 
assign R2278_U166 = U2784 | INSTADDRPOINTER_REG_3__SCAN_IN; 
assign R2278_U171 = ~R2278_U99; 
assign R2278_U173 = ~(R2278_U99 & R2278_U299); 
assign R2278_U175 = ~(U2784 & INSTADDRPOINTER_REG_3__SCAN_IN); 
assign R2278_U402 = ~(R2278_U271 & R2278_U19); 
assign R2358_U23 = ~U2643; 
assign R2358_U25 = ~U2645; 
assign R2358_U26 = ~U2646; 
assign R2358_U64 = ~(R2358_U233 & R2358_U270); 
assign R2358_U82 = ~(R2358_U654 & R2358_U653); 
assign R2358_U229 = ~(R2358_U480 & R2358_U479 & R2358_U28); 
assign R2358_U231 = ~(R2358_U482 & R2358_U481 & R2358_U30); 
assign R2358_U239 = ~(R2358_U238 & R2358_U233 & R2358_U234); 
assign R2358_U245 = ~(U2643 & R2358_U450); 
assign R2358_U246 = ~(U2645 & R2358_U458); 
assign R2358_U247 = ~(U2646 & R2358_U461); 
assign R2358_U504 = ~(U2352 & R2358_U179); 
assign R2358_U506 = ~(U2352 & R2358_U179); 
assign R2358_U580 = ~(R2358_U579 & R2358_U578); 
assign R2358_U634 = ~(R2358_U111 & R2358_U269); 
assign R2144_U26 = ~(R2144_U65 & R2144_U141); 
assign R2144_U80 = R2144_U211 & R2144_U210; 
assign R2144_U95 = ~(R2144_U141 & R2144_U34); 
assign R2144_U145 = ~R2144_U144; 
assign R2144_U146 = ~(R2144_U101 & R2144_U12); 
assign R2144_U208 = ~(R2144_U122 & R2144_U207); 
assign R2144_U253 = ~(R2144_U231 & R2144_U141); 
assign R2144_U255 = ~(R2144_U140 & R2144_U234); 
assign R2144_U257 = ~(R2144_U139 & R2144_U237); 
assign R2099_U76 = ~(R2099_U326 & R2099_U325); 
assign R2099_U171 = ~R2099_U16; 
assign R2099_U317 = ~(R2099_U53 & R2099_U16); 
assign R2096_U81 = ~(R2096_U162 & R2096_U161); 
assign R2096_U112 = ~R2096_U42; 
assign R2096_U159 = ~(R2096_U42 & REIP_REG_21__SCAN_IN); 
assign ADD_405_U80 = ~(ADD_405_U164 & ADD_405_U163); 
assign ADD_405_U115 = ~ADD_405_U42; 
assign ADD_405_U161 = ~(ADD_405_U42 & INSTADDRPOINTER_REG_21__SCAN_IN); 
assign ADD_515_U81 = ~(ADD_515_U162 & ADD_515_U161); 
assign ADD_515_U112 = ~ADD_515_U42; 
assign ADD_515_U159 = ~(ADD_515_U42 & INSTADDRPOINTER_REG_21__SCAN_IN); 
assign U2620 = R2144_U145 & U6734; 
assign U2621 = R2144_U145 & U6734; 
assign U2622 = R2144_U145 & U6734; 
assign U2623 = R2144_U145 & U6734; 
assign U2624 = R2144_U145 & U6734; 
assign U2625 = R2144_U145 & U6734; 
assign U2626 = R2144_U145 & U6734; 
assign U2627 = R2144_U145 & U6734; 
assign U2628 = R2144_U145 & U6734; 
assign U2629 = R2144_U145 & U6734; 
assign U2630 = R2144_U145 & U6734; 
assign U2631 = R2144_U145 & U6734; 
assign U2632 = R2144_U145 & U6734; 
assign U2633 = R2144_U145 & U6734; 
assign U2642 = R2144_U80 & U6734; 
assign U2769 = R2144_U145 & U4147; 
assign U2770 = U4147 & R2144_U145; 
assign U2781 = ~(U6864 & U6863); 
assign U3345 = ~(U3329 & U4518 & U3344); 
assign U3391 = ~(U4230 & U3287 & U5524); 
assign U4226 = ~U3344; 
assign U4233 = ~(U2428 & U3390); 
assign U4499 = ~U3280; 
assign U4511 = ~(U2368 & U3280); 
assign U4781 = ~(U2491 & U2413); 
assign U4786 = ~(U2491 & U2411); 
assign U4791 = ~(U2491 & U2409); 
assign U4796 = ~(U2491 & U2407); 
assign U4801 = ~(U2491 & U2405); 
assign U4806 = ~(U2491 & U2403); 
assign U4811 = ~(U2491 & U2401); 
assign U4816 = ~(U2491 & U2399); 
assign U4838 = ~(U2493 & U2413); 
assign U4843 = ~(U2493 & U2411); 
assign U4848 = ~(U2493 & U2409); 
assign U4853 = ~(U2493 & U2407); 
assign U4858 = ~(U2493 & U2405); 
assign U4863 = ~(U2493 & U2403); 
assign U4868 = ~(U2493 & U2401); 
assign U4873 = ~(U2493 & U2399); 
assign U4896 = ~(U2495 & U2413); 
assign U4901 = ~(U2495 & U2411); 
assign U4906 = ~(U2495 & U2409); 
assign U4911 = ~(U2495 & U2407); 
assign U4916 = ~(U2495 & U2405); 
assign U4921 = ~(U2495 & U2403); 
assign U4926 = ~(U2495 & U2401); 
assign U4931 = ~(U2495 & U2399); 
assign U4953 = ~(U2497 & U2413); 
assign U4958 = ~(U2497 & U2411); 
assign U4963 = ~(U2497 & U2409); 
assign U4968 = ~(U2497 & U2407); 
assign U4973 = ~(U2497 & U2405); 
assign U4978 = ~(U2497 & U2403); 
assign U4983 = ~(U2497 & U2401); 
assign U4988 = ~(U2497 & U2399); 
assign U5066 = ~(U2501 & U2413); 
assign U5071 = ~(U2501 & U2411); 
assign U5076 = ~(U2501 & U2409); 
assign U5081 = ~(U2501 & U2407); 
assign U5086 = ~(U2501 & U2405); 
assign U5091 = ~(U2501 & U2403); 
assign U5096 = ~(U2501 & U2401); 
assign U5101 = ~(U2501 & U2399); 
assign U5124 = ~(U2503 & U2413); 
assign U5129 = ~(U2503 & U2411); 
assign U5134 = ~(U2503 & U2409); 
assign U5139 = ~(U2503 & U2407); 
assign U5144 = ~(U2503 & U2405); 
assign U5149 = ~(U2503 & U2403); 
assign U5154 = ~(U2503 & U2401); 
assign U5159 = ~(U2503 & U2399); 
assign U5181 = ~(U2505 & U2413); 
assign U5186 = ~(U2505 & U2411); 
assign U5191 = ~(U2505 & U2409); 
assign U5196 = ~(U2505 & U2407); 
assign U5201 = ~(U2505 & U2405); 
assign U5206 = ~(U2505 & U2403); 
assign U5211 = ~(U2505 & U2401); 
assign U5216 = ~(U2505 & U2399); 
assign U5539 = ~(U2388 & U5538); 
assign U5691 = ~(R2099_U76 & U2380); 
assign U5701 = ~(ADD_405_U80 & U2375); 
assign U5702 = ~(ADD_515_U81 & U2374); 
assign U5790 = ~(R2358_U82 & U2364); 
assign U6143 = ~(U2386 & R2358_U82); 
assign U6253 = ~(U2383 & R2358_U82); 
assign U6311 = ~(U2371 & R2099_U76); 
assign U6359 = ~(U2429 & R2358_U82); 
assign U6495 = ~(U2604 & R2099_U76); 
assign U6503 = ~(R2096_U81 & U7473); 
assign U6859 = ~(U4147 & R2144_U80); 
assign U7719 = ~(U7681 & U4515); 
assign R2278_U18 = ~(U2783 & INSTADDRPOINTER_REG_4__SCAN_IN); 
assign R2278_U20 = ~(U2782 & INSTADDRPOINTER_REG_5__SCAN_IN); 
assign R2278_U42 = ~(R2278_U402 & R2278_U401); 
assign R2278_U90 = ~(R2278_U172 & R2278_U173); 
assign R2278_U91 = ~(R2278_U166 & R2278_U175); 
assign R2278_U162 = U2780 | INSTADDRPOINTER_REG_7__SCAN_IN; 
assign R2278_U163 = ~(U2780 & INSTADDRPOINTER_REG_7__SCAN_IN); 
assign R2278_U178 = U2783 | INSTADDRPOINTER_REG_4__SCAN_IN; 
assign R2278_U179 = U2782 | INSTADDRPOINTER_REG_5__SCAN_IN; 
assign R2278_U262 = ~R2278_U100; 
assign R2278_U300 = ~(R2278_U172 & R2278_U173); 
assign R2278_U373 = ~(R2278_U171 & R2278_U100); 
assign R2358_U24 = ~U2644; 
assign R2358_U31 = ~(U2644 & R2358_U77); 
assign R2358_U65 = ~(R2358_U64 & R2358_U229); 
assign R2358_U112 = ~(R2358_U634 & R2358_U633); 
assign R2358_U124 = R2358_U231 & R2358_U229; 
assign R2358_U129 = R2358_U231 & R2358_U230; 
assign R2358_U180 = R2358_U505 & R2358_U504; 
assign R2358_U242 = ~(R2358_U452 & R2358_U451 & R2358_U23); 
assign R2358_U243 = ~(R2358_U463 & R2358_U462 & R2358_U25); 
assign R2358_U244 = ~(R2358_U465 & R2358_U464 & R2358_U26); 
assign R2358_U248 = ~(R2358_U247 & R2358_U246); 
assign R2358_U271 = ~R2358_U64; 
assign R2358_U275 = ~(R2358_U231 & R2358_U230); 
assign R2358_U334 = ~(R2358_U234 & R2358_U229); 
assign R2358_U495 = ~(R2358_U455 & U2644); 
assign R2358_U508 = ~(R2358_U507 & R2358_U506); 
assign R2144_U11 = ~(R2144_U144 & R2144_U146); 
assign R2144_U30 = ~(R2144_U209 & R2144_U208); 
assign R2144_U40 = ~(R2144_U254 & R2144_U253); 
assign R2144_U41 = ~(R2144_U256 & R2144_U255); 
assign R2144_U42 = ~(R2144_U258 & R2144_U257); 
assign R2144_U142 = ~R2144_U95; 
assign R2144_U143 = ~R2144_U26; 
assign R2144_U250 = ~(R2144_U32 & R2144_U26); 
assign R2144_U252 = ~(R2144_U33 & R2144_U95); 
assign R2099_U17 = ~(R2099_U171 & R2099_U53); 
assign R2099_U316 = ~(R2099_U252 & R2099_U171); 
assign R2096_U44 = ~(R2096_U112 & REIP_REG_21__SCAN_IN); 
assign R2096_U160 = ~(R2096_U112 & R2096_U43); 
assign ADD_405_U44 = ~(ADD_405_U115 & INSTADDRPOINTER_REG_21__SCAN_IN); 
assign ADD_405_U162 = ~(ADD_405_U115 & ADD_405_U43); 
assign ADD_515_U44 = ~(ADD_515_U112 & INSTADDRPOINTER_REG_21__SCAN_IN); 
assign ADD_515_U160 = ~(ADD_515_U112 & ADD_515_U43); 
assign U2475 = U3441 & U3345; 
assign U2490 = U7681 & U3345; 
assign U2634 = R2144_U11 & U6734; 
assign U2638 = R2144_U40 & U6734; 
assign U2639 = R2144_U41 & U6734; 
assign U2640 = R2144_U42 & U6734; 
assign U2641 = R2144_U30 & U6734; 
assign U2771 = U4147 & R2144_U11; 
assign U2775 = U4147 & R2144_U40; 
assign U2776 = U4147 & R2144_U41; 
assign U2777 = U4147 & R2144_U42; 
assign U2778 = U4147 & R2144_U30; 
assign U2779 = ~(U6860 & U6859); 
assign U2859 = ~(U6254 & U6253 & U6255); 
assign U2891 = ~(U6143 & U6142 & U6144); 
assign U2986 = ~(U5788 & U5787 & U5789 & U5791 & U5790); 
assign U3574 = U3573 & U4511; 
assign U3814 = U5699 & U5701; 
assign U3816 = U3815 & U5702; 
assign U3878 = U6361 & U6360 & U6363 & U6362 & U6359; 
assign U3914 = U6505 & U6503; 
assign U4500 = ~(U4499 & U3249); 
assign U4519 = ~U3345; 
assign U5009 = ~(U4226 & U2413); 
assign U5014 = ~(U4226 & U2411); 
assign U5019 = ~(U4226 & U2409); 
assign U5024 = ~(U4226 & U2407); 
assign U5029 = ~(U4226 & U2405); 
assign U5034 = ~(U4226 & U2403); 
assign U5039 = ~(U4226 & U2401); 
assign U5044 = ~(U4226 & U2399); 
assign U5525 = ~U3391; 
assign U5528 = ~(U3345 & U5527); 
assign U5542 = ~(U3741 & U5539); 
assign U5545 = ~(U5543 & U5544 & U4233); 
assign U5567 = ~(R2278_U42 & U2377); 
assign U5793 = ~(U2372 & R2278_U42); 
assign U5795 = ~(R2358_U112 & U2364); 
assign U6146 = ~(U2386 & R2358_U112); 
assign U6256 = ~(U2383 & R2358_U112); 
assign U6367 = ~(U2429 & R2358_U112); 
assign U7721 = ~(U7720 & U7719); 
assign R2278_U22 = ~U2770; 
assign R2278_U23 = ~(U2770 & INSTADDRPOINTER_REG_19__SCAN_IN); 
assign R2278_U33 = ~U2770; 
assign R2278_U35 = ~U2770; 
assign R2278_U36 = ~(U2770 & INSTADDRPOINTER_REG_26__SCAN_IN); 
assign R2278_U43 = R2278_U178 & R2278_U162; 
assign R2278_U47 = U2770 & INSTADDRPOINTER_REG_20__SCAN_IN; 
assign R2278_U48 = R2278_U178 & R2278_U162; 
assign R2278_U79 = ~(R2278_U162 & R2278_U163); 
assign R2278_U85 = ~(R2278_U179 & R2278_U20); 
assign R2278_U88 = ~(R2278_U178 & R2278_U18); 
assign R2278_U93 = ~U2769; 
assign R2278_U164 = U2781 | INSTADDRPOINTER_REG_6__SCAN_IN; 
assign R2278_U165 = ~(U2781 & INSTADDRPOINTER_REG_6__SCAN_IN); 
assign R2278_U174 = ~R2278_U90; 
assign R2278_U176 = ~(R2278_U300 & R2278_U166); 
assign R2278_U180 = ~R2278_U20; 
assign R2278_U181 = ~R2278_U18; 
assign R2278_U203 = ~R2278_U91; 
assign R2278_U204 = U2770 | INSTADDRPOINTER_REG_25__SCAN_IN; 
assign R2278_U205 = U2770 | INSTADDRPOINTER_REG_23__SCAN_IN; 
assign R2278_U206 = U2770 | INSTADDRPOINTER_REG_22__SCAN_IN; 
assign R2278_U207 = U2770 | INSTADDRPOINTER_REG_19__SCAN_IN; 
assign R2278_U208 = U2770 | INSTADDRPOINTER_REG_18__SCAN_IN; 
assign R2278_U227 = U2770 | INSTADDRPOINTER_REG_17__SCAN_IN; 
assign R2278_U228 = ~(U2770 & INSTADDRPOINTER_REG_17__SCAN_IN); 
assign R2278_U229 = ~(U2770 & INSTADDRPOINTER_REG_18__SCAN_IN); 
assign R2278_U231 = U2770 | INSTADDRPOINTER_REG_20__SCAN_IN; 
assign R2278_U232 = ~(U2770 & INSTADDRPOINTER_REG_20__SCAN_IN); 
assign R2278_U235 = U2770 | INSTADDRPOINTER_REG_21__SCAN_IN; 
assign R2278_U236 = ~(U2770 & INSTADDRPOINTER_REG_21__SCAN_IN); 
assign R2278_U238 = ~(U2770 & INSTADDRPOINTER_REG_22__SCAN_IN); 
assign R2278_U240 = ~(U2770 & INSTADDRPOINTER_REG_23__SCAN_IN); 
assign R2278_U242 = U2770 | INSTADDRPOINTER_REG_24__SCAN_IN; 
assign R2278_U243 = ~(U2770 & INSTADDRPOINTER_REG_24__SCAN_IN); 
assign R2278_U245 = ~(U2770 & INSTADDRPOINTER_REG_25__SCAN_IN); 
assign R2278_U246 = U2770 | INSTADDRPOINTER_REG_26__SCAN_IN; 
assign R2278_U250 = U2770 | INSTADDRPOINTER_REG_27__SCAN_IN; 
assign R2278_U251 = ~(U2770 & INSTADDRPOINTER_REG_27__SCAN_IN); 
assign R2278_U253 = U2770 | INSTADDRPOINTER_REG_28__SCAN_IN; 
assign R2278_U254 = ~(U2770 & INSTADDRPOINTER_REG_28__SCAN_IN); 
assign R2278_U256 = U2770 | INSTADDRPOINTER_REG_29__SCAN_IN; 
assign R2278_U257 = ~(U2770 & INSTADDRPOINTER_REG_29__SCAN_IN); 
assign R2278_U259 = U2770 | INSTADDRPOINTER_REG_30__SCAN_IN; 
assign R2278_U260 = ~(U2770 & INSTADDRPOINTER_REG_30__SCAN_IN); 
assign R2278_U301 = ~(R2278_U162 & U2781 & INSTADDRPOINTER_REG_6__SCAN_IN); 
assign R2278_U303 = U2781 | INSTADDRPOINTER_REG_6__SCAN_IN; 
assign R2278_U337 = U2781 | INSTADDRPOINTER_REG_6__SCAN_IN; 
assign R2278_U363 = ~(U2769 & R2278_U94); 
assign R2278_U368 = ~(U2770 & R2278_U21); 
assign R2278_U374 = ~(R2278_U262 & R2278_U99); 
assign R2278_U375 = ~(U2770 & R2278_U32); 
assign R2278_U380 = ~(U2770 & R2278_U34); 
assign R2358_U32 = ~U2642; 
assign R2358_U35 = ~U2620; 
assign R2358_U36 = ~U2625; 
assign R2358_U37 = ~U2624; 
assign R2358_U38 = ~U2622; 
assign R2358_U39 = ~U2623; 
assign R2358_U40 = ~U2621; 
assign R2358_U41 = ~U2626; 
assign R2358_U42 = ~U2627; 
assign R2358_U43 = ~U2628; 
assign R2358_U44 = ~U2629; 
assign R2358_U45 = ~U2630; 
assign R2358_U46 = ~(U2630 & R2358_U78); 
assign R2358_U49 = ~(U2642 & R2358_U490); 
assign R2358_U56 = ~U2631; 
assign R2358_U57 = ~U2632; 
assign R2358_U58 = ~U2633; 
assign R2358_U59 = ~(U2633 & R2358_U607); 
assign R2358_U87 = R2358_U246 & R2358_U243; 
assign R2358_U89 = R2358_U247 & R2358_U244; 
assign R2358_U125 = R2358_U244 & R2358_U243; 
assign R2358_U228 = ~R2358_U31; 
assign R2358_U240 = ~(R2358_U124 & R2358_U239); 
assign R2358_U263 = ~(R2358_U455 & R2358_U24); 
assign R2358_U265 = ~(R2358_U245 & R2358_U242); 
assign R2358_U267 = ~(R2358_U455 & R2358_U24); 
assign R2358_U272 = ~R2358_U65; 
assign R2358_U273 = ~(R2358_U65 & R2358_U234); 
assign R2358_U276 = ~(R2358_U65 & R2358_U234 & R2358_U275); 
assign R2358_U278 = ~(U2620 & R2358_U580); 
assign R2358_U280 = ~(U2621 & R2358_U595); 
assign R2358_U283 = ~(U2625 & R2358_U583); 
assign R2358_U284 = ~(U2624 & R2358_U586); 
assign R2358_U288 = ~(U2622 & R2358_U592); 
assign R2358_U289 = ~(U2623 & R2358_U589); 
assign R2358_U295 = ~(U2632 & R2358_U604); 
assign R2358_U316 = ~(U2631 & R2358_U598); 
assign R2358_U320 = ~(U2626 & R2358_U568); 
assign R2358_U321 = ~(U2627 & R2358_U571); 
assign R2358_U323 = ~(U2628 & R2358_U574); 
assign R2358_U326 = ~(U2629 & R2358_U577); 
assign R2358_U335 = ~(R2358_U271 & R2358_U334); 
assign R2358_U383 = ~(R2358_U246 & R2358_U243); 
assign R2358_U384 = ~(R2358_U247 & R2358_U244); 
assign R2358_U403 = ~(R2358_U77 & R2358_U242); 
assign R2358_U404 = ~(U2644 & R2358_U242); 
assign R2358_U496 = ~(R2358_U77 & R2358_U24); 
assign R2358_U628 = ~(R2358_U553 & U2630); 
assign R2144_U94 = ~(R2144_U143 & R2144_U32); 
assign R2144_U249 = ~(R2144_U222 & R2144_U143); 
assign R2144_U251 = ~(R2144_U142 & R2144_U228); 
assign R2099_U75 = ~(R2099_U317 & R2099_U316); 
assign R2099_U172 = ~R2099_U17; 
assign R2099_U315 = ~(R2099_U52 & R2099_U17); 
assign R2096_U80 = ~(R2096_U160 & R2096_U159); 
assign R2096_U113 = ~R2096_U44; 
assign R2096_U157 = ~(R2096_U44 & REIP_REG_22__SCAN_IN); 
assign ADD_405_U79 = ~(ADD_405_U162 & ADD_405_U161); 
assign ADD_405_U116 = ~ADD_405_U44; 
assign ADD_405_U159 = ~(ADD_405_U44 & INSTADDRPOINTER_REG_22__SCAN_IN); 
assign ADD_515_U80 = ~(ADD_515_U160 & ADD_515_U159); 
assign ADD_515_U113 = ~ADD_515_U44; 
assign ADD_515_U157 = ~(ADD_515_U44 & INSTADDRPOINTER_REG_22__SCAN_IN); 
assign U2499 = U4519 & U3441; 
assign U2507 = U4519 & U7681; 
assign U2827 = ~(U6357 & U6356 & U6358 & U3878); 
assign U2858 = ~(U6257 & U6258 & U6256); 
assign U2890 = ~(U6146 & U6145 & U6147); 
assign U2985 = ~(U5793 & U5792 & U5794 & U5796 & U5795); 
assign U3019 = U5525 & INSTQUEUEWR_ADDR_REG_4__SCAN_IN; 
assign U3302 = ~(U4515 & U2475); 
assign U3314 = ~(U4588 & U2475); 
assign U3321 = ~(U4646 & U2475); 
assign U3325 = ~(U2485 & U2475); 
assign U3330 = ~(U2490 & U4515); 
assign U3334 = ~(U2490 & U4588); 
assign U3337 = ~(U2490 & U4646); 
assign U3341 = ~(U2490 & U2485); 
assign U3756 = U5568 & U5567; 
assign U3879 = U6369 & U6368 & U6371 & U6370 & U6367; 
assign U5534 = ~(U2388 & U7721); 
assign U5698 = ~(R2099_U75 & U2380); 
assign U5708 = ~(ADD_405_U79 & U2375); 
assign U5709 = ~(ADD_515_U80 & U2374); 
assign U6314 = ~(U2371 & R2099_U75); 
assign U6502 = ~(U2604 & R2099_U75); 
assign U6510 = ~(R2096_U80 & U7473); 
assign U7671 = ~(U4500 & STATE2_REG_0__SCAN_IN); 
assign U7717 = ~(U5525 & INSTQUEUEWR_ADDR_REG_3__SCAN_IN); 
assign U7722 = ~(U5525 & INSTQUEUEWR_ADDR_REG_2__SCAN_IN); 
assign U7724 = ~(U5525 & INSTQUEUEWR_ADDR_REG_1__SCAN_IN); 
assign U7725 = ~(U5542 & U3391); 
assign U7726 = ~(U5525 & INSTQUEUEWR_ADDR_REG_0__SCAN_IN); 
assign U7727 = ~(U5545 & U3391); 
assign R2278_U9 = R2278_U235 & R2278_U231; 
assign R2278_U14 = R2278_U250 & R2278_U246; 
assign R2278_U24 = ~(U2771 & INSTADDRPOINTER_REG_16__SCAN_IN); 
assign R2278_U26 = ~(U2779 & INSTADDRPOINTER_REG_8__SCAN_IN); 
assign R2278_U27 = ~(U2778 & INSTADDRPOINTER_REG_9__SCAN_IN); 
assign R2278_U28 = ~(U2777 & INSTADDRPOINTER_REG_10__SCAN_IN); 
assign R2278_U29 = ~(U2775 & INSTADDRPOINTER_REG_12__SCAN_IN); 
assign R2278_U44 = R2278_U303 & R2278_U179; 
assign R2278_U49 = R2278_U337 & R2278_U179; 
assign R2278_U82 = ~(R2278_U165 & R2278_U164); 
assign R2278_U87 = ~(R2278_U175 & R2278_U176); 
assign R2278_U101 = R2278_U374 & R2278_U373; 
assign R2278_U107 = ~(R2278_U250 & R2278_U251); 
assign R2278_U109 = ~(R2278_U246 & R2278_U36); 
assign R2278_U113 = ~(R2278_U204 & R2278_U245); 
assign R2278_U116 = ~(R2278_U243 & R2278_U242); 
assign R2278_U119 = ~(R2278_U240 & R2278_U205); 
assign R2278_U122 = ~(R2278_U238 & R2278_U206); 
assign R2278_U125 = ~(R2278_U236 & R2278_U235); 
assign R2278_U127 = ~(R2278_U231 & R2278_U232); 
assign R2278_U131 = ~(R2278_U207 & R2278_U23); 
assign R2278_U134 = ~(R2278_U208 & R2278_U229); 
assign R2278_U137 = ~(R2278_U227 & R2278_U228); 
assign R2278_U182 = ~(R2278_U181 & R2278_U179 & R2278_U164 & R2278_U162); 
assign R2278_U185 = U2779 | INSTADDRPOINTER_REG_8__SCAN_IN; 
assign R2278_U189 = U2778 | INSTADDRPOINTER_REG_9__SCAN_IN; 
assign R2278_U199 = ~R2278_U79; 
assign R2278_U201 = ~R2278_U85; 
assign R2278_U202 = ~R2278_U88; 
assign R2278_U215 = U2776 | INSTADDRPOINTER_REG_11__SCAN_IN; 
assign R2278_U216 = ~(U2776 & INSTADDRPOINTER_REG_11__SCAN_IN); 
assign R2278_U217 = U2777 | INSTADDRPOINTER_REG_10__SCAN_IN; 
assign R2278_U221 = U2775 | INSTADDRPOINTER_REG_12__SCAN_IN; 
assign R2278_U225 = U2771 | INSTADDRPOINTER_REG_16__SCAN_IN; 
assign R2278_U230 = ~R2278_U23; 
assign R2278_U247 = ~R2278_U36; 
assign R2278_U302 = ~(R2278_U180 & R2278_U162 & R2278_U164); 
assign R2278_U310 = ~(R2278_U47 & R2278_U235); 
assign R2278_U361 = ~(R2278_U174 & R2278_U91); 
assign R2278_U362 = ~(R2278_U203 & R2278_U90); 
assign R2278_U364 = ~(R2278_U93 & INSTADDRPOINTER_REG_31__SCAN_IN); 
assign R2278_U369 = ~(R2278_U22 & INSTADDRPOINTER_REG_30__SCAN_IN); 
assign R2278_U376 = ~(R2278_U33 & INSTADDRPOINTER_REG_29__SCAN_IN); 
assign R2278_U381 = ~(R2278_U35 & INSTADDRPOINTER_REG_28__SCAN_IN); 
assign R2358_U33 = ~U2641; 
assign R2358_U47 = ~U2639; 
assign R2358_U48 = ~U2640; 
assign R2358_U52 = ~U2638; 
assign R2358_U53 = ~(U2638 & R2358_U531); 
assign R2358_U60 = ~U2634; 
assign R2358_U61 = ~(U2634 & R2358_U601); 
assign R2358_U128 = R2358_U265 & R2358_U31; 
assign R2358_U131 = R2358_U288 & R2358_U289; 
assign R2358_U133 = R2358_U326 & R2358_U323; 
assign R2358_U154 = R2358_U284 & R2358_U283; 
assign R2358_U178 = ~(R2358_U230 & R2358_U240); 
assign R2358_U222 = ~(R2358_U404 & R2358_U403); 
assign R2358_U225 = ~R2358_U46; 
assign R2358_U251 = ~(R2358_U228 & R2358_U242); 
assign R2358_U253 = ~(R2358_U487 & R2358_U486 & R2358_U32); 
assign R2358_U254 = ~R2358_U49; 
assign R2358_U274 = ~(R2358_U129 & R2358_U273); 
assign R2358_U277 = ~(R2358_U563 & R2358_U562 & R2358_U35); 
assign R2358_U279 = ~(R2358_U565 & R2358_U564 & R2358_U40); 
assign R2358_U281 = ~(R2358_U555 & R2358_U554 & R2358_U38); 
assign R2358_U282 = ~(R2358_U557 & R2358_U556 & R2358_U39); 
assign R2358_U285 = ~(R2358_U559 & R2358_U558 & R2358_U37); 
assign R2358_U286 = ~(R2358_U284 & R2358_U283); 
assign R2358_U293 = ~(R2358_U561 & R2358_U560 & R2358_U36); 
assign R2358_U294 = ~(R2358_U536 & R2358_U535 & R2358_U57); 
assign R2358_U296 = ~(R2358_U538 & R2358_U537 & R2358_U58); 
assign R2358_U297 = ~R2358_U59; 
assign R2358_U302 = ~(U2639 & R2358_U515); 
assign R2358_U305 = ~(U2641 & R2358_U76); 
assign R2358_U307 = ~(U2640 & R2358_U518); 
assign R2358_U317 = ~(R2358_U542 & R2358_U541 & R2358_U56); 
assign R2358_U319 = ~(R2358_U544 & R2358_U543 & R2358_U41); 
assign R2358_U322 = ~(R2358_U546 & R2358_U545 & R2358_U42); 
assign R2358_U324 = ~(R2358_U548 & R2358_U547 & R2358_U43); 
assign R2358_U325 = ~(R2358_U550 & R2358_U549 & R2358_U44); 
assign R2358_U329 = ~(R2358_U553 & R2358_U45); 
assign R2358_U336 = ~(R2358_U272 & R2358_U234); 
assign R2358_U382 = ~(R2358_U267 & R2358_U31); 
assign R2358_U405 = ~(U2640 & R2358_U518); 
assign R2358_U443 = ~(R2358_U442 & U2641); 
assign R2358_U445 = ~(R2358_U442 & U2641); 
assign R2358_U497 = ~(R2358_U496 & R2358_U495); 
assign R2358_U629 = ~(R2358_U78 & R2358_U45); 
assign R2144_U38 = ~(R2144_U250 & R2144_U249); 
assign R2144_U39 = ~(R2144_U252 & R2144_U251); 
assign R2144_U147 = ~R2144_U94; 
assign R2144_U248 = ~(R2144_U31 & R2144_U94); 
assign R2099_U18 = ~(R2099_U172 & R2099_U52); 
assign R2099_U314 = ~(R2099_U249 & R2099_U172); 
assign R2096_U46 = ~(R2096_U113 & REIP_REG_22__SCAN_IN); 
assign R2096_U158 = ~(R2096_U113 & R2096_U45); 
assign ADD_405_U46 = ~(ADD_405_U116 & INSTADDRPOINTER_REG_22__SCAN_IN); 
assign ADD_405_U160 = ~(ADD_405_U116 & ADD_405_U45); 
assign ADD_515_U46 = ~(ADD_515_U113 & INSTADDRPOINTER_REG_22__SCAN_IN); 
assign ADD_515_U158 = ~(ADD_515_U113 & ADD_515_U45); 
assign U2480 = U3302 & U4536; 
assign U2482 = U3314 & U4594; 
assign U2484 = U3321 & U4653; 
assign U2489 = U3325 & U4710; 
assign U2492 = U3330 & U4768; 
assign U2494 = U3334 & U4825; 
assign U2496 = U3337 & U4883; 
assign U2498 = U3341 & U4940; 
assign U2636 = R2144_U38 & U6734; 
assign U2637 = R2144_U39 & U6734; 
assign U2773 = U4147 & R2144_U38; 
assign U2774 = U4147 & R2144_U39; 
assign U2826 = ~(U6365 & U6364 & U6366 & U3879); 
assign U3017 = ~(U3756 & U3755 & U3758); 
assign U3346 = ~(U2499 & U4515); 
assign U3351 = ~(U2499 & U4588); 
assign U3354 = ~(U2499 & U4646); 
assign U3358 = ~(U2499 & U2485); 
assign U3361 = ~(U2507 & U4515); 
assign U3365 = ~(U2507 & U4588); 
assign U3368 = ~(U2507 & U4646); 
assign U3372 = ~(U2507 & U2485); 
assign U3464 = ~(U7725 & U7724); 
assign U3465 = ~(U7727 & U7726); 
assign U3817 = U5706 & U5708; 
assign U3819 = U3818 & U5709; 
assign U3916 = U6512 & U6510; 
assign U4520 = ~U3302; 
assign U4589 = ~U3314; 
assign U4647 = ~U3321; 
assign U4705 = ~U3325; 
assign U4762 = ~U3330; 
assign U4820 = ~U3334; 
assign U4877 = ~U3337; 
assign U4935 = ~U3341; 
assign U5537 = ~(U3740 & U5534); 
assign U5574 = ~(R2278_U101 & U2377); 
assign U5798 = ~(U2372 & R2278_U101); 
assign U7592 = ~(U7672 & U7671 & U3569); 
assign R2278_U5 = R2278_U217 & R2278_U215; 
assign R2278_U6 = R2278_U227 & R2278_U225; 
assign R2278_U10 = R2278_U9 & R2278_U206; 
assign R2278_U15 = R2278_U14 & R2278_U253; 
assign R2278_U45 = R2278_U182 & R2278_U163; 
assign R2278_U46 = R2278_U302 & R2278_U301; 
assign R2278_U50 = R2278_U301 & R2278_U163 & R2278_U182; 
assign R2278_U51 = R2278_U189 & R2278_U185; 
assign R2278_U62 = ~(R2278_U364 & R2278_U363); 
assign R2278_U63 = ~(R2278_U369 & R2278_U368); 
assign R2278_U64 = ~(R2278_U376 & R2278_U375); 
assign R2278_U65 = ~(R2278_U381 & R2278_U380); 
assign R2278_U70 = R2278_U310 & R2278_U236; 
assign R2278_U73 = ~(R2278_U189 & R2278_U27); 
assign R2278_U76 = ~(R2278_U185 & R2278_U26); 
assign R2278_U92 = R2278_U362 & R2278_U361; 
assign R2278_U141 = ~(R2278_U225 & R2278_U24); 
assign R2278_U153 = ~(R2278_U221 & R2278_U29); 
assign R2278_U156 = ~(R2278_U215 & R2278_U216); 
assign R2278_U159 = ~(R2278_U28 & R2278_U217); 
assign R2278_U177 = ~R2278_U87; 
assign R2278_U183 = ~(R2278_U43 & R2278_U87 & R2278_U44); 
assign R2278_U186 = ~R2278_U26; 
assign R2278_U190 = ~R2278_U27; 
assign R2278_U193 = ~(R2278_U178 & R2278_U87); 
assign R2278_U200 = ~R2278_U82; 
assign R2278_U218 = ~R2278_U28; 
assign R2278_U222 = ~R2278_U29; 
assign R2278_U226 = ~R2278_U24; 
assign R2278_U263 = ~R2278_U107; 
assign R2278_U264 = ~R2278_U109; 
assign R2278_U265 = ~R2278_U113; 
assign R2278_U266 = ~R2278_U116; 
assign R2278_U267 = ~R2278_U119; 
assign R2278_U268 = ~R2278_U122; 
assign R2278_U269 = ~R2278_U125; 
assign R2278_U270 = ~R2278_U127; 
assign R2278_U272 = ~R2278_U131; 
assign R2278_U273 = ~R2278_U134; 
assign R2278_U274 = ~R2278_U137; 
assign R2278_U322 = ~(R2278_U247 & R2278_U250); 
assign R2278_U334 = ~(R2278_U310 & R2278_U236); 
assign R2278_U336 = ~(R2278_U48 & R2278_U87 & R2278_U49); 
assign R2278_U360 = ~(R2278_U202 & R2278_U87); 
assign R2358_U5 = R2358_U293 & R2358_U285 & R2358_U282 & R2358_U281; 
assign R2358_U6 = R2358_U329 & R2358_U325; 
assign R2358_U9 = R2358_U296 & R2358_U294; 
assign R2358_U19 = R2358_U336 & R2358_U335; 
assign R2358_U20 = R2358_U276 & R2358_U274; 
assign R2358_U84 = R2358_U49 & R2358_U253; 
assign R2358_U92 = R2358_U278 & R2358_U277; 
assign R2358_U94 = R2358_U280 & R2358_U279; 
assign R2358_U96 = R2358_U288 & R2358_U281; 
assign R2358_U98 = R2358_U289 & R2358_U282; 
assign R2358_U100 = R2358_U285 & R2358_U284; 
assign R2358_U102 = R2358_U293 & R2358_U283; 
assign R2358_U104 = R2358_U320 & R2358_U319; 
assign R2358_U106 = R2358_U322 & R2358_U321; 
assign R2358_U108 = R2358_U324 & R2358_U323; 
assign R2358_U113 = R2358_U317 & R2358_U316; 
assign R2358_U115 = R2358_U295 & R2358_U294; 
assign R2358_U117 = R2358_U59 & R2358_U296; 
assign R2358_U127 = R2358_U245 & R2358_U222; 
assign R2358_U130 = R2358_U285 & R2358_U282; 
assign R2358_U132 = R2358_U281 & R2358_U279; 
assign R2358_U134 = R2358_U322 & R2358_U319; 
assign R2358_U135 = R2358_U279 & R2358_U277; 
assign R2358_U141 = R2358_U322 & R2358_U319; 
assign R2358_U152 = R2358_U285 & R2358_U282 & R2358_U293; 
assign R2358_U241 = ~R2358_U178; 
assign R2358_U249 = ~(R2358_U243 & R2358_U248 & R2358_U222); 
assign R2358_U250 = ~(R2358_U178 & R2358_U125 & R2358_U222); 
assign R2358_U257 = ~(R2358_U244 & R2358_U178); 
assign R2358_U298 = ~R2358_U61; 
assign R2358_U301 = ~(R2358_U510 & R2358_U509 & R2358_U48); 
assign R2358_U303 = ~(R2358_U512 & R2358_U511 & R2358_U47); 
assign R2358_U304 = ~(R2358_U442 & R2358_U33); 
assign R2358_U309 = ~R2358_U53; 
assign R2358_U310 = ~(R2358_U523 & R2358_U522 & R2358_U52); 
assign R2358_U313 = ~(R2358_U540 & R2358_U539 & R2358_U60); 
assign R2358_U327 = ~(R2358_U225 & R2358_U325); 
assign R2358_U353 = ~(R2358_U326 & R2358_U325); 
assign R2358_U381 = ~(R2358_U49 & R2358_U253); 
assign R2358_U385 = ~(R2358_U278 & R2358_U277); 
assign R2358_U386 = ~(R2358_U280 & R2358_U279); 
assign R2358_U387 = ~(R2358_U288 & R2358_U281); 
assign R2358_U388 = ~(R2358_U289 & R2358_U282); 
assign R2358_U389 = ~(R2358_U285 & R2358_U284); 
assign R2358_U390 = ~(R2358_U293 & R2358_U283); 
assign R2358_U391 = ~(R2358_U320 & R2358_U319); 
assign R2358_U392 = ~(R2358_U322 & R2358_U321); 
assign R2358_U393 = ~(R2358_U324 & R2358_U323); 
assign R2358_U394 = ~(R2358_U329 & R2358_U46); 
assign R2358_U396 = ~(R2358_U317 & R2358_U316); 
assign R2358_U397 = ~(R2358_U295 & R2358_U294); 
assign R2358_U398 = ~(R2358_U59 & R2358_U296); 
assign R2358_U424 = ~(R2358_U405 & R2358_U302); 
assign R2358_U444 = ~(R2358_U76 & R2358_U33); 
assign R2358_U446 = ~(R2358_U76 & R2358_U33); 
assign R2358_U502 = ~(R2358_U384 & R2358_U178); 
assign R2358_U630 = ~(R2358_U629 & R2358_U628); 
assign R2144_U247 = ~(R2144_U147 & R2144_U225); 
assign R2099_U74 = ~(R2099_U315 & R2099_U314); 
assign R2099_U173 = ~R2099_U18; 
assign R2099_U313 = ~(R2099_U51 & R2099_U18); 
assign R2096_U79 = ~(R2096_U158 & R2096_U157); 
assign R2096_U114 = ~R2096_U46; 
assign R2096_U155 = ~(R2096_U46 & REIP_REG_23__SCAN_IN); 
assign ADD_405_U78 = ~(ADD_405_U160 & ADD_405_U159); 
assign ADD_405_U117 = ~ADD_405_U46; 
assign ADD_405_U157 = ~(ADD_405_U46 & INSTADDRPOINTER_REG_23__SCAN_IN); 
assign ADD_515_U79 = ~(ADD_515_U158 & ADD_515_U157); 
assign ADD_515_U114 = ~ADD_515_U46; 
assign ADD_515_U155 = ~(ADD_515_U46 & INSTADDRPOINTER_REG_23__SCAN_IN); 
assign U2500 = U3346 & U3344; 
assign U2502 = U3351 & U5053; 
assign U2504 = U3354 & U5111; 
assign U2506 = U3358 & U5168; 
assign U2511 = U3361 & U5226; 
assign U2513 = U3365 & U5283; 
assign U2515 = U3368 & U5341; 
assign U2517 = U3372 & U5398; 
assign U3282 = ~(U7592 & STATE2_REG_0__SCAN_IN); 
assign U3760 = U5575 & U5574; 
assign U4505 = ~(U7592 & U4234); 
assign U4508 = ~(U2368 & U7592); 
assign U4510 = ~(U7592 & U4233); 
assign U4537 = ~(U2480 & U2358); 
assign U4543 = ~(U2480 & U2388); 
assign U4550 = ~(U2412 & U4520); 
assign U4555 = ~(U2410 & U4520); 
assign U4560 = ~(U2408 & U4520); 
assign U4565 = ~(U2406 & U4520); 
assign U4570 = ~(U2404 & U4520); 
assign U4575 = ~(U2402 & U4520); 
assign U4580 = ~(U2400 & U4520); 
assign U4585 = ~(U2398 & U4520); 
assign U4595 = ~(U2482 & U2358); 
assign U4601 = ~(U2482 & U2388); 
assign U4608 = ~(U4589 & U2412); 
assign U4613 = ~(U4589 & U2410); 
assign U4618 = ~(U4589 & U2408); 
assign U4623 = ~(U4589 & U2406); 
assign U4628 = ~(U4589 & U2404); 
assign U4633 = ~(U4589 & U2402); 
assign U4638 = ~(U4589 & U2400); 
assign U4643 = ~(U4589 & U2398); 
assign U4654 = ~(U2484 & U2358); 
assign U4660 = ~(U2484 & U2388); 
assign U4667 = ~(U4647 & U2412); 
assign U4672 = ~(U4647 & U2410); 
assign U4677 = ~(U4647 & U2408); 
assign U4682 = ~(U4647 & U2406); 
assign U4687 = ~(U4647 & U2404); 
assign U4692 = ~(U4647 & U2402); 
assign U4697 = ~(U4647 & U2400); 
assign U4702 = ~(U4647 & U2398); 
assign U4711 = ~(U2489 & U2358); 
assign U4717 = ~(U2489 & U2388); 
assign U4724 = ~(U4705 & U2412); 
assign U4729 = ~(U4705 & U2410); 
assign U4734 = ~(U4705 & U2408); 
assign U4739 = ~(U4705 & U2406); 
assign U4744 = ~(U4705 & U2404); 
assign U4749 = ~(U4705 & U2402); 
assign U4754 = ~(U4705 & U2400); 
assign U4759 = ~(U4705 & U2398); 
assign U4769 = ~(U2492 & U2358); 
assign U4775 = ~(U2492 & U2388); 
assign U4782 = ~(U4762 & U2412); 
assign U4787 = ~(U4762 & U2410); 
assign U4792 = ~(U4762 & U2408); 
assign U4797 = ~(U4762 & U2406); 
assign U4802 = ~(U4762 & U2404); 
assign U4807 = ~(U4762 & U2402); 
assign U4812 = ~(U4762 & U2400); 
assign U4817 = ~(U4762 & U2398); 
assign U4826 = ~(U2494 & U2358); 
assign U4832 = ~(U2494 & U2388); 
assign U4839 = ~(U4820 & U2412); 
assign U4844 = ~(U4820 & U2410); 
assign U4849 = ~(U4820 & U2408); 
assign U4854 = ~(U4820 & U2406); 
assign U4859 = ~(U4820 & U2404); 
assign U4864 = ~(U4820 & U2402); 
assign U4869 = ~(U4820 & U2400); 
assign U4874 = ~(U4820 & U2398); 
assign U4884 = ~(U2496 & U2358); 
assign U4890 = ~(U2496 & U2388); 
assign U4897 = ~(U4877 & U2412); 
assign U4902 = ~(U4877 & U2410); 
assign U4907 = ~(U4877 & U2408); 
assign U4912 = ~(U4877 & U2406); 
assign U4917 = ~(U4877 & U2404); 
assign U4922 = ~(U4877 & U2402); 
assign U4927 = ~(U4877 & U2400); 
assign U4932 = ~(U4877 & U2398); 
assign U4941 = ~(U2498 & U2358); 
assign U4947 = ~(U2498 & U2388); 
assign U4954 = ~(U4935 & U2412); 
assign U4959 = ~(U4935 & U2410); 
assign U4964 = ~(U4935 & U2408); 
assign U4969 = ~(U4935 & U2406); 
assign U4974 = ~(U4935 & U2404); 
assign U4979 = ~(U4935 & U2402); 
assign U4984 = ~(U4935 & U2400); 
assign U4989 = ~(U4935 & U2398); 
assign U4992 = ~U3346; 
assign U5048 = ~U3351; 
assign U5105 = ~U3354; 
assign U5163 = ~U3358; 
assign U5220 = ~U3361; 
assign U5278 = ~U3365; 
assign U5335 = ~U3368; 
assign U5393 = ~U3372; 
assign U5529 = ~(U3346 & U5528); 
assign U5581 = ~(R2278_U92 & U2377); 
assign U5705 = ~(R2099_U74 & U2380); 
assign U5715 = ~(ADD_405_U78 & U2375); 
assign U5716 = ~(ADD_515_U79 & U2374); 
assign U5800 = ~(R2358_U19 & U2364); 
assign U5803 = ~(U2372 & R2278_U92); 
assign U5805 = ~(R2358_U20 & U2364); 
assign U6149 = ~(U2386 & R2358_U19); 
assign U6152 = ~(U2386 & R2358_U20); 
assign U6259 = ~(U2383 & R2358_U19); 
assign U6262 = ~(U2383 & R2358_U20); 
assign U6317 = ~(U2371 & R2099_U74); 
assign U6375 = ~(U2429 & R2358_U19); 
assign U6383 = ~(U2429 & R2358_U20); 
assign U6509 = ~(U2604 & R2099_U74); 
assign U6517 = ~(R2096_U79 & U7473); 
assign U7678 = ~(U7592 & U4509 & U3281); 
assign U7723 = ~(U5537 & U3391); 
assign R2278_U7 = R2278_U6 & R2278_U208; 
assign R2278_U11 = R2278_U10 & R2278_U205; 
assign R2278_U16 = R2278_U15 & R2278_U256; 
assign R2278_U30 = ~(U2773 & INSTADDRPOINTER_REG_14__SCAN_IN); 
assign R2278_U31 = ~(U2774 & INSTADDRPOINTER_REG_13__SCAN_IN); 
assign R2278_U39 = ~(R2278_U322 & R2278_U251); 
assign R2278_U52 = R2278_U5 & R2278_U51; 
assign R2278_U53 = R2278_U186 & R2278_U189; 
assign R2278_U75 = ~(R2278_U46 & R2278_U183 & R2278_U45); 
assign R2278_U84 = ~(R2278_U18 & R2278_U193); 
assign R2278_U191 = ~R2278_U73; 
assign R2278_U192 = ~R2278_U76; 
assign R2278_U211 = U2773 | INSTADDRPOINTER_REG_14__SCAN_IN; 
assign R2278_U213 = U2774 | INSTADDRPOINTER_REG_13__SCAN_IN; 
assign R2278_U275 = ~R2278_U141; 
assign R2278_U285 = ~R2278_U153; 
assign R2278_U290 = ~R2278_U156; 
assign R2278_U291 = ~R2278_U159; 
assign R2278_U295 = ~(R2278_U190 & R2278_U5); 
assign R2278_U296 = ~(R2278_U218 & R2278_U5); 
assign R2278_U304 = ~(R2278_U226 & R2278_U227); 
assign R2278_U312 = ~(R2278_U334 & R2278_U206); 
assign R2278_U335 = ~(R2278_U336 & R2278_U302 & R2278_U50); 
assign R2278_U359 = ~(R2278_U177 & R2278_U88); 
assign R2278_U365 = ~R2278_U62; 
assign R2278_U370 = ~R2278_U63; 
assign R2278_U377 = ~R2278_U64; 
assign R2278_U382 = ~R2278_U65; 
assign R2358_U7 = R2358_U6 & R2358_U324 & R2358_U141; 
assign R2358_U8 = R2358_U135 & R2358_U5; 
assign R2358_U10 = R2358_U304 & R2358_U253; 
assign R2358_U11 = R2358_U303 & R2358_U301; 
assign R2358_U50 = ~U2637; 
assign R2358_U51 = ~(U2637 & R2358_U80); 
assign R2358_U54 = ~U2636; 
assign R2358_U121 = R2358_U310 & R2358_U53; 
assign R2358_U126 = R2358_U249 & R2358_U245; 
assign R2358_U142 = R2358_U317 & R2358_U313; 
assign R2358_U147 = R2358_U313 & R2358_U317; 
assign R2358_U151 = R2358_U5 & R2358_U279; 
assign R2358_U156 = R2358_U6 & R2358_U324; 
assign R2358_U158 = R2358_U6 & R2358_U326; 
assign R2358_U159 = R2358_U313 & R2358_U9; 
assign R2358_U162 = R2358_U303 & R2358_U302; 
assign R2358_U165 = R2358_U444 & R2358_U443; 
assign R2358_U177 = ~(R2358_U247 & R2358_U257); 
assign R2358_U227 = ~(U2636 & R2358_U79); 
assign R2358_U287 = ~(R2358_U130 & R2358_U286); 
assign R2358_U358 = ~(R2358_U313 & R2358_U61); 
assign R2358_U375 = ~(R2358_U303 & R2358_U302); 
assign R2358_U377 = ~(R2358_U307 & R2358_U301); 
assign R2358_U401 = ~(R2358_U310 & R2358_U53); 
assign R2358_U407 = ~(R2358_U297 & R2358_U9); 
assign R2358_U408 = ~(R2358_U298 & R2358_U9); 
assign R2358_U414 = ~(R2358_U254 & R2358_U304); 
assign R2358_U425 = ~(R2358_U424 & R2358_U303); 
assign R2358_U436 = ~(R2358_U133 & R2358_U327); 
assign R2358_U447 = ~(R2358_U446 & R2358_U445); 
assign R2358_U503 = ~(R2358_U89 & R2358_U241); 
assign R2358_U641 = ~(R2358_U521 & U2636); 
assign R2358_U646 = ~(R2358_U526 & U2637); 
assign R2144_U37 = ~(R2144_U248 & R2144_U247); 
assign R2099_U19 = ~(R2099_U173 & R2099_U51); 
assign R2099_U312 = ~(R2099_U246 & R2099_U173); 
assign R2096_U48 = ~(R2096_U114 & REIP_REG_23__SCAN_IN); 
assign R2096_U156 = ~(R2096_U114 & R2096_U47); 
assign ADD_405_U48 = ~(ADD_405_U117 & INSTADDRPOINTER_REG_23__SCAN_IN); 
assign ADD_405_U158 = ~(ADD_405_U117 & ADD_405_U47); 
assign ADD_515_U48 = ~(ADD_515_U114 & INSTADDRPOINTER_REG_23__SCAN_IN); 
assign ADD_515_U156 = ~(ADD_515_U114 & ADD_515_U47); 
assign U2635 = R2144_U37 & U6734; 
assign U2772 = U4147 & R2144_U37; 
assign U2856 = ~(U6263 & U6264 & U6262); 
assign U2857 = ~(U6260 & U6261 & U6259); 
assign U2888 = ~(U6153 & U6151 & U6152); 
assign U2889 = ~(U6150 & U6148 & U6149); 
assign U2983 = ~(U5804 & U5802 & U5803 & U5806 & U5805); 
assign U2984 = ~(U5799 & U5797 & U5798 & U5801 & U5800); 
assign U3016 = ~(U3760 & U3759 & U3762); 
assign U3463 = ~(U7723 & U7722); 
assign U3576 = U4549 & U4548 & U4550; 
assign U3577 = U4554 & U4553 & U4555; 
assign U3578 = U4559 & U4558 & U4560; 
assign U3579 = U4564 & U4563 & U4565; 
assign U3580 = U4569 & U4568 & U4570; 
assign U3581 = U4574 & U4573 & U4575; 
assign U3582 = U4579 & U4578 & U4580; 
assign U3583 = U4584 & U4583 & U4585; 
assign U3585 = U4607 & U4606 & U4608; 
assign U3586 = U4612 & U4611 & U4613; 
assign U3587 = U4617 & U4616 & U4618; 
assign U3588 = U4622 & U4621 & U4623; 
assign U3589 = U4627 & U4626 & U4628; 
assign U3590 = U4632 & U4631 & U4633; 
assign U3591 = U4637 & U4636 & U4638; 
assign U3592 = U4642 & U4641 & U4643; 
assign U3594 = U4666 & U4665 & U4667; 
assign U3595 = U4671 & U4670 & U4672; 
assign U3596 = U4676 & U4675 & U4677; 
assign U3597 = U4681 & U4680 & U4682; 
assign U3598 = U4686 & U4685 & U4687; 
assign U3599 = U4691 & U4690 & U4692; 
assign U3600 = U4696 & U4695 & U4697; 
assign U3601 = U4701 & U4700 & U4702; 
assign U3603 = U4723 & U4722 & U4724; 
assign U3604 = U4728 & U4727 & U4729; 
assign U3605 = U4733 & U4732 & U4734; 
assign U3606 = U4738 & U4737 & U4739; 
assign U3607 = U4743 & U4742 & U4744; 
assign U3608 = U4748 & U4747 & U4749; 
assign U3609 = U4753 & U4752 & U4754; 
assign U3610 = U4758 & U4757 & U4759; 
assign U3612 = U4781 & U4780 & U4782; 
assign U3613 = U4786 & U4785 & U4787; 
assign U3614 = U4791 & U4790 & U4792; 
assign U3615 = U4796 & U4795 & U4797; 
assign U3616 = U4801 & U4800 & U4802; 
assign U3617 = U4806 & U4805 & U4807; 
assign U3618 = U4811 & U4810 & U4812; 
assign U3619 = U4816 & U4815 & U4817; 
assign U3621 = U4838 & U4837 & U4839; 
assign U3622 = U4843 & U4842 & U4844; 
assign U3623 = U4848 & U4847 & U4849; 
assign U3624 = U4853 & U4852 & U4854; 
assign U3625 = U4858 & U4857 & U4859; 
assign U3626 = U4863 & U4862 & U4864; 
assign U3627 = U4868 & U4867 & U4869; 
assign U3628 = U4873 & U4872 & U4874; 
assign U3630 = U4896 & U4895 & U4897; 
assign U3631 = U4901 & U4900 & U4902; 
assign U3632 = U4906 & U4905 & U4907; 
assign U3633 = U4911 & U4910 & U4912; 
assign U3634 = U4916 & U4915 & U4917; 
assign U3635 = U4921 & U4920 & U4922; 
assign U3636 = U4926 & U4925 & U4927; 
assign U3637 = U4931 & U4930 & U4932; 
assign U3639 = U4953 & U4952 & U4954; 
assign U3640 = U4958 & U4957 & U4959; 
assign U3641 = U4963 & U4962 & U4964; 
assign U3642 = U4968 & U4967 & U4969; 
assign U3643 = U4973 & U4972 & U4974; 
assign U3644 = U4978 & U4977 & U4979; 
assign U3645 = U4983 & U4982 & U4984; 
assign U3646 = U4988 & U4987 & U4989; 
assign U3764 = U3765 & U5583 & U5581; 
assign U3820 = U5713 & U5715; 
assign U3822 = U3821 & U5716; 
assign U3880 = U6377 & U6376 & U6379 & U6378 & U6375; 
assign U3881 = U6385 & U6384 & U6387 & U6386 & U6383; 
assign U3918 = U6519 & U6517; 
assign U4502 = ~U3282; 
assign U4504 = ~(U3282 & STATE2_REG_2__SCAN_IN); 
assign U4507 = ~(U4505 & STATE2_REG_1__SCAN_IN); 
assign U4538 = ~(U3307 & U4537); 
assign U4544 = ~(U3307 & U4543); 
assign U4596 = ~(U3307 & U4595); 
assign U4602 = ~(U3307 & U4601); 
assign U4655 = ~(U3307 & U4654); 
assign U4661 = ~(U3307 & U4660); 
assign U4712 = ~(U3307 & U4711); 
assign U4718 = ~(U3307 & U4717); 
assign U4770 = ~(U3307 & U4769); 
assign U4776 = ~(U3307 & U4775); 
assign U4827 = ~(U3307 & U4826); 
assign U4833 = ~(U3307 & U4832); 
assign U4885 = ~(U3307 & U4884); 
assign U4891 = ~(U3307 & U4890); 
assign U4942 = ~(U3307 & U4941); 
assign U4948 = ~(U3307 & U4947); 
assign U4997 = ~(U2500 & U2358); 
assign U5003 = ~(U2500 & U2388); 
assign U5010 = ~(U4992 & U2412); 
assign U5015 = ~(U4992 & U2410); 
assign U5020 = ~(U4992 & U2408); 
assign U5025 = ~(U4992 & U2406); 
assign U5030 = ~(U4992 & U2404); 
assign U5035 = ~(U4992 & U2402); 
assign U5040 = ~(U4992 & U2400); 
assign U5045 = ~(U4992 & U2398); 
assign U5054 = ~(U2502 & U2358); 
assign U5060 = ~(U2502 & U2388); 
assign U5067 = ~(U5048 & U2412); 
assign U5072 = ~(U5048 & U2410); 
assign U5077 = ~(U5048 & U2408); 
assign U5082 = ~(U5048 & U2406); 
assign U5087 = ~(U5048 & U2404); 
assign U5092 = ~(U5048 & U2402); 
assign U5097 = ~(U5048 & U2400); 
assign U5102 = ~(U5048 & U2398); 
assign U5112 = ~(U2504 & U2358); 
assign U5118 = ~(U2504 & U2388); 
assign U5125 = ~(U5105 & U2412); 
assign U5130 = ~(U5105 & U2410); 
assign U5135 = ~(U5105 & U2408); 
assign U5140 = ~(U5105 & U2406); 
assign U5145 = ~(U5105 & U2404); 
assign U5150 = ~(U5105 & U2402); 
assign U5155 = ~(U5105 & U2400); 
assign U5160 = ~(U5105 & U2398); 
assign U5169 = ~(U2506 & U2358); 
assign U5175 = ~(U2506 & U2388); 
assign U5182 = ~(U5163 & U2412); 
assign U5187 = ~(U5163 & U2410); 
assign U5192 = ~(U5163 & U2408); 
assign U5197 = ~(U5163 & U2406); 
assign U5202 = ~(U5163 & U2404); 
assign U5207 = ~(U5163 & U2402); 
assign U5212 = ~(U5163 & U2400); 
assign U5217 = ~(U5163 & U2398); 
assign U5227 = ~(U2511 & U2358); 
assign U5233 = ~(U2511 & U2388); 
assign U5240 = ~(U5220 & U2412); 
assign U5245 = ~(U5220 & U2410); 
assign U5250 = ~(U5220 & U2408); 
assign U5255 = ~(U5220 & U2406); 
assign U5260 = ~(U5220 & U2404); 
assign U5265 = ~(U5220 & U2402); 
assign U5270 = ~(U5220 & U2400); 
assign U5275 = ~(U5220 & U2398); 
assign U5284 = ~(U2513 & U2358); 
assign U5290 = ~(U2513 & U2388); 
assign U5297 = ~(U5278 & U2412); 
assign U5302 = ~(U5278 & U2410); 
assign U5307 = ~(U5278 & U2408); 
assign U5312 = ~(U5278 & U2406); 
assign U5317 = ~(U5278 & U2404); 
assign U5322 = ~(U5278 & U2402); 
assign U5327 = ~(U5278 & U2400); 
assign U5332 = ~(U5278 & U2398); 
assign U5342 = ~(U2515 & U2358); 
assign U5348 = ~(U2515 & U2388); 
assign U5355 = ~(U5335 & U2412); 
assign U5360 = ~(U5335 & U2410); 
assign U5365 = ~(U5335 & U2408); 
assign U5370 = ~(U5335 & U2406); 
assign U5375 = ~(U5335 & U2404); 
assign U5380 = ~(U5335 & U2402); 
assign U5385 = ~(U5335 & U2400); 
assign U5390 = ~(U5335 & U2398); 
assign U5399 = ~(U2517 & U2358); 
assign U5405 = ~(U2517 & U2388); 
assign U5412 = ~(U5393 & U2412); 
assign U5417 = ~(U5393 & U2410); 
assign U5422 = ~(U5393 & U2408); 
assign U5427 = ~(U5393 & U2406); 
assign U5431 = ~(U5393 & U2404); 
assign U5436 = ~(U5393 & U2402); 
assign U5441 = ~(U5393 & U2400); 
assign U5446 = ~(U5393 & U2398); 
assign U5530 = ~(U2388 & U5529); 
assign U7673 = ~(U3282 & STATE2_REG_3__SCAN_IN); 
assign U7677 = ~(U4510 & STATE2_REG_0__SCAN_IN); 
assign R2278_U8 = R2278_U7 & R2278_U207; 
assign R2278_U12 = R2278_U11 & R2278_U242; 
assign R2278_U41 = ~(R2278_U304 & R2278_U228); 
assign R2278_U60 = R2278_U16 & R2278_U259; 
assign R2278_U69 = R2278_U312 & R2278_U238; 
assign R2278_U89 = R2278_U360 & R2278_U359; 
assign R2278_U147 = ~(R2278_U30 & R2278_U211); 
assign R2278_U150 = ~(R2278_U213 & R2278_U31); 
assign R2278_U184 = ~R2278_U75; 
assign R2278_U187 = ~(R2278_U185 & R2278_U75); 
assign R2278_U194 = ~R2278_U84; 
assign R2278_U195 = ~(R2278_U84 & R2278_U179); 
assign R2278_U212 = ~R2278_U30; 
assign R2278_U214 = ~R2278_U31; 
assign R2278_U219 = ~(R2278_U52 & R2278_U335); 
assign R2278_U293 = ~(R2278_U53 & R2278_U5); 
assign R2278_U314 = ~(R2278_U312 & R2278_U238); 
assign R2278_U323 = ~R2278_U39; 
assign R2278_U325 = ~(R2278_U39 & R2278_U253); 
assign R2278_U352 = ~(R2278_U192 & R2278_U75); 
assign R2278_U358 = ~(R2278_U201 & R2278_U84); 
assign R2358_U12 = R2358_U8 & R2358_U7; 
assign R2358_U55 = ~(R2358_U142 & R2358_U9); 
assign R2358_U69 = ~(R2358_U407 & R2358_U295 & R2358_U408); 
assign R2358_U73 = ~(R2358_U414 & R2358_U305); 
assign R2358_U90 = ~(R2358_U503 & R2358_U502); 
assign R2358_U136 = R2358_U11 & R2358_U10; 
assign R2358_U149 = R2358_U9 & R2358_U147; 
assign R2358_U153 = R2358_U289 & R2358_U287; 
assign R2358_U163 = R2358_U375 & R2358_U307; 
assign R2358_U176 = ~(R2358_U251 & R2358_U250 & R2358_U126); 
assign R2358_U223 = ~R2358_U51; 
assign R2358_U224 = ~(R2358_U521 & R2358_U54); 
assign R2358_U258 = ~R2358_U177; 
assign R2358_U259 = ~(R2358_U177 & R2358_U243); 
assign R2358_U290 = ~(R2358_U131 & R2358_U287); 
assign R2358_U311 = ~(R2358_U526 & R2358_U50); 
assign R2358_U363 = ~(R2358_U526 & R2358_U50); 
assign R2358_U371 = ~(R2358_U526 & R2358_U50); 
assign R2358_U428 = ~(R2358_U534 & R2358_U227); 
assign R2358_U437 = ~(R2358_U436 & R2358_U324); 
assign R2358_U500 = ~(R2358_U383 & R2358_U177); 
assign R2358_U642 = ~(R2358_U79 & R2358_U54); 
assign R2358_U647 = ~(R2358_U80 & R2358_U50); 
assign R2099_U73 = ~(R2099_U313 & R2099_U312); 
assign R2099_U174 = ~R2099_U19; 
assign R2099_U311 = ~(R2099_U50 & R2099_U19); 
assign R2096_U78 = ~(R2096_U156 & R2096_U155); 
assign R2096_U115 = ~R2096_U48; 
assign R2096_U153 = ~(R2096_U48 & REIP_REG_24__SCAN_IN); 
assign ADD_405_U77 = ~(ADD_405_U158 & ADD_405_U157); 
assign ADD_405_U118 = ~ADD_405_U48; 
assign ADD_405_U155 = ~(ADD_405_U48 & INSTADDRPOINTER_REG_24__SCAN_IN); 
assign ADD_515_U78 = ~(ADD_515_U156 & ADD_515_U155); 
assign ADD_515_U115 = ~ADD_515_U48; 
assign ADD_515_U153 = ~(ADD_515_U48 & INSTADDRPOINTER_REG_24__SCAN_IN); 
assign U2824 = ~(U6381 & U6380 & U6382 & U3881); 
assign U2825 = ~(U6373 & U6372 & U6374 & U3880); 
assign U3015 = ~(U3763 & U3764); 
assign U3148 = ~(U7678 & U7677 & U3574); 
assign U3150 = ~(U3570 & U4504); 
assign U3648 = U5009 & U5008 & U5010; 
assign U3649 = U5014 & U5013 & U5015; 
assign U3650 = U5019 & U5018 & U5020; 
assign U3651 = U5024 & U5023 & U5025; 
assign U3652 = U5029 & U5028 & U5030; 
assign U3653 = U5034 & U5033 & U5035; 
assign U3654 = U5039 & U5038 & U5040; 
assign U3655 = U5044 & U5043 & U5045; 
assign U3657 = U5066 & U5065 & U5067; 
assign U3658 = U5071 & U5070 & U5072; 
assign U3659 = U5076 & U5075 & U5077; 
assign U3660 = U5081 & U5080 & U5082; 
assign U3661 = U5086 & U5085 & U5087; 
assign U3662 = U5091 & U5090 & U5092; 
assign U3663 = U5096 & U5095 & U5097; 
assign U3664 = U5101 & U5100 & U5102; 
assign U3666 = U5124 & U5123 & U5125; 
assign U3667 = U5129 & U5128 & U5130; 
assign U3668 = U5134 & U5133 & U5135; 
assign U3669 = U5139 & U5138 & U5140; 
assign U3670 = U5144 & U5143 & U5145; 
assign U3671 = U5149 & U5148 & U5150; 
assign U3672 = U5154 & U5153 & U5155; 
assign U3673 = U5159 & U5158 & U5160; 
assign U3675 = U5181 & U5180 & U5182; 
assign U3676 = U5186 & U5185 & U5187; 
assign U3677 = U5191 & U5190 & U5192; 
assign U3678 = U5196 & U5195 & U5197; 
assign U3679 = U5201 & U5200 & U5202; 
assign U3680 = U5206 & U5205 & U5207; 
assign U3681 = U5211 & U5210 & U5212; 
assign U3682 = U5216 & U5215 & U5217; 
assign U3684 = U5239 & U5238 & U5240; 
assign U3685 = U5244 & U5243 & U5245; 
assign U3686 = U5249 & U5248 & U5250; 
assign U3687 = U5254 & U5253 & U5255; 
assign U3688 = U5259 & U5258 & U5260; 
assign U3689 = U5264 & U5263 & U5265; 
assign U3690 = U5269 & U5268 & U5270; 
assign U3691 = U5274 & U5273 & U5275; 
assign U3693 = U5296 & U5295 & U5297; 
assign U3694 = U5301 & U5300 & U5302; 
assign U3695 = U5306 & U5305 & U5307; 
assign U3696 = U5311 & U5310 & U5312; 
assign U3697 = U5316 & U5315 & U5317; 
assign U3698 = U5321 & U5320 & U5322; 
assign U3699 = U5326 & U5325 & U5327; 
assign U3700 = U5331 & U5330 & U5332; 
assign U3702 = U5354 & U5353 & U5355; 
assign U3703 = U5359 & U5358 & U5360; 
assign U3704 = U5364 & U5363 & U5365; 
assign U3705 = U5369 & U5368 & U5370; 
assign U3706 = U5374 & U5373 & U5375; 
assign U3707 = U5379 & U5378 & U5380; 
assign U3708 = U5384 & U5383 & U5385; 
assign U3709 = U5389 & U5388 & U5390; 
assign U3711 = U5411 & U5410 & U5412; 
assign U3712 = U5416 & U5415 & U5417; 
assign U3713 = U5421 & U5420 & U5422; 
assign U3714 = U5426 & U5425 & U5427; 
assign U3715 = U5430 & U5429 & U5431; 
assign U3716 = U5435 & U5434 & U5436; 
assign U3717 = U5440 & U5439 & U5441; 
assign U3718 = U5445 & U5444 & U5446; 
assign U4506 = ~(U3571 & U4502); 
assign U4539 = ~(U4524 & U4538); 
assign U4545 = ~(U4544 & U3308); 
assign U4597 = ~(U4592 & U4596); 
assign U4603 = ~(U4602 & U3315); 
assign U4656 = ~(U4650 & U4655); 
assign U4662 = ~(U4661 & U3322); 
assign U4713 = ~(U4708 & U4712); 
assign U4719 = ~(U4718 & U3326); 
assign U4771 = ~(U4765 & U4770); 
assign U4777 = ~(U4776 & U3331); 
assign U4828 = ~(U4823 & U4827); 
assign U4834 = ~(U4833 & U3335); 
assign U4886 = ~(U4880 & U4885); 
assign U4892 = ~(U4891 & U3338); 
assign U4943 = ~(U4938 & U4942); 
assign U4949 = ~(U4948 & U3342); 
assign U4998 = ~(U3307 & U4997); 
assign U5004 = ~(U3307 & U5003); 
assign U5055 = ~(U3307 & U5054); 
assign U5061 = ~(U3307 & U5060); 
assign U5113 = ~(U3307 & U5112); 
assign U5119 = ~(U3307 & U5118); 
assign U5170 = ~(U3307 & U5169); 
assign U5176 = ~(U3307 & U5175); 
assign U5228 = ~(U3307 & U5227); 
assign U5234 = ~(U3307 & U5233); 
assign U5285 = ~(U3307 & U5284); 
assign U5291 = ~(U3307 & U5290); 
assign U5343 = ~(U3307 & U5342); 
assign U5349 = ~(U3307 & U5348); 
assign U5400 = ~(U3307 & U5399); 
assign U5406 = ~(U3307 & U5405); 
assign U5533 = ~(U3739 & U5530); 
assign U5588 = ~(R2278_U89 & U2377); 
assign U5712 = ~(R2099_U73 & U2380); 
assign U5722 = ~(ADD_405_U77 & U2375); 
assign U5723 = ~(ADD_515_U78 & U2374); 
assign U5808 = ~(U2372 & R2278_U89); 
assign U5810 = ~(R2358_U90 & U2364); 
assign U6155 = ~(U2386 & R2358_U90); 
assign U6265 = ~(U2383 & R2358_U90); 
assign U6320 = ~(U2371 & R2099_U73); 
assign U6391 = ~(U2429 & R2358_U90); 
assign U6516 = ~(U2604 & R2099_U73); 
assign U6524 = ~(R2096_U78 & U7473); 
assign U7674 = ~(U2428 & U4502); 
assign R2278_U13 = R2278_U12 & R2278_U204; 
assign R2278_U38 = ~(R2278_U325 & R2278_U254); 
assign R2278_U54 = R2278_U293 & R2278_U216 & R2278_U296 & R2278_U295; 
assign R2278_U71 = R2278_U293 & R2278_U216 & R2278_U296 & R2278_U295; 
assign R2278_U72 = ~(R2278_U26 & R2278_U187); 
assign R2278_U81 = ~(R2278_U20 & R2278_U195); 
assign R2278_U209 = U2772 | INSTADDRPOINTER_REG_15__SCAN_IN; 
assign R2278_U210 = ~(U2772 & INSTADDRPOINTER_REG_15__SCAN_IN); 
assign R2278_U283 = ~R2278_U147; 
assign R2278_U284 = ~R2278_U150; 
assign R2278_U305 = ~R2278_U41; 
assign R2278_U306 = ~(R2278_U41 & R2278_U208); 
assign R2278_U315 = ~(R2278_U314 & R2278_U205); 
assign R2278_U351 = ~(R2278_U184 & R2278_U76); 
assign R2278_U357 = ~(R2278_U194 & R2278_U85); 
assign R2358_U34 = ~(R2358_U246 & R2358_U259); 
assign R2358_U71 = ~U2635; 
assign R2358_U138 = R2358_U310 & R2358_U224; 
assign R2358_U148 = R2358_U7 & R2358_U149; 
assign R2358_U252 = ~R2358_U176; 
assign R2358_U255 = ~(R2358_U253 & R2358_U176); 
assign R2358_U291 = ~(R2358_U132 & R2358_U290); 
assign R2358_U300 = ~(U2635 & R2358_U81); 
assign R2358_U328 = ~(R2358_U437 & R2358_U321); 
assign R2358_U337 = ~(R2358_U290 & R2358_U281); 
assign R2358_U399 = ~(R2358_U227 & R2358_U224); 
assign R2358_U400 = ~(R2358_U371 & R2358_U51); 
assign R2358_U412 = ~R2358_U69; 
assign R2358_U413 = ~(R2358_U10 & R2358_U176); 
assign R2358_U417 = ~(R2358_U69 & R2358_U317); 
assign R2358_U423 = ~R2358_U73; 
assign R2358_U426 = ~R2358_U55; 
assign R2358_U431 = ~(R2358_U136 & R2358_U176); 
assign R2358_U432 = ~(R2358_U11 & R2358_U73); 
assign R2358_U493 = ~(R2358_U381 & R2358_U176); 
assign R2358_U501 = ~(R2358_U87 & R2358_U258); 
assign R2358_U643 = ~(R2358_U642 & R2358_U641); 
assign R2358_U648 = ~(R2358_U647 & R2358_U646); 
assign R2099_U20 = ~(R2099_U174 & R2099_U50); 
assign R2099_U310 = ~(R2099_U243 & R2099_U174); 
assign R2096_U50 = ~(R2096_U115 & REIP_REG_24__SCAN_IN); 
assign R2096_U154 = ~(R2096_U115 & R2096_U49); 
assign ADD_405_U50 = ~(ADD_405_U118 & INSTADDRPOINTER_REG_24__SCAN_IN); 
assign ADD_405_U156 = ~(ADD_405_U118 & ADD_405_U49); 
assign ADD_515_U50 = ~(ADD_515_U115 & INSTADDRPOINTER_REG_24__SCAN_IN); 
assign ADD_515_U154 = ~(ADD_515_U115 & ADD_515_U49); 
assign U2823 = ~(U3882 & U6389 & U3883 & U6391 & U6390); 
assign U2855 = ~(U6266 & U6267 & U6265); 
assign U2887 = ~(U6156 & U6154 & U6155); 
assign U2982 = ~(U5809 & U5807 & U5808 & U5811 & U5810); 
assign U3014 = ~(U3766 & U3768 & U5588); 
assign U3149 = ~(U4508 & U4507 & U4506 & U4232); 
assign U3453 = ~(U7674 & U7673); 
assign U3823 = U5720 & U5722; 
assign U3825 = U3824 & U5723; 
assign U3920 = U6526 & U6524; 
assign U4542 = ~(U4539 & U3575); 
assign U4547 = ~(U4546 & U4545); 
assign U4600 = ~(U4597 & U3584); 
assign U4605 = ~(U4604 & U4603); 
assign U4659 = ~(U4656 & U3593); 
assign U4664 = ~(U4663 & U4662); 
assign U4716 = ~(U4713 & U3602); 
assign U4721 = ~(U4720 & U4719); 
assign U4774 = ~(U4771 & U3611); 
assign U4779 = ~(U4778 & U4777); 
assign U4831 = ~(U4828 & U3620); 
assign U4836 = ~(U4835 & U4834); 
assign U4889 = ~(U4886 & U3629); 
assign U4894 = ~(U4893 & U4892); 
assign U4946 = ~(U4943 & U3638); 
assign U4951 = ~(U4950 & U4949); 
assign U4999 = ~(U4994 & U4998); 
assign U5005 = ~(U5004 & U3348); 
assign U5056 = ~(U5051 & U5055); 
assign U5062 = ~(U5061 & U3352); 
assign U5114 = ~(U5108 & U5113); 
assign U5120 = ~(U5119 & U3355); 
assign U5171 = ~(U5166 & U5170); 
assign U5177 = ~(U5176 & U3359); 
assign U5229 = ~(U5223 & U5228); 
assign U5235 = ~(U5234 & U3362); 
assign U5286 = ~(U5281 & U5285); 
assign U5292 = ~(U5291 & U3366); 
assign U5344 = ~(U5338 & U5343); 
assign U5350 = ~(U5349 & U3369); 
assign U5401 = ~(U5396 & U5400); 
assign U5407 = ~(U5406 & U3373); 
assign U7718 = ~(U5533 & U3391); 
assign R2278_U40 = ~(R2278_U306 & R2278_U229); 
assign R2278_U55 = R2278_U211 & R2278_U213 & R2278_U221 & R2278_U209; 
assign R2278_U57 = R2278_U13 & R2278_U8; 
assign R2278_U68 = R2278_U315 & R2278_U240; 
assign R2278_U77 = R2278_U352 & R2278_U351; 
assign R2278_U86 = R2278_U358 & R2278_U357; 
assign R2278_U144 = ~(R2278_U209 & R2278_U210); 
assign R2278_U152 = ~(R2278_U219 & R2278_U71); 
assign R2278_U188 = ~R2278_U72; 
assign R2278_U196 = ~R2278_U81; 
assign R2278_U197 = ~(R2278_U81 & R2278_U164); 
assign R2278_U286 = ~(R2278_U189 & R2278_U72); 
assign R2278_U294 = ~(R2278_U222 & R2278_U213 & R2278_U211 & R2278_U209); 
assign R2278_U297 = ~(R2278_U212 & R2278_U209); 
assign R2278_U298 = ~(R2278_U211 & R2278_U214 & R2278_U209); 
assign R2278_U317 = ~(R2278_U315 & R2278_U240); 
assign R2278_U326 = ~R2278_U38; 
assign R2278_U328 = ~(R2278_U38 & R2278_U256); 
assign R2278_U332 = ~(R2278_U230 & R2278_U13); 
assign R2278_U338 = ~(R2278_U219 & R2278_U54); 
assign R2278_U350 = ~(R2278_U191 & R2278_U72); 
assign R2278_U356 = ~(R2278_U200 & R2278_U81); 
assign R2358_U63 = ~(R2358_U280 & R2358_U291); 
assign R2358_U66 = ~(R2358_U417 & R2358_U316); 
assign R2358_U74 = ~(R2358_U423 & R2358_U413); 
assign R2358_U88 = ~(R2358_U501 & R2358_U500); 
assign R2358_U137 = R2358_U432 & R2358_U425; 
assign R2358_U143 = R2358_U12 & R2358_U426; 
assign R2358_U175 = ~(R2358_U49 & R2358_U255); 
assign R2358_U260 = ~R2358_U34; 
assign R2358_U264 = ~(R2358_U263 & R2358_U34); 
assign R2358_U299 = ~(R2358_U13 & R2358_U71); 
assign R2358_U415 = ~(R2358_U13 & R2358_U71); 
assign R2358_U419 = ~(R2358_U13 & R2358_U71); 
assign R2358_U427 = ~(R2358_U227 & R2358_U71); 
assign R2358_U438 = ~(R2358_U134 & R2358_U328); 
assign R2358_U494 = ~(R2358_U84 & R2358_U252); 
assign R2358_U498 = ~(R2358_U382 & R2358_U34); 
assign R2099_U72 = ~(R2099_U311 & R2099_U310); 
assign R2099_U175 = ~R2099_U20; 
assign R2099_U309 = ~(R2099_U49 & R2099_U20); 
assign R2096_U77 = ~(R2096_U154 & R2096_U153); 
assign R2096_U116 = ~R2096_U50; 
assign R2096_U151 = ~(R2096_U50 & REIP_REG_25__SCAN_IN); 
assign ADD_405_U76 = ~(ADD_405_U156 & ADD_405_U155); 
assign ADD_405_U119 = ~ADD_405_U50; 
assign ADD_405_U153 = ~(ADD_405_U50 & INSTADDRPOINTER_REG_25__SCAN_IN); 
assign ADD_515_U77 = ~(ADD_515_U154 & ADD_515_U153); 
assign ADD_515_U116 = ~ADD_515_U50; 
assign ADD_515_U151 = ~(ADD_515_U50 & INSTADDRPOINTER_REG_25__SCAN_IN); 
assign U3462 = ~(U7718 & U7717); 
assign U4551 = ~(U2397 & U4547); 
assign U4552 = ~(U4542 & INSTQUEUE_REG_15__7__SCAN_IN); 
assign U4556 = ~(U2396 & U4547); 
assign U4557 = ~(U4542 & INSTQUEUE_REG_15__6__SCAN_IN); 
assign U4561 = ~(U2395 & U4547); 
assign U4562 = ~(U4542 & INSTQUEUE_REG_15__5__SCAN_IN); 
assign U4566 = ~(U2394 & U4547); 
assign U4567 = ~(U4542 & INSTQUEUE_REG_15__4__SCAN_IN); 
assign U4571 = ~(U2393 & U4547); 
assign U4572 = ~(U4542 & INSTQUEUE_REG_15__3__SCAN_IN); 
assign U4576 = ~(U2392 & U4547); 
assign U4577 = ~(U4542 & INSTQUEUE_REG_15__2__SCAN_IN); 
assign U4581 = ~(U2391 & U4547); 
assign U4582 = ~(U4542 & INSTQUEUE_REG_15__1__SCAN_IN); 
assign U4586 = ~(U2390 & U4547); 
assign U4587 = ~(U4542 & INSTQUEUE_REG_15__0__SCAN_IN); 
assign U4609 = ~(U2397 & U4605); 
assign U4610 = ~(U4600 & INSTQUEUE_REG_14__7__SCAN_IN); 
assign U4614 = ~(U2396 & U4605); 
assign U4615 = ~(U4600 & INSTQUEUE_REG_14__6__SCAN_IN); 
assign U4619 = ~(U2395 & U4605); 
assign U4620 = ~(U4600 & INSTQUEUE_REG_14__5__SCAN_IN); 
assign U4624 = ~(U2394 & U4605); 
assign U4625 = ~(U4600 & INSTQUEUE_REG_14__4__SCAN_IN); 
assign U4629 = ~(U2393 & U4605); 
assign U4630 = ~(U4600 & INSTQUEUE_REG_14__3__SCAN_IN); 
assign U4634 = ~(U2392 & U4605); 
assign U4635 = ~(U4600 & INSTQUEUE_REG_14__2__SCAN_IN); 
assign U4639 = ~(U2391 & U4605); 
assign U4640 = ~(U4600 & INSTQUEUE_REG_14__1__SCAN_IN); 
assign U4644 = ~(U2390 & U4605); 
assign U4645 = ~(U4600 & INSTQUEUE_REG_14__0__SCAN_IN); 
assign U4668 = ~(U2397 & U4664); 
assign U4669 = ~(U4659 & INSTQUEUE_REG_13__7__SCAN_IN); 
assign U4673 = ~(U2396 & U4664); 
assign U4674 = ~(U4659 & INSTQUEUE_REG_13__6__SCAN_IN); 
assign U4678 = ~(U2395 & U4664); 
assign U4679 = ~(U4659 & INSTQUEUE_REG_13__5__SCAN_IN); 
assign U4683 = ~(U2394 & U4664); 
assign U4684 = ~(U4659 & INSTQUEUE_REG_13__4__SCAN_IN); 
assign U4688 = ~(U2393 & U4664); 
assign U4689 = ~(U4659 & INSTQUEUE_REG_13__3__SCAN_IN); 
assign U4693 = ~(U2392 & U4664); 
assign U4694 = ~(U4659 & INSTQUEUE_REG_13__2__SCAN_IN); 
assign U4698 = ~(U2391 & U4664); 
assign U4699 = ~(U4659 & INSTQUEUE_REG_13__1__SCAN_IN); 
assign U4703 = ~(U2390 & U4664); 
assign U4704 = ~(U4659 & INSTQUEUE_REG_13__0__SCAN_IN); 
assign U4725 = ~(U2397 & U4721); 
assign U4726 = ~(U4716 & INSTQUEUE_REG_12__7__SCAN_IN); 
assign U4730 = ~(U2396 & U4721); 
assign U4731 = ~(U4716 & INSTQUEUE_REG_12__6__SCAN_IN); 
assign U4735 = ~(U2395 & U4721); 
assign U4736 = ~(U4716 & INSTQUEUE_REG_12__5__SCAN_IN); 
assign U4740 = ~(U2394 & U4721); 
assign U4741 = ~(U4716 & INSTQUEUE_REG_12__4__SCAN_IN); 
assign U4745 = ~(U2393 & U4721); 
assign U4746 = ~(U4716 & INSTQUEUE_REG_12__3__SCAN_IN); 
assign U4750 = ~(U2392 & U4721); 
assign U4751 = ~(U4716 & INSTQUEUE_REG_12__2__SCAN_IN); 
assign U4755 = ~(U2391 & U4721); 
assign U4756 = ~(U4716 & INSTQUEUE_REG_12__1__SCAN_IN); 
assign U4760 = ~(U2390 & U4721); 
assign U4761 = ~(U4716 & INSTQUEUE_REG_12__0__SCAN_IN); 
assign U4783 = ~(U2397 & U4779); 
assign U4784 = ~(U4774 & INSTQUEUE_REG_11__7__SCAN_IN); 
assign U4788 = ~(U2396 & U4779); 
assign U4789 = ~(U4774 & INSTQUEUE_REG_11__6__SCAN_IN); 
assign U4793 = ~(U2395 & U4779); 
assign U4794 = ~(U4774 & INSTQUEUE_REG_11__5__SCAN_IN); 
assign U4798 = ~(U2394 & U4779); 
assign U4799 = ~(U4774 & INSTQUEUE_REG_11__4__SCAN_IN); 
assign U4803 = ~(U2393 & U4779); 
assign U4804 = ~(U4774 & INSTQUEUE_REG_11__3__SCAN_IN); 
assign U4808 = ~(U2392 & U4779); 
assign U4809 = ~(U4774 & INSTQUEUE_REG_11__2__SCAN_IN); 
assign U4813 = ~(U2391 & U4779); 
assign U4814 = ~(U4774 & INSTQUEUE_REG_11__1__SCAN_IN); 
assign U4818 = ~(U2390 & U4779); 
assign U4819 = ~(U4774 & INSTQUEUE_REG_11__0__SCAN_IN); 
assign U4840 = ~(U2397 & U4836); 
assign U4841 = ~(U4831 & INSTQUEUE_REG_10__7__SCAN_IN); 
assign U4845 = ~(U2396 & U4836); 
assign U4846 = ~(U4831 & INSTQUEUE_REG_10__6__SCAN_IN); 
assign U4850 = ~(U2395 & U4836); 
assign U4851 = ~(U4831 & INSTQUEUE_REG_10__5__SCAN_IN); 
assign U4855 = ~(U2394 & U4836); 
assign U4856 = ~(U4831 & INSTQUEUE_REG_10__4__SCAN_IN); 
assign U4860 = ~(U2393 & U4836); 
assign U4861 = ~(U4831 & INSTQUEUE_REG_10__3__SCAN_IN); 
assign U4865 = ~(U2392 & U4836); 
assign U4866 = ~(U4831 & INSTQUEUE_REG_10__2__SCAN_IN); 
assign U4870 = ~(U2391 & U4836); 
assign U4871 = ~(U4831 & INSTQUEUE_REG_10__1__SCAN_IN); 
assign U4875 = ~(U2390 & U4836); 
assign U4876 = ~(U4831 & INSTQUEUE_REG_10__0__SCAN_IN); 
assign U4898 = ~(U2397 & U4894); 
assign U4899 = ~(U4889 & INSTQUEUE_REG_9__7__SCAN_IN); 
assign U4903 = ~(U2396 & U4894); 
assign U4904 = ~(U4889 & INSTQUEUE_REG_9__6__SCAN_IN); 
assign U4908 = ~(U2395 & U4894); 
assign U4909 = ~(U4889 & INSTQUEUE_REG_9__5__SCAN_IN); 
assign U4913 = ~(U2394 & U4894); 
assign U4914 = ~(U4889 & INSTQUEUE_REG_9__4__SCAN_IN); 
assign U4918 = ~(U2393 & U4894); 
assign U4919 = ~(U4889 & INSTQUEUE_REG_9__3__SCAN_IN); 
assign U4923 = ~(U2392 & U4894); 
assign U4924 = ~(U4889 & INSTQUEUE_REG_9__2__SCAN_IN); 
assign U4928 = ~(U2391 & U4894); 
assign U4929 = ~(U4889 & INSTQUEUE_REG_9__1__SCAN_IN); 
assign U4933 = ~(U2390 & U4894); 
assign U4934 = ~(U4889 & INSTQUEUE_REG_9__0__SCAN_IN); 
assign U4955 = ~(U2397 & U4951); 
assign U4956 = ~(U4946 & INSTQUEUE_REG_8__7__SCAN_IN); 
assign U4960 = ~(U2396 & U4951); 
assign U4961 = ~(U4946 & INSTQUEUE_REG_8__6__SCAN_IN); 
assign U4965 = ~(U2395 & U4951); 
assign U4966 = ~(U4946 & INSTQUEUE_REG_8__5__SCAN_IN); 
assign U4970 = ~(U2394 & U4951); 
assign U4971 = ~(U4946 & INSTQUEUE_REG_8__4__SCAN_IN); 
assign U4975 = ~(U2393 & U4951); 
assign U4976 = ~(U4946 & INSTQUEUE_REG_8__3__SCAN_IN); 
assign U4980 = ~(U2392 & U4951); 
assign U4981 = ~(U4946 & INSTQUEUE_REG_8__2__SCAN_IN); 
assign U4985 = ~(U2391 & U4951); 
assign U4986 = ~(U4946 & INSTQUEUE_REG_8__1__SCAN_IN); 
assign U4990 = ~(U2390 & U4951); 
assign U4991 = ~(U4946 & INSTQUEUE_REG_8__0__SCAN_IN); 
assign U5002 = ~(U4999 & U3647); 
assign U5007 = ~(U5006 & U5005); 
assign U5059 = ~(U5056 & U3656); 
assign U5064 = ~(U5063 & U5062); 
assign U5117 = ~(U5114 & U3665); 
assign U5122 = ~(U5121 & U5120); 
assign U5174 = ~(U5171 & U3674); 
assign U5179 = ~(U5178 & U5177); 
assign U5232 = ~(U5229 & U3683); 
assign U5237 = ~(U5236 & U5235); 
assign U5289 = ~(U5286 & U3692); 
assign U5294 = ~(U5293 & U5292); 
assign U5347 = ~(U5344 & U3701); 
assign U5352 = ~(U5351 & U5350); 
assign U5404 = ~(U5401 & U3710); 
assign U5409 = ~(U5408 & U5407); 
assign U5595 = ~(R2278_U86 & U2377); 
assign U5616 = ~(R2278_U77 & U2377); 
assign U5719 = ~(R2099_U72 & U2380); 
assign U5729 = ~(ADD_405_U76 & U2375); 
assign U5730 = ~(ADD_515_U77 & U2374); 
assign U5813 = ~(U2372 & R2278_U86); 
assign U5815 = ~(R2358_U88 & U2364); 
assign U5828 = ~(U2372 & R2278_U77); 
assign U6158 = ~(U2386 & R2358_U88); 
assign U6268 = ~(U2383 & R2358_U88); 
assign U6323 = ~(U2371 & R2099_U72); 
assign U6399 = ~(U2429 & R2358_U88); 
assign U6523 = ~(U2604 & R2099_U72); 
assign U6531 = ~(R2096_U77 & U7473); 
assign R2278_U25 = ~(R2278_U40 & R2278_U207); 
assign R2278_U37 = ~(R2278_U328 & R2278_U257); 
assign R2278_U56 = R2278_U294 & R2278_U210 & R2278_U298 & R2278_U297; 
assign R2278_U58 = R2278_U332 & R2278_U245; 
assign R2278_U78 = ~(R2278_U197 & R2278_U165); 
assign R2278_U158 = ~(R2278_U27 & R2278_U286); 
assign R2278_U220 = ~R2278_U152; 
assign R2278_U223 = ~(R2278_U55 & R2278_U338); 
assign R2278_U276 = ~(R2278_U221 & R2278_U152); 
assign R2278_U282 = ~R2278_U144; 
assign R2278_U307 = ~R2278_U40; 
assign R2278_U318 = ~(R2278_U317 & R2278_U242); 
assign R2278_U349 = ~(R2278_U188 & R2278_U73); 
assign R2278_U355 = ~(R2278_U196 & R2278_U82); 
assign R2278_U418 = ~(R2278_U285 & R2278_U152); 
assign R2358_U62 = ~(R2358_U438 & R2358_U320); 
assign R2358_U75 = ~(R2358_U74 & R2358_U301); 
assign R2358_U85 = ~(R2358_U494 & R2358_U493); 
assign R2358_U139 = R2358_U415 & R2358_U311; 
assign R2358_U160 = R2358_U299 & R2358_U224 & R2358_U300; 
assign R2358_U217 = ~(R2358_U137 & R2358_U431); 
assign R2358_U256 = ~R2358_U175; 
assign R2358_U261 = ~(R2358_U260 & R2358_U31); 
assign R2358_U266 = ~(R2358_U128 & R2358_U264); 
assign R2358_U292 = ~R2358_U63; 
assign R2358_U306 = ~R2358_U74; 
assign R2358_U369 = ~(R2358_U300 & R2358_U299); 
assign R2358_U402 = ~(R2358_U63 & R2358_U277); 
assign R2358_U410 = ~(R2358_U223 & R2358_U224 & R2358_U299); 
assign R2358_U411 = ~(R2358_U309 & R2358_U311 & R2358_U224 & R2358_U299); 
assign R2358_U418 = ~R2358_U66; 
assign R2358_U420 = ~(R2358_U427 & R2358_U419 & R2358_U428); 
assign R2358_U422 = ~(R2358_U66 & R2358_U7); 
assign R2358_U430 = ~(R2358_U12 & R2358_U66); 
assign R2358_U491 = ~(R2358_U165 & R2358_U175); 
assign R2358_U499 = ~(R2358_U497 & R2358_U260); 
assign R2099_U21 = ~(R2099_U175 & R2099_U49); 
assign R2099_U308 = ~(R2099_U240 & R2099_U175); 
assign R2096_U52 = ~(R2096_U116 & REIP_REG_25__SCAN_IN); 
assign R2096_U152 = ~(R2096_U116 & R2096_U51); 
assign ADD_405_U52 = ~(ADD_405_U119 & INSTADDRPOINTER_REG_25__SCAN_IN); 
assign ADD_405_U154 = ~(ADD_405_U119 & ADD_405_U51); 
assign ADD_515_U52 = ~(ADD_515_U116 & INSTADDRPOINTER_REG_25__SCAN_IN); 
assign ADD_515_U152 = ~(ADD_515_U116 & ADD_515_U51); 
assign U2854 = ~(U6269 & U6270 & U6268); 
assign U2886 = ~(U6159 & U6157 & U6158); 
assign U2981 = ~(U5814 & U5812 & U5813 & U5816 & U5815); 
assign U3010 = ~(U3778 & U3780 & U5616); 
assign U3013 = ~(U3769 & U3771 & U5595); 
assign U3084 = ~(U4991 & U4990 & U3646); 
assign U3085 = ~(U4986 & U4985 & U3645); 
assign U3086 = ~(U4981 & U4980 & U3644); 
assign U3087 = ~(U4976 & U4975 & U3643); 
assign U3088 = ~(U4971 & U4970 & U3642); 
assign U3089 = ~(U4966 & U4965 & U3641); 
assign U3090 = ~(U4961 & U4960 & U3640); 
assign U3091 = ~(U4956 & U4955 & U3639); 
assign U3092 = ~(U4934 & U4933 & U3637); 
assign U3093 = ~(U4929 & U4928 & U3636); 
assign U3094 = ~(U4924 & U4923 & U3635); 
assign U3095 = ~(U4919 & U4918 & U3634); 
assign U3096 = ~(U4914 & U4913 & U3633); 
assign U3097 = ~(U4909 & U4908 & U3632); 
assign U3098 = ~(U4904 & U4903 & U3631); 
assign U3099 = ~(U4899 & U4898 & U3630); 
assign U3100 = ~(U4876 & U4875 & U3628); 
assign U3101 = ~(U4871 & U4870 & U3627); 
assign U3102 = ~(U4866 & U4865 & U3626); 
assign U3103 = ~(U4861 & U4860 & U3625); 
assign U3104 = ~(U4856 & U4855 & U3624); 
assign U3105 = ~(U4851 & U4850 & U3623); 
assign U3106 = ~(U4846 & U4845 & U3622); 
assign U3107 = ~(U4841 & U4840 & U3621); 
assign U3108 = ~(U4819 & U4818 & U3619); 
assign U3109 = ~(U4814 & U4813 & U3618); 
assign U3110 = ~(U4809 & U4808 & U3617); 
assign U3111 = ~(U4804 & U4803 & U3616); 
assign U3112 = ~(U4799 & U4798 & U3615); 
assign U3113 = ~(U4794 & U4793 & U3614); 
assign U3114 = ~(U4789 & U4788 & U3613); 
assign U3115 = ~(U4784 & U4783 & U3612); 
assign U3116 = ~(U4761 & U4760 & U3610); 
assign U3117 = ~(U4756 & U4755 & U3609); 
assign U3118 = ~(U4751 & U4750 & U3608); 
assign U3119 = ~(U4746 & U4745 & U3607); 
assign U3120 = ~(U4741 & U4740 & U3606); 
assign U3121 = ~(U4736 & U4735 & U3605); 
assign U3122 = ~(U4731 & U4730 & U3604); 
assign U3123 = ~(U4726 & U4725 & U3603); 
assign U3124 = ~(U4704 & U4703 & U3601); 
assign U3125 = ~(U4699 & U4698 & U3600); 
assign U3126 = ~(U4694 & U4693 & U3599); 
assign U3127 = ~(U4689 & U4688 & U3598); 
assign U3128 = ~(U4684 & U4683 & U3597); 
assign U3129 = ~(U4679 & U4678 & U3596); 
assign U3130 = ~(U4674 & U4673 & U3595); 
assign U3131 = ~(U4669 & U4668 & U3594); 
assign U3132 = ~(U4645 & U4644 & U3592); 
assign U3133 = ~(U4640 & U4639 & U3591); 
assign U3134 = ~(U4635 & U4634 & U3590); 
assign U3135 = ~(U4630 & U4629 & U3589); 
assign U3136 = ~(U4625 & U4624 & U3588); 
assign U3137 = ~(U4620 & U4619 & U3587); 
assign U3138 = ~(U4615 & U4614 & U3586); 
assign U3139 = ~(U4610 & U4609 & U3585); 
assign U3140 = ~(U4587 & U4586 & U3583); 
assign U3141 = ~(U4582 & U4581 & U3582); 
assign U3142 = ~(U4577 & U4576 & U3581); 
assign U3143 = ~(U4572 & U4571 & U3580); 
assign U3144 = ~(U4567 & U4566 & U3579); 
assign U3145 = ~(U4562 & U4561 & U3578); 
assign U3146 = ~(U4557 & U4556 & U3577); 
assign U3147 = ~(U4552 & U4551 & U3576); 
assign U3826 = U5727 & U5729; 
assign U3828 = U3827 & U5730; 
assign U3885 = U6401 & U6400 & U6403 & U6402 & U6399; 
assign U3922 = U6533 & U6531; 
assign U5011 = ~(U2397 & U5007); 
assign U5012 = ~(U5002 & INSTQUEUE_REG_7__7__SCAN_IN); 
assign U5016 = ~(U2396 & U5007); 
assign U5017 = ~(U5002 & INSTQUEUE_REG_7__6__SCAN_IN); 
assign U5021 = ~(U2395 & U5007); 
assign U5022 = ~(U5002 & INSTQUEUE_REG_7__5__SCAN_IN); 
assign U5026 = ~(U2394 & U5007); 
assign U5027 = ~(U5002 & INSTQUEUE_REG_7__4__SCAN_IN); 
assign U5031 = ~(U2393 & U5007); 
assign U5032 = ~(U5002 & INSTQUEUE_REG_7__3__SCAN_IN); 
assign U5036 = ~(U2392 & U5007); 
assign U5037 = ~(U5002 & INSTQUEUE_REG_7__2__SCAN_IN); 
assign U5041 = ~(U2391 & U5007); 
assign U5042 = ~(U5002 & INSTQUEUE_REG_7__1__SCAN_IN); 
assign U5046 = ~(U2390 & U5007); 
assign U5047 = ~(U5002 & INSTQUEUE_REG_7__0__SCAN_IN); 
assign U5068 = ~(U2397 & U5064); 
assign U5069 = ~(U5059 & INSTQUEUE_REG_6__7__SCAN_IN); 
assign U5073 = ~(U2396 & U5064); 
assign U5074 = ~(U5059 & INSTQUEUE_REG_6__6__SCAN_IN); 
assign U5078 = ~(U2395 & U5064); 
assign U5079 = ~(U5059 & INSTQUEUE_REG_6__5__SCAN_IN); 
assign U5083 = ~(U2394 & U5064); 
assign U5084 = ~(U5059 & INSTQUEUE_REG_6__4__SCAN_IN); 
assign U5088 = ~(U2393 & U5064); 
assign U5089 = ~(U5059 & INSTQUEUE_REG_6__3__SCAN_IN); 
assign U5093 = ~(U2392 & U5064); 
assign U5094 = ~(U5059 & INSTQUEUE_REG_6__2__SCAN_IN); 
assign U5098 = ~(U2391 & U5064); 
assign U5099 = ~(U5059 & INSTQUEUE_REG_6__1__SCAN_IN); 
assign U5103 = ~(U2390 & U5064); 
assign U5104 = ~(U5059 & INSTQUEUE_REG_6__0__SCAN_IN); 
assign U5126 = ~(U2397 & U5122); 
assign U5127 = ~(U5117 & INSTQUEUE_REG_5__7__SCAN_IN); 
assign U5131 = ~(U2396 & U5122); 
assign U5132 = ~(U5117 & INSTQUEUE_REG_5__6__SCAN_IN); 
assign U5136 = ~(U2395 & U5122); 
assign U5137 = ~(U5117 & INSTQUEUE_REG_5__5__SCAN_IN); 
assign U5141 = ~(U2394 & U5122); 
assign U5142 = ~(U5117 & INSTQUEUE_REG_5__4__SCAN_IN); 
assign U5146 = ~(U2393 & U5122); 
assign U5147 = ~(U5117 & INSTQUEUE_REG_5__3__SCAN_IN); 
assign U5151 = ~(U2392 & U5122); 
assign U5152 = ~(U5117 & INSTQUEUE_REG_5__2__SCAN_IN); 
assign U5156 = ~(U2391 & U5122); 
assign U5157 = ~(U5117 & INSTQUEUE_REG_5__1__SCAN_IN); 
assign U5161 = ~(U2390 & U5122); 
assign U5162 = ~(U5117 & INSTQUEUE_REG_5__0__SCAN_IN); 
assign U5183 = ~(U2397 & U5179); 
assign U5184 = ~(U5174 & INSTQUEUE_REG_4__7__SCAN_IN); 
assign U5188 = ~(U2396 & U5179); 
assign U5189 = ~(U5174 & INSTQUEUE_REG_4__6__SCAN_IN); 
assign U5193 = ~(U2395 & U5179); 
assign U5194 = ~(U5174 & INSTQUEUE_REG_4__5__SCAN_IN); 
assign U5198 = ~(U2394 & U5179); 
assign U5199 = ~(U5174 & INSTQUEUE_REG_4__4__SCAN_IN); 
assign U5203 = ~(U2393 & U5179); 
assign U5204 = ~(U5174 & INSTQUEUE_REG_4__3__SCAN_IN); 
assign U5208 = ~(U2392 & U5179); 
assign U5209 = ~(U5174 & INSTQUEUE_REG_4__2__SCAN_IN); 
assign U5213 = ~(U2391 & U5179); 
assign U5214 = ~(U5174 & INSTQUEUE_REG_4__1__SCAN_IN); 
assign U5218 = ~(U2390 & U5179); 
assign U5219 = ~(U5174 & INSTQUEUE_REG_4__0__SCAN_IN); 
assign U5241 = ~(U2397 & U5237); 
assign U5242 = ~(U5232 & INSTQUEUE_REG_3__7__SCAN_IN); 
assign U5246 = ~(U2396 & U5237); 
assign U5247 = ~(U5232 & INSTQUEUE_REG_3__6__SCAN_IN); 
assign U5251 = ~(U2395 & U5237); 
assign U5252 = ~(U5232 & INSTQUEUE_REG_3__5__SCAN_IN); 
assign U5256 = ~(U2394 & U5237); 
assign U5257 = ~(U5232 & INSTQUEUE_REG_3__4__SCAN_IN); 
assign U5261 = ~(U2393 & U5237); 
assign U5262 = ~(U5232 & INSTQUEUE_REG_3__3__SCAN_IN); 
assign U5266 = ~(U2392 & U5237); 
assign U5267 = ~(U5232 & INSTQUEUE_REG_3__2__SCAN_IN); 
assign U5271 = ~(U2391 & U5237); 
assign U5272 = ~(U5232 & INSTQUEUE_REG_3__1__SCAN_IN); 
assign U5276 = ~(U2390 & U5237); 
assign U5277 = ~(U5232 & INSTQUEUE_REG_3__0__SCAN_IN); 
assign U5298 = ~(U2397 & U5294); 
assign U5299 = ~(U5289 & INSTQUEUE_REG_2__7__SCAN_IN); 
assign U5303 = ~(U2396 & U5294); 
assign U5304 = ~(U5289 & INSTQUEUE_REG_2__6__SCAN_IN); 
assign U5308 = ~(U2395 & U5294); 
assign U5309 = ~(U5289 & INSTQUEUE_REG_2__5__SCAN_IN); 
assign U5313 = ~(U2394 & U5294); 
assign U5314 = ~(U5289 & INSTQUEUE_REG_2__4__SCAN_IN); 
assign U5318 = ~(U2393 & U5294); 
assign U5319 = ~(U5289 & INSTQUEUE_REG_2__3__SCAN_IN); 
assign U5323 = ~(U2392 & U5294); 
assign U5324 = ~(U5289 & INSTQUEUE_REG_2__2__SCAN_IN); 
assign U5328 = ~(U2391 & U5294); 
assign U5329 = ~(U5289 & INSTQUEUE_REG_2__1__SCAN_IN); 
assign U5333 = ~(U2390 & U5294); 
assign U5334 = ~(U5289 & INSTQUEUE_REG_2__0__SCAN_IN); 
assign U5356 = ~(U2397 & U5352); 
assign U5357 = ~(U5347 & INSTQUEUE_REG_1__7__SCAN_IN); 
assign U5361 = ~(U2396 & U5352); 
assign U5362 = ~(U5347 & INSTQUEUE_REG_1__6__SCAN_IN); 
assign U5366 = ~(U2395 & U5352); 
assign U5367 = ~(U5347 & INSTQUEUE_REG_1__5__SCAN_IN); 
assign U5371 = ~(U2394 & U5352); 
assign U5372 = ~(U5347 & INSTQUEUE_REG_1__4__SCAN_IN); 
assign U5376 = ~(U2393 & U5352); 
assign U5377 = ~(U5347 & INSTQUEUE_REG_1__3__SCAN_IN); 
assign U5381 = ~(U2392 & U5352); 
assign U5382 = ~(U5347 & INSTQUEUE_REG_1__2__SCAN_IN); 
assign U5386 = ~(U2391 & U5352); 
assign U5387 = ~(U5347 & INSTQUEUE_REG_1__1__SCAN_IN); 
assign U5391 = ~(U2390 & U5352); 
assign U5392 = ~(U5347 & INSTQUEUE_REG_1__0__SCAN_IN); 
assign U5413 = ~(U2397 & U5409); 
assign U5414 = ~(U5404 & INSTQUEUE_REG_0__7__SCAN_IN); 
assign U5418 = ~(U2396 & U5409); 
assign U5419 = ~(U5404 & INSTQUEUE_REG_0__6__SCAN_IN); 
assign U5423 = ~(U2395 & U5409); 
assign U5424 = ~(U5404 & INSTQUEUE_REG_0__5__SCAN_IN); 
assign U5428 = ~(U2394 & U5409); 
assign U5432 = ~(U2393 & U5409); 
assign U5433 = ~(U5404 & INSTQUEUE_REG_0__3__SCAN_IN); 
assign U5437 = ~(U2392 & U5409); 
assign U5438 = ~(U5404 & INSTQUEUE_REG_0__2__SCAN_IN); 
assign U5442 = ~(U2391 & U5409); 
assign U5443 = ~(U5404 & INSTQUEUE_REG_0__1__SCAN_IN); 
assign U5447 = ~(U2390 & U5409); 
assign U5448 = ~(U5404 & INSTQUEUE_REG_0__0__SCAN_IN); 
assign U5830 = ~(R2358_U85 & U2364); 
assign U6167 = ~(U2386 & R2358_U85); 
assign U6277 = ~(U2383 & R2358_U85); 
assign U6422 = ~(U2367 & R2358_U85); 
assign U7600 = ~(U5404 & INSTQUEUE_REG_0__4__SCAN_IN); 
assign R2278_U66 = R2278_U25 & R2278_U23; 
assign R2278_U67 = R2278_U318 & R2278_U243; 
assign R2278_U74 = R2278_U350 & R2278_U349; 
assign R2278_U83 = R2278_U356 & R2278_U355; 
assign R2278_U140 = ~(R2278_U223 & R2278_U56); 
assign R2278_U149 = ~(R2278_U29 & R2278_U276); 
assign R2278_U198 = ~R2278_U78; 
assign R2278_U287 = ~R2278_U158; 
assign R2278_U288 = ~(R2278_U158 & R2278_U217); 
assign R2278_U308 = ~R2278_U25; 
assign R2278_U319 = ~(R2278_U318 & R2278_U243); 
assign R2278_U329 = ~R2278_U37; 
assign R2278_U331 = ~(R2278_U37 & R2278_U259); 
assign R2278_U354 = ~(R2278_U199 & R2278_U78); 
assign R2278_U417 = ~(R2278_U220 & R2278_U153); 
assign R2278_U422 = ~(R2278_U291 & R2278_U158); 
assign R2358_U86 = ~(R2358_U499 & R2358_U498); 
assign R2358_U140 = R2358_U420 & R2358_U411; 
assign R2358_U144 = R2358_U402 & R2358_U278; 
assign R2358_U146 = R2358_U420 & R2358_U411; 
assign R2358_U157 = R2358_U418 & R2358_U46; 
assign R2358_U161 = R2358_U369 & R2358_U227; 
assign R2358_U219 = ~(R2358_U138 & R2358_U217 & R2358_U139); 
assign R2358_U262 = ~(R2358_U127 & R2358_U261); 
assign R2358_U308 = ~R2358_U217; 
assign R2358_U361 = ~(R2358_U310 & R2358_U217); 
assign R2358_U372 = ~R2358_U75; 
assign R2358_U373 = ~(R2358_U75 & R2358_U307); 
assign R2358_U376 = ~(R2358_U163 & R2358_U75); 
assign R2358_U378 = ~(R2358_U306 & R2358_U377); 
assign R2358_U406 = ~(R2358_U8 & R2358_U62); 
assign R2358_U434 = ~(R2358_U418 & R2358_U55); 
assign R2358_U439 = ~R2358_U62; 
assign R2358_U492 = ~(R2358_U256 & R2358_U447); 
assign R2358_U651 = ~(R2358_U401 & R2358_U217); 
assign R2099_U71 = ~(R2099_U309 & R2099_U308); 
assign R2099_U176 = ~R2099_U21; 
assign R2099_U307 = ~(R2099_U48 & R2099_U21); 
assign R2096_U76 = ~(R2096_U152 & R2096_U151); 
assign R2096_U117 = ~R2096_U52; 
assign R2096_U149 = ~(R2096_U52 & REIP_REG_26__SCAN_IN); 
assign ADD_405_U75 = ~(ADD_405_U154 & ADD_405_U153); 
assign ADD_405_U120 = ~ADD_405_U52; 
assign ADD_405_U151 = ~(ADD_405_U52 & INSTADDRPOINTER_REG_26__SCAN_IN); 
assign ADD_515_U76 = ~(ADD_515_U152 & ADD_515_U151); 
assign ADD_515_U117 = ~ADD_515_U52; 
assign ADD_515_U149 = ~(ADD_515_U52 & INSTADDRPOINTER_REG_26__SCAN_IN); 
assign U2819 = ~(U3891 & U6420 & U3890 & U6419 & U6422); 
assign U2822 = ~(U3884 & U6397 & U6398 & U3885); 
assign U2851 = ~(U6278 & U6279 & U6277); 
assign U2883 = ~(U6168 & U6166 & U6167); 
assign U2978 = ~(U5829 & U5827 & U5831 & U5828 & U5830); 
assign U3020 = ~(U5448 & U5447 & U3718); 
assign U3021 = ~(U5443 & U5442 & U3717); 
assign U3022 = ~(U5438 & U5437 & U3716); 
assign U3023 = ~(U5433 & U5432 & U3715); 
assign U3024 = ~(U7600 & U5428 & U3714); 
assign U3025 = ~(U5424 & U5423 & U3713); 
assign U3026 = ~(U5419 & U5418 & U3712); 
assign U3027 = ~(U5414 & U5413 & U3711); 
assign U3028 = ~(U5392 & U5391 & U3709); 
assign U3029 = ~(U5387 & U5386 & U3708); 
assign U3030 = ~(U5382 & U5381 & U3707); 
assign U3031 = ~(U5377 & U5376 & U3706); 
assign U3032 = ~(U5372 & U5371 & U3705); 
assign U3033 = ~(U5367 & U5366 & U3704); 
assign U3034 = ~(U5362 & U5361 & U3703); 
assign U3035 = ~(U5357 & U5356 & U3702); 
assign U3036 = ~(U5334 & U5333 & U3700); 
assign U3037 = ~(U5329 & U5328 & U3699); 
assign U3038 = ~(U5324 & U5323 & U3698); 
assign U3039 = ~(U5319 & U5318 & U3697); 
assign U3040 = ~(U5314 & U5313 & U3696); 
assign U3041 = ~(U5309 & U5308 & U3695); 
assign U3042 = ~(U5304 & U5303 & U3694); 
assign U3043 = ~(U5299 & U5298 & U3693); 
assign U3044 = ~(U5277 & U5276 & U3691); 
assign U3045 = ~(U5272 & U5271 & U3690); 
assign U3046 = ~(U5267 & U5266 & U3689); 
assign U3047 = ~(U5262 & U5261 & U3688); 
assign U3048 = ~(U5257 & U5256 & U3687); 
assign U3049 = ~(U5252 & U5251 & U3686); 
assign U3050 = ~(U5247 & U5246 & U3685); 
assign U3051 = ~(U5242 & U5241 & U3684); 
assign U3052 = ~(U5219 & U5218 & U3682); 
assign U3053 = ~(U5214 & U5213 & U3681); 
assign U3054 = ~(U5209 & U5208 & U3680); 
assign U3055 = ~(U5204 & U5203 & U3679); 
assign U3056 = ~(U5199 & U5198 & U3678); 
assign U3057 = ~(U5194 & U5193 & U3677); 
assign U3058 = ~(U5189 & U5188 & U3676); 
assign U3059 = ~(U5184 & U5183 & U3675); 
assign U3060 = ~(U5162 & U5161 & U3673); 
assign U3061 = ~(U5157 & U5156 & U3672); 
assign U3062 = ~(U5152 & U5151 & U3671); 
assign U3063 = ~(U5147 & U5146 & U3670); 
assign U3064 = ~(U5142 & U5141 & U3669); 
assign U3065 = ~(U5137 & U5136 & U3668); 
assign U3066 = ~(U5132 & U5131 & U3667); 
assign U3067 = ~(U5127 & U5126 & U3666); 
assign U3068 = ~(U5104 & U5103 & U3664); 
assign U3069 = ~(U5099 & U5098 & U3663); 
assign U3070 = ~(U5094 & U5093 & U3662); 
assign U3071 = ~(U5089 & U5088 & U3661); 
assign U3072 = ~(U5084 & U5083 & U3660); 
assign U3073 = ~(U5079 & U5078 & U3659); 
assign U3074 = ~(U5074 & U5073 & U3658); 
assign U3075 = ~(U5069 & U5068 & U3657); 
assign U3076 = ~(U5047 & U5046 & U3655); 
assign U3077 = ~(U5042 & U5041 & U3654); 
assign U3078 = ~(U5037 & U5036 & U3653); 
assign U3079 = ~(U5032 & U5031 & U3652); 
assign U3080 = ~(U5027 & U5026 & U3651); 
assign U3081 = ~(U5022 & U5021 & U3650); 
assign U3082 = ~(U5017 & U5016 & U3649); 
assign U3083 = ~(U5012 & U5011 & U3648); 
assign U5602 = ~(R2278_U83 & U2377); 
assign U5623 = ~(R2278_U74 & U2377); 
assign U5726 = ~(R2099_U71 & U2380); 
assign U5736 = ~(ADD_405_U75 & U2375); 
assign U5737 = ~(ADD_515_U76 & U2374); 
assign U5818 = ~(U2372 & R2278_U83); 
assign U5820 = ~(R2358_U86 & U2364); 
assign U5833 = ~(U2372 & R2278_U74); 
assign U6161 = ~(U2386 & R2358_U86); 
assign U6271 = ~(U2383 & R2358_U86); 
assign U6326 = ~(U2371 & R2099_U71); 
assign U6408 = ~(U2367 & R2358_U86); 
assign U6530 = ~(U2604 & R2099_U71); 
assign U6538 = ~(R2096_U76 & U7473); 
assign R2278_U61 = R2278_U331 & R2278_U260; 
assign R2278_U154 = R2278_U418 & R2278_U417; 
assign R2278_U155 = ~(R2278_U288 & R2278_U28); 
assign R2278_U224 = ~R2278_U140; 
assign R2278_U277 = ~R2278_U149; 
assign R2278_U278 = ~(R2278_U149 & R2278_U213); 
assign R2278_U320 = ~(R2278_U319 & R2278_U204); 
assign R2278_U333 = ~(R2278_U308 & R2278_U13); 
assign R2278_U339 = ~(R2278_U225 & R2278_U140); 
assign R2278_U341 = ~(R2278_U6 & R2278_U140); 
assign R2278_U343 = ~(R2278_U7 & R2278_U140); 
assign R2278_U345 = ~(R2278_U8 & R2278_U140); 
assign R2278_U347 = ~(R2278_U57 & R2278_U140); 
assign R2278_U353 = ~(R2278_U198 & R2278_U79); 
assign R2278_U410 = ~(R2278_U275 & R2278_U140); 
assign R2278_U416 = ~(R2278_U284 & R2278_U149); 
assign R2278_U421 = ~(R2278_U287 & R2278_U159); 
assign R2358_U21 = R2358_U266 & R2358_U262; 
assign R2358_U67 = ~(R2358_U410 & R2358_U219 & R2358_U146); 
assign R2358_U83 = ~(R2358_U492 & R2358_U491); 
assign R2358_U145 = R2358_U144 & R2358_U406 & R2358_U430; 
assign R2358_U150 = R2358_U422 & R2358_U439; 
assign R2358_U155 = R2358_U156 & R2358_U434; 
assign R2358_U216 = ~(R2358_U53 & R2358_U361); 
assign R2358_U374 = ~(R2358_U162 & R2358_U373); 
assign R2358_U379 = ~(R2358_U372 & R2358_U307); 
assign R2358_U435 = ~(R2358_U410 & R2358_U219 & R2358_U140); 
assign R2358_U652 = ~(R2358_U121 & R2358_U308); 
assign R2099_U22 = ~(R2099_U176 & R2099_U48); 
assign R2099_U306 = ~(R2099_U237 & R2099_U176); 
assign R2096_U54 = ~(R2096_U117 & REIP_REG_26__SCAN_IN); 
assign R2096_U150 = ~(R2096_U117 & R2096_U53); 
assign ADD_405_U54 = ~(ADD_405_U120 & INSTADDRPOINTER_REG_26__SCAN_IN); 
assign ADD_405_U152 = ~(ADD_405_U120 & ADD_405_U53); 
assign ADD_515_U54 = ~(ADD_515_U117 & INSTADDRPOINTER_REG_26__SCAN_IN); 
assign ADD_515_U150 = ~(ADD_515_U117 & ADD_515_U53); 
assign U2821 = ~(U3887 & U6406 & U3886 & U6405 & U6408); 
assign U2853 = ~(U6272 & U6273 & U6271); 
assign U2885 = ~(U6162 & U6160 & U6161); 
assign U2980 = ~(U5819 & U5817 & U5818 & U5821 & U5820); 
assign U3009 = ~(U3781 & U3783 & U5623); 
assign U3012 = ~(U3772 & U3774 & U5602); 
assign U3829 = U5734 & U5736; 
assign U3831 = U3830 & U5737; 
assign U3924 = U6540 & U6538; 
assign U5644 = ~(R2278_U154 & U2377); 
assign U5825 = ~(R2358_U21 & U2364); 
assign U5835 = ~(R2358_U83 & U2364); 
assign U5848 = ~(U2372 & R2278_U154); 
assign U6164 = ~(U2386 & R2358_U21); 
assign U6170 = ~(U2386 & R2358_U83); 
assign U6274 = ~(U2383 & R2358_U21); 
assign U6280 = ~(U2383 & R2358_U83); 
assign U6415 = ~(U2367 & R2358_U21); 
assign U6429 = ~(U2367 & R2358_U83); 
assign R2278_U59 = R2278_U333 & R2278_U320 & R2278_U58; 
assign R2278_U80 = R2278_U354 & R2278_U353; 
assign R2278_U128 = ~(R2278_U66 & R2278_U345); 
assign R2278_U132 = ~(R2278_U307 & R2278_U343); 
assign R2278_U135 = ~(R2278_U305 & R2278_U341); 
assign R2278_U138 = ~(R2278_U339 & R2278_U24); 
assign R2278_U146 = ~(R2278_U31 & R2278_U278); 
assign R2278_U160 = R2278_U422 & R2278_U421; 
assign R2278_U289 = ~R2278_U155; 
assign R2278_U409 = ~(R2278_U224 & R2278_U141); 
assign R2278_U415 = ~(R2278_U277 & R2278_U150); 
assign R2278_U420 = ~(R2278_U290 & R2278_U155); 
assign R2358_U14 = R2358_U379 & R2358_U378; 
assign R2358_U15 = R2358_U376 & R2358_U374; 
assign R2358_U70 = ~(R2358_U313 & R2358_U67); 
assign R2358_U122 = ~(R2358_U652 & R2358_U651); 
assign R2358_U312 = ~R2358_U67; 
assign R2358_U362 = ~R2358_U216; 
assign R2358_U364 = ~(R2358_U363 & R2358_U216); 
assign R2358_U409 = ~(R2358_U159 & R2358_U67); 
assign R2358_U416 = ~(R2358_U426 & R2358_U67); 
assign R2358_U421 = ~(R2358_U67 & R2358_U148); 
assign R2358_U429 = ~(R2358_U143 & R2358_U435); 
assign R2358_U649 = ~(R2358_U400 & R2358_U216); 
assign R2099_U70 = ~(R2099_U307 & R2099_U306); 
assign R2099_U177 = ~R2099_U22; 
assign R2099_U305 = ~(R2099_U47 & R2099_U22); 
assign R2096_U75 = ~(R2096_U150 & R2096_U149); 
assign R2096_U118 = ~R2096_U54; 
assign R2096_U147 = ~(R2096_U54 & REIP_REG_27__SCAN_IN); 
assign ADD_405_U74 = ~(ADD_405_U152 & ADD_405_U151); 
assign ADD_405_U121 = ~ADD_405_U54; 
assign ADD_405_U149 = ~(ADD_405_U54 & INSTADDRPOINTER_REG_27__SCAN_IN); 
assign ADD_515_U75 = ~(ADD_515_U150 & ADD_515_U149); 
assign ADD_515_U118 = ~ADD_515_U54; 
assign ADD_515_U147 = ~(ADD_515_U54 & INSTADDRPOINTER_REG_27__SCAN_IN); 
assign U2818 = ~(U3893 & U6427 & U3892 & U6426 & U6429); 
assign U2820 = ~(U3889 & U6413 & U3888 & U6412 & U6415); 
assign U2850 = ~(U6281 & U6282 & U6280); 
assign U2852 = ~(U6275 & U6276 & U6274); 
assign U2882 = ~(U6171 & U6169 & U6170); 
assign U2884 = ~(U6165 & U6163 & U6164); 
assign U2977 = ~(U5834 & U5832 & U5836 & U5833 & U5835); 
assign U3006 = ~(U3790 & U3792 & U5644); 
assign U5609 = ~(R2278_U80 & U2377); 
assign U5630 = ~(R2278_U160 & U2377); 
assign U5733 = ~(R2099_U70 & U2380); 
assign U5743 = ~(ADD_405_U74 & U2375); 
assign U5744 = ~(ADD_515_U75 & U2374); 
assign U5823 = ~(U2372 & R2278_U80); 
assign U5838 = ~(U2372 & R2278_U160); 
assign U5840 = ~(R2358_U14 & U2364); 
assign U5845 = ~(R2358_U15 & U2364); 
assign U5850 = ~(R2358_U122 & U2364); 
assign U6173 = ~(U2386 & R2358_U14); 
assign U6176 = ~(U2386 & R2358_U15); 
assign U6179 = ~(U2386 & R2358_U122); 
assign U6283 = ~(U2383 & R2358_U14); 
assign U6286 = ~(U2383 & R2358_U15); 
assign U6289 = ~(U2383 & R2358_U122); 
assign U6329 = ~(U2371 & R2099_U70); 
assign U6436 = ~(U2367 & R2358_U14); 
assign U6443 = ~(U2367 & R2358_U15); 
assign U6450 = ~(U2367 & R2358_U122); 
assign U6537 = ~(U2604 & R2099_U70); 
assign U6545 = ~(R2096_U75 & U7473); 
assign R2278_U110 = ~(R2278_U59 & R2278_U347); 
assign R2278_U142 = R2278_U410 & R2278_U409; 
assign R2278_U151 = R2278_U416 & R2278_U415; 
assign R2278_U233 = ~(R2278_U231 & R2278_U128); 
assign R2278_U279 = ~R2278_U146; 
assign R2278_U280 = ~(R2278_U146 & R2278_U211); 
assign R2278_U309 = ~(R2278_U9 & R2278_U128); 
assign R2278_U311 = ~(R2278_U10 & R2278_U128); 
assign R2278_U313 = ~(R2278_U11 & R2278_U128); 
assign R2278_U316 = ~(R2278_U12 & R2278_U128); 
assign R2278_U340 = ~R2278_U138; 
assign R2278_U342 = ~R2278_U135; 
assign R2278_U344 = ~R2278_U132; 
assign R2278_U346 = ~R2278_U128; 
assign R2278_U399 = ~(R2278_U270 & R2278_U128); 
assign R2278_U403 = ~(R2278_U272 & R2278_U132); 
assign R2278_U405 = ~(R2278_U273 & R2278_U135); 
assign R2278_U407 = ~(R2278_U274 & R2278_U138); 
assign R2278_U414 = ~(R2278_U283 & R2278_U146); 
assign R2278_U419 = ~(R2278_U289 & R2278_U156); 
assign R2358_U68 = ~(R2358_U418 & R2358_U416); 
assign R2358_U72 = ~(R2358_U51 & R2358_U364); 
assign R2358_U202 = ~(R2358_U145 & R2358_U429); 
assign R2358_U208 = ~(R2358_U150 & R2358_U421); 
assign R2358_U213 = ~(R2358_U412 & R2358_U409); 
assign R2358_U215 = ~(R2358_U61 & R2358_U70); 
assign R2358_U314 = ~R2358_U70; 
assign R2358_U349 = ~(R2358_U157 & R2358_U416); 
assign R2358_U359 = ~(R2358_U312 & R2358_U358); 
assign R2358_U433 = ~(R2358_U312 & R2358_U418); 
assign R2358_U650 = ~(R2358_U362 & R2358_U648); 
assign R2099_U23 = ~(R2099_U177 & R2099_U47); 
assign R2099_U304 = ~(R2099_U234 & R2099_U177); 
assign R2096_U56 = ~(R2096_U118 & REIP_REG_27__SCAN_IN); 
assign R2096_U148 = ~(R2096_U118 & R2096_U55); 
assign ADD_405_U56 = ~(ADD_405_U121 & INSTADDRPOINTER_REG_27__SCAN_IN); 
assign ADD_405_U150 = ~(ADD_405_U121 & ADD_405_U55); 
assign ADD_515_U56 = ~(ADD_515_U118 & INSTADDRPOINTER_REG_27__SCAN_IN); 
assign ADD_515_U148 = ~(ADD_515_U118 & ADD_515_U55); 
assign U2815 = ~(U3899 & U6448 & U3898 & U6447 & U6450); 
assign U2816 = ~(U3897 & U6441 & U3896 & U6440 & U6443); 
assign U2817 = ~(U3895 & U6434 & U3894 & U6433 & U6436); 
assign U2847 = ~(U6290 & U6291 & U6289); 
assign U2848 = ~(U6287 & U6288 & U6286); 
assign U2849 = ~(U6284 & U6285 & U6283); 
assign U2879 = ~(U6180 & U6178 & U6179); 
assign U2880 = ~(U6177 & U6175 & U6176); 
assign U2881 = ~(U6174 & U6172 & U6173); 
assign U2974 = ~(U5849 & U5847 & U5851 & U5848 & U5850); 
assign U2976 = ~(U5839 & U5837 & U5841 & U5838 & U5840); 
assign U2979 = ~(U5824 & U5822 & U5823 & U5826 & U5825); 
assign U3008 = ~(U3784 & U3786 & U5630); 
assign U3011 = ~(U3775 & U3777 & U5609); 
assign U3832 = U5741 & U5743; 
assign U3834 = U3833 & U5744; 
assign U3926 = U6547 & U6545; 
assign U5651 = ~(R2278_U151 & U2377); 
assign U5672 = ~(R2278_U142 & U2377); 
assign U5853 = ~(U2372 & R2278_U151); 
assign U5868 = ~(U2372 & R2278_U142); 
assign R2278_U112 = ~(R2278_U67 & R2278_U316); 
assign R2278_U115 = ~(R2278_U68 & R2278_U313); 
assign R2278_U118 = ~(R2278_U69 & R2278_U311); 
assign R2278_U121 = ~(R2278_U70 & R2278_U309); 
assign R2278_U124 = ~(R2278_U232 & R2278_U233); 
assign R2278_U143 = ~(R2278_U280 & R2278_U30); 
assign R2278_U157 = R2278_U420 & R2278_U419; 
assign R2278_U248 = ~(R2278_U246 & R2278_U110); 
assign R2278_U321 = ~(R2278_U14 & R2278_U110); 
assign R2278_U324 = ~(R2278_U15 & R2278_U110); 
assign R2278_U327 = ~(R2278_U16 & R2278_U110); 
assign R2278_U330 = ~(R2278_U60 & R2278_U110); 
assign R2278_U348 = ~R2278_U110; 
assign R2278_U387 = ~(R2278_U264 & R2278_U110); 
assign R2278_U400 = ~(R2278_U346 & R2278_U127); 
assign R2278_U404 = ~(R2278_U344 & R2278_U131); 
assign R2278_U406 = ~(R2278_U342 & R2278_U134); 
assign R2278_U408 = ~(R2278_U340 & R2278_U137); 
assign R2278_U413 = ~(R2278_U279 & R2278_U147); 
assign R2358_U120 = ~(R2358_U650 & R2358_U649); 
assign R2358_U226 = ~(R2358_U349 & R2358_U329); 
assign R2358_U315 = ~R2358_U213; 
assign R2358_U318 = ~R2358_U68; 
assign R2358_U330 = ~R2358_U202; 
assign R2358_U331 = ~R2358_U208; 
assign R2358_U332 = ~(R2358_U151 & R2358_U208); 
assign R2358_U338 = ~(R2358_U5 & R2358_U208); 
assign R2358_U340 = ~(R2358_U152 & R2358_U208); 
assign R2358_U342 = ~(R2358_U208 & R2358_U293); 
assign R2358_U345 = ~(R2358_U433 & R2358_U155); 
assign R2358_U355 = ~R2358_U215; 
assign R2358_U356 = ~(R2358_U215 & R2358_U296); 
assign R2358_U360 = ~(R2358_U314 & R2358_U61); 
assign R2358_U365 = ~R2358_U72; 
assign R2358_U368 = ~(R2358_U72 & R2358_U224); 
assign R2358_U608 = ~(R2358_U180 & R2358_U202); 
assign R2358_U620 = ~(R2358_U390 & R2358_U208); 
assign R2358_U631 = ~(R2358_U394 & R2358_U68); 
assign R2358_U635 = ~(R2358_U396 & R2358_U213); 
assign R2358_U639 = ~(R2358_U398 & R2358_U215); 
assign R2358_U644 = ~(R2358_U399 & R2358_U72); 
assign R2099_U69 = ~(R2099_U305 & R2099_U304); 
assign R2099_U178 = ~R2099_U23; 
assign R2099_U303 = ~(R2099_U46 & R2099_U23); 
assign R2096_U74 = ~(R2096_U148 & R2096_U147); 
assign R2096_U119 = ~R2096_U56; 
assign R2096_U145 = ~(R2096_U56 & REIP_REG_28__SCAN_IN); 
assign ADD_405_U73 = ~(ADD_405_U150 & ADD_405_U149); 
assign ADD_405_U122 = ~ADD_405_U56; 
assign ADD_405_U147 = ~(ADD_405_U56 & INSTADDRPOINTER_REG_28__SCAN_IN); 
assign ADD_515_U74 = ~(ADD_515_U148 & ADD_515_U147); 
assign ADD_515_U119 = ~ADD_515_U56; 
assign ADD_515_U145 = ~(ADD_515_U56 & INSTADDRPOINTER_REG_28__SCAN_IN); 
assign U3002 = ~(U3804 & U3802 & U5670 & U5672); 
assign U3005 = ~(U3795 & U3793 & U5649 & U5651); 
assign U5637 = ~(R2278_U157 & U2377); 
assign U5740 = ~(R2099_U69 & U2380); 
assign U5750 = ~(ADD_405_U73 & U2375); 
assign U5751 = ~(ADD_515_U74 & U2374); 
assign U5843 = ~(U2372 & R2278_U157); 
assign U5855 = ~(R2358_U120 & U2364); 
assign U6182 = ~(U2386 & R2358_U120); 
assign U6292 = ~(U2383 & R2358_U120); 
assign U6332 = ~(U2371 & R2099_U69); 
assign U6457 = ~(U2367 & R2358_U120); 
assign U6544 = ~(U2604 & R2099_U69); 
assign U6552 = ~(R2096_U74 & U7473); 
assign R2278_U95 = ~(R2278_U61 & R2278_U330); 
assign R2278_U97 = ~(R2278_U329 & R2278_U327); 
assign R2278_U102 = ~(R2278_U326 & R2278_U324); 
assign R2278_U104 = ~(R2278_U323 & R2278_U321); 
assign R2278_U106 = ~(R2278_U36 & R2278_U248); 
assign R2278_U129 = R2278_U400 & R2278_U399; 
assign R2278_U133 = R2278_U404 & R2278_U403; 
assign R2278_U136 = R2278_U406 & R2278_U405; 
assign R2278_U139 = R2278_U408 & R2278_U407; 
assign R2278_U148 = R2278_U414 & R2278_U413; 
assign R2278_U234 = ~R2278_U124; 
assign R2278_U237 = ~R2278_U121; 
assign R2278_U239 = ~R2278_U118; 
assign R2278_U241 = ~R2278_U115; 
assign R2278_U244 = ~R2278_U112; 
assign R2278_U281 = ~R2278_U143; 
assign R2278_U388 = ~(R2278_U348 & R2278_U109); 
assign R2278_U390 = ~(R2278_U265 & R2278_U112); 
assign R2278_U392 = ~(R2278_U266 & R2278_U115); 
assign R2278_U394 = ~(R2278_U267 & R2278_U118); 
assign R2278_U396 = ~(R2278_U268 & R2278_U121); 
assign R2278_U398 = ~(R2278_U269 & R2278_U124); 
assign R2278_U412 = ~(R2278_U282 & R2278_U143); 
assign R2358_U17 = R2358_U360 & R2358_U359; 
assign R2358_U203 = ~(R2358_U292 & R2358_U332); 
assign R2358_U204 = ~(R2358_U338 & R2358_U337); 
assign R2358_U205 = ~(R2358_U153 & R2358_U340); 
assign R2358_U207 = ~(R2358_U283 & R2358_U342); 
assign R2358_U210 = ~(R2358_U345 & R2358_U437); 
assign R2358_U214 = ~(R2358_U356 & R2358_U59); 
assign R2358_U344 = ~(R2358_U154 & R2358_U342); 
assign R2358_U350 = ~(R2358_U326 & R2358_U226); 
assign R2358_U351 = ~(R2358_U318 & R2358_U46); 
assign R2358_U354 = ~(R2358_U226 & R2358_U353); 
assign R2358_U366 = ~(R2358_U365 & R2358_U227); 
assign R2358_U370 = ~(R2358_U161 & R2358_U368); 
assign R2358_U609 = ~(R2358_U330 & R2358_U508); 
assign R2358_U621 = ~(R2358_U102 & R2358_U331); 
assign R2358_U632 = ~(R2358_U630 & R2358_U318); 
assign R2358_U636 = ~(R2358_U113 & R2358_U315); 
assign R2358_U640 = ~(R2358_U117 & R2358_U355); 
assign R2358_U645 = ~(R2358_U643 & R2358_U365); 
assign R2099_U24 = ~(R2099_U178 & R2099_U46); 
assign R2099_U302 = ~(R2099_U231 & R2099_U178); 
assign R2096_U58 = ~(R2096_U119 & REIP_REG_28__SCAN_IN); 
assign R2096_U146 = ~(R2096_U119 & R2096_U57); 
assign ADD_405_U58 = ~(ADD_405_U122 & INSTADDRPOINTER_REG_28__SCAN_IN); 
assign ADD_405_U148 = ~(ADD_405_U122 & ADD_405_U57); 
assign ADD_515_U58 = ~(ADD_515_U119 & INSTADDRPOINTER_REG_28__SCAN_IN); 
assign ADD_515_U146 = ~(ADD_515_U119 & ADD_515_U57); 
assign U2814 = ~(U3901 & U6455 & U3900 & U6454 & U6457); 
assign U2846 = ~(U6293 & U6294 & U6292); 
assign U2878 = ~(U6183 & U6181 & U6182); 
assign U2973 = ~(U5854 & U5852 & U5856 & U5853 & U5855); 
assign U2975 = ~(U5844 & U5842 & U5846 & U5843 & U5845); 
assign U3007 = ~(U3787 & U3789 & U5637); 
assign U3835 = U5748 & U5750; 
assign U3837 = U3836 & U5751; 
assign U3928 = U6554 & U6552; 
assign U5658 = ~(R2278_U148 & U2377); 
assign U5679 = ~(R2278_U139 & U2377); 
assign U5686 = ~(R2278_U136 & U2377); 
assign U5693 = ~(R2278_U133 & U2377); 
assign U5700 = ~(R2278_U129 & U2377); 
assign U5858 = ~(U2372 & R2278_U148); 
assign U5870 = ~(R2358_U17 & U2364); 
assign U5873 = ~(U2372 & R2278_U139); 
assign U5878 = ~(U2372 & R2278_U136); 
assign U5883 = ~(U2372 & R2278_U133); 
assign U5888 = ~(U2372 & R2278_U129); 
assign U6192 = ~(U2386 & R2358_U17); 
assign U6301 = ~(U2383 & R2358_U17); 
assign U6478 = ~(U2367 & R2358_U17); 
assign R2278_U111 = R2278_U388 & R2278_U387; 
assign R2278_U249 = ~R2278_U106; 
assign R2278_U252 = ~R2278_U104; 
assign R2278_U255 = ~R2278_U102; 
assign R2278_U258 = ~R2278_U97; 
assign R2278_U261 = ~R2278_U95; 
assign R2278_U367 = ~(R2278_U62 & R2278_U95); 
assign R2278_U372 = ~(R2278_U63 & R2278_U97); 
assign R2278_U379 = ~(R2278_U64 & R2278_U102); 
assign R2278_U384 = ~(R2278_U65 & R2278_U104); 
assign R2278_U386 = ~(R2278_U263 & R2278_U106); 
assign R2278_U389 = ~(R2278_U244 & R2278_U113); 
assign R2278_U391 = ~(R2278_U241 & R2278_U116); 
assign R2278_U393 = ~(R2278_U239 & R2278_U119); 
assign R2278_U395 = ~(R2278_U237 & R2278_U122); 
assign R2278_U397 = ~(R2278_U234 & R2278_U125); 
assign R2278_U411 = ~(R2278_U281 & R2278_U144); 
assign R2358_U91 = ~(R2358_U609 & R2358_U608); 
assign R2358_U103 = ~(R2358_U621 & R2358_U620); 
assign R2358_U110 = ~(R2358_U632 & R2358_U631); 
assign R2358_U114 = ~(R2358_U636 & R2358_U635); 
assign R2358_U118 = ~(R2358_U640 & R2358_U639); 
assign R2358_U119 = ~(R2358_U645 & R2358_U644); 
assign R2358_U206 = ~(R2358_U344 & R2358_U285); 
assign R2358_U211 = ~(R2358_U350 & R2358_U325); 
assign R2358_U333 = ~R2358_U203; 
assign R2358_U339 = ~R2358_U204; 
assign R2358_U341 = ~R2358_U205; 
assign R2358_U343 = ~R2358_U207; 
assign R2358_U346 = ~R2358_U210; 
assign R2358_U347 = ~(R2358_U210 & R2358_U322); 
assign R2358_U352 = ~(R2358_U158 & R2358_U351); 
assign R2358_U357 = ~R2358_U214; 
assign R2358_U367 = ~(R2358_U160 & R2358_U366); 
assign R2358_U610 = ~(R2358_U385 & R2358_U203); 
assign R2358_U612 = ~(R2358_U386 & R2358_U204); 
assign R2358_U614 = ~(R2358_U387 & R2358_U205); 
assign R2358_U618 = ~(R2358_U389 & R2358_U207); 
assign R2358_U624 = ~(R2358_U392 & R2358_U210); 
assign R2358_U637 = ~(R2358_U397 & R2358_U214); 
assign R2099_U68 = ~(R2099_U303 & R2099_U302); 
assign R2099_U179 = ~R2099_U24; 
assign R2099_U301 = ~(R2099_U45 & R2099_U24); 
assign R2096_U73 = ~(R2096_U146 & R2096_U145); 
assign R2096_U120 = ~R2096_U58; 
assign R2096_U143 = ~(R2096_U58 & REIP_REG_29__SCAN_IN); 
assign ADD_405_U72 = ~(ADD_405_U148 & ADD_405_U147); 
assign ADD_405_U123 = ~ADD_405_U58; 
assign ADD_405_U145 = ~(ADD_405_U58 & INSTADDRPOINTER_REG_29__SCAN_IN); 
assign ADD_515_U73 = ~(ADD_515_U146 & ADD_515_U145); 
assign ADD_515_U120 = ~ADD_515_U58; 
assign ADD_515_U143 = ~(ADD_515_U58 & INSTADDRPOINTER_REG_29__SCAN_IN); 
assign U2811 = ~(U6476 & U6475 & U3907 & U3906 & U6478); 
assign U2843 = ~(U6302 & U6303 & U6301); 
assign U2875 = ~(U6191 & U6190 & U6193 & U6192); 
assign U2970 = ~(U5869 & U5867 & U5871 & U5868 & U5870); 
assign U2998 = ~(U3816 & U3814 & U5698 & U5700); 
assign U2999 = ~(U3813 & U3811 & U5691 & U5693); 
assign U3000 = ~(U3810 & U3808 & U5684 & U5686); 
assign U3001 = ~(U3807 & U3805 & U5677 & U5679); 
assign U3004 = ~(U3798 & U3796 & U5656 & U5658); 
assign U3466 = R2358_U91 & U4437; 
assign U5742 = ~(R2278_U111 & U2377); 
assign U5747 = ~(R2099_U68 & U2380); 
assign U5757 = ~(ADD_405_U72 & U2375); 
assign U5758 = ~(ADD_515_U73 & U2374); 
assign U5860 = ~(R2358_U119 & U2364); 
assign U5875 = ~(R2358_U118 & U2364); 
assign U5885 = ~(R2358_U114 & U2364); 
assign U5890 = ~(R2358_U110 & U2364); 
assign U5915 = ~(R2358_U103 & U2364); 
assign U5918 = ~(U2372 & R2278_U111); 
assign U5945 = ~(R2358_U91 & U2364); 
assign U6185 = ~(U2386 & R2358_U119); 
assign U6196 = ~(U2386 & R2358_U118); 
assign U6204 = ~(U2386 & R2358_U114); 
assign U6208 = ~(U2386 & R2358_U110); 
assign U6228 = ~(U2386 & R2358_U103); 
assign U6295 = ~(U2383 & R2358_U119); 
assign U6304 = ~(U2383 & R2358_U118); 
assign U6310 = ~(U2383 & R2358_U114); 
assign U6313 = ~(U2383 & R2358_U110); 
assign U6328 = ~(U2383 & R2358_U103); 
assign U6335 = ~(U2371 & R2099_U68); 
assign U6464 = ~(U2367 & R2358_U119); 
assign U6485 = ~(U2367 & R2358_U118); 
assign U6499 = ~(U2367 & R2358_U114); 
assign U6506 = ~(U2367 & R2358_U110); 
assign U6541 = ~(U2367 & R2358_U103); 
assign U6551 = ~(U2604 & R2099_U68); 
assign U6559 = ~(R2096_U73 & U7473); 
assign U6583 = ~(U2367 & R2358_U91); 
assign R2278_U114 = R2278_U390 & R2278_U389; 
assign R2278_U117 = R2278_U392 & R2278_U391; 
assign R2278_U120 = R2278_U394 & R2278_U393; 
assign R2278_U123 = R2278_U396 & R2278_U395; 
assign R2278_U126 = R2278_U398 & R2278_U397; 
assign R2278_U145 = R2278_U412 & R2278_U411; 
assign R2278_U366 = ~(R2278_U261 & R2278_U365); 
assign R2278_U371 = ~(R2278_U258 & R2278_U370); 
assign R2278_U378 = ~(R2278_U255 & R2278_U377); 
assign R2278_U383 = ~(R2278_U252 & R2278_U382); 
assign R2278_U385 = ~(R2278_U249 & R2278_U107); 
assign R2358_U16 = R2358_U370 & R2358_U367; 
assign R2358_U18 = R2358_U354 & R2358_U352; 
assign R2358_U209 = ~(R2358_U321 & R2358_U347); 
assign R2358_U220 = ~R2358_U211; 
assign R2358_U221 = ~R2358_U206; 
assign R2358_U611 = ~(R2358_U92 & R2358_U333); 
assign R2358_U613 = ~(R2358_U94 & R2358_U339); 
assign R2358_U615 = ~(R2358_U96 & R2358_U341); 
assign R2358_U617 = ~(R2358_U98 & R2358_U206); 
assign R2358_U619 = ~(R2358_U100 & R2358_U343); 
assign R2358_U625 = ~(R2358_U106 & R2358_U346); 
assign R2358_U627 = ~(R2358_U108 & R2358_U211); 
assign R2358_U638 = ~(R2358_U115 & R2358_U357); 
assign R2099_U25 = ~(R2099_U179 & R2099_U45); 
assign R2099_U300 = ~(R2099_U228 & R2099_U179); 
assign R2096_U60 = ~(R2096_U120 & REIP_REG_29__SCAN_IN); 
assign R2096_U144 = ~(R2096_U120 & R2096_U59); 
assign ADD_405_U60 = ~(ADD_405_U123 & INSTADDRPOINTER_REG_29__SCAN_IN); 
assign ADD_405_U146 = ~(ADD_405_U123 & ADD_405_U59); 
assign ADD_515_U60 = ~(ADD_515_U120 & INSTADDRPOINTER_REG_29__SCAN_IN); 
assign ADD_515_U144 = ~(ADD_515_U120 & ADD_515_U59); 
assign U2802 = ~(U6539 & U3924 & U3925 & U6537 & U6541); 
assign U2807 = ~(U6504 & U3914 & U3915 & U6502 & U6506); 
assign U2808 = ~(U3912 & U6497 & U3913 & U6495 & U6499); 
assign U2810 = ~(U3908 & U6483 & U3909 & U6481 & U6485); 
assign U2813 = ~(U3903 & U6462 & U3902 & U6461 & U6464); 
assign U2834 = ~(U6329 & U6330 & U6328); 
assign U2839 = ~(U6314 & U6315 & U6313); 
assign U2840 = ~(U6311 & U6312 & U6310); 
assign U2842 = ~(U6305 & U6306 & U6304); 
assign U2845 = ~(U6296 & U6297 & U6295); 
assign U2866 = ~(U6227 & U6226 & U6229 & U6228); 
assign U2871 = ~(U6207 & U6206 & U6209 & U6208); 
assign U2872 = ~(U6203 & U6202 & U6205 & U6204); 
assign U2874 = ~(U6195 & U6194 & U6197 & U6196); 
assign U2877 = ~(U6186 & U6184 & U6185); 
assign U2966 = ~(U5889 & U5887 & U5891 & U5888 & U5890); 
assign U2967 = ~(U5884 & U5882 & U5886 & U5883 & U5885); 
assign U2969 = ~(U5874 & U5872 & U5876 & U5873 & U5875); 
assign U2972 = ~(U5859 & U5857 & U5861 & U5858 & U5860); 
assign U2992 = ~(U3834 & U3832 & U5740 & U5742); 
assign U3838 = U5755 & U5757; 
assign U3840 = U3839 & U5758; 
assign U3930 = U6561 & U6559; 
assign U5665 = ~(R2278_U145 & U2377); 
assign U5707 = ~(R2278_U126 & U2377); 
assign U5714 = ~(R2278_U123 & U2377); 
assign U5721 = ~(R2278_U120 & U2377); 
assign U5728 = ~(R2278_U117 & U2377); 
assign U5735 = ~(R2278_U114 & U2377); 
assign U5863 = ~(U2372 & R2278_U145); 
assign U5865 = ~(R2358_U16 & U2364); 
assign U5893 = ~(U2372 & R2278_U126); 
assign U5895 = ~(R2358_U18 & U2364); 
assign U5898 = ~(U2372 & R2278_U123); 
assign U5903 = ~(U2372 & R2278_U120); 
assign U5908 = ~(U2372 & R2278_U117); 
assign U5913 = ~(U2372 & R2278_U114); 
assign U6188 = ~(U2386 & R2358_U16); 
assign U6212 = ~(U2386 & R2358_U18); 
assign U6298 = ~(U2383 & R2358_U16); 
assign U6316 = ~(U2383 & R2358_U18); 
assign U6471 = ~(U2367 & R2358_U16); 
assign U6513 = ~(U2367 & R2358_U18); 
assign U7733 = ~(U3466 & U4211); 
assign R2278_U96 = R2278_U367 & R2278_U366; 
assign R2278_U98 = R2278_U372 & R2278_U371; 
assign R2278_U103 = R2278_U379 & R2278_U378; 
assign R2278_U105 = R2278_U384 & R2278_U383; 
assign R2278_U108 = R2278_U386 & R2278_U385; 
assign R2358_U93 = ~(R2358_U611 & R2358_U610); 
assign R2358_U95 = ~(R2358_U613 & R2358_U612); 
assign R2358_U97 = ~(R2358_U615 & R2358_U614); 
assign R2358_U101 = ~(R2358_U619 & R2358_U618); 
assign R2358_U107 = ~(R2358_U625 & R2358_U624); 
assign R2358_U116 = ~(R2358_U638 & R2358_U637); 
assign R2358_U348 = ~R2358_U209; 
assign R2358_U616 = ~(R2358_U221 & R2358_U388); 
assign R2358_U622 = ~(R2358_U391 & R2358_U209); 
assign R2358_U626 = ~(R2358_U220 & R2358_U393); 
assign R2099_U67 = ~(R2099_U301 & R2099_U300); 
assign R2099_U180 = ~R2099_U25; 
assign R2099_U299 = ~(R2099_U44 & R2099_U25); 
assign R2096_U72 = ~(R2096_U144 & R2096_U143); 
assign R2096_U121 = ~R2096_U60; 
assign R2096_U139 = ~(R2096_U60 & REIP_REG_30__SCAN_IN); 
assign ADD_405_U71 = ~(ADD_405_U146 & ADD_405_U145); 
assign ADD_405_U124 = ~ADD_405_U60; 
assign ADD_405_U143 = ~(ADD_405_U60 & INSTADDRPOINTER_REG_30__SCAN_IN); 
assign ADD_515_U72 = ~(ADD_515_U144 & ADD_515_U143); 
assign ADD_515_U121 = ~ADD_515_U60; 
assign ADD_515_U139 = ~(ADD_515_U60 & INSTADDRPOINTER_REG_30__SCAN_IN); 
assign U2806 = ~(U6511 & U3916 & U3917 & U6509 & U6513); 
assign U2812 = ~(U6469 & U6468 & U3905 & U3904 & U6471); 
assign U2838 = ~(U6317 & U6318 & U6316); 
assign U2844 = ~(U6299 & U6300 & U6298); 
assign U2870 = ~(U6211 & U6210 & U6213 & U6212); 
assign U2876 = ~(U6189 & U6187 & U6188); 
assign U2961 = ~(U5914 & U5912 & U5916 & U5913 & U5915); 
assign U2965 = ~(U5894 & U5892 & U5896 & U5893 & U5895); 
assign U2971 = ~(U5864 & U5862 & U5866 & U5863 & U5865); 
assign U2993 = ~(U3831 & U3829 & U5733 & U5735); 
assign U2994 = ~(U3828 & U3826 & U5726 & U5728); 
assign U2995 = ~(U3825 & U3823 & U5719 & U5721); 
assign U2996 = ~(U3822 & U3820 & U5712 & U5714); 
assign U2997 = ~(U3819 & U3817 & U5705 & U5707); 
assign U3003 = ~(U3801 & U3799 & U5663 & U5665); 
assign U4164 = U7733 & U7732; 
assign U5749 = ~(R2278_U108 & U2377); 
assign U5754 = ~(R2099_U67 & U2380); 
assign U5756 = ~(R2278_U105 & U2377); 
assign U5763 = ~(R2278_U103 & U2377); 
assign U5764 = ~(ADD_405_U71 & U2375); 
assign U5765 = ~(ADD_515_U72 & U2374); 
assign U5770 = ~(R2278_U98 & U2377); 
assign U5777 = ~(R2278_U96 & U2377); 
assign U5880 = ~(R2358_U116 & U2364); 
assign U5905 = ~(R2358_U107 & U2364); 
assign U5920 = ~(R2358_U101 & U2364); 
assign U5923 = ~(U2372 & R2278_U108); 
assign U5928 = ~(U2372 & R2278_U105); 
assign U5930 = ~(R2358_U97 & U2364); 
assign U5933 = ~(U2372 & R2278_U103); 
assign U5935 = ~(R2358_U95 & U2364); 
assign U5938 = ~(U2372 & R2278_U98); 
assign U5940 = ~(R2358_U93 & U2364); 
assign U5943 = ~(U2372 & R2278_U96); 
assign U6200 = ~(U2386 & R2358_U116); 
assign U6220 = ~(U2386 & R2358_U107); 
assign U6232 = ~(U2386 & R2358_U101); 
assign U6240 = ~(U2386 & R2358_U97); 
assign U6244 = ~(U2386 & R2358_U95); 
assign U6248 = ~(U2386 & R2358_U93); 
assign U6307 = ~(U2383 & R2358_U116); 
assign U6322 = ~(U2383 & R2358_U107); 
assign U6331 = ~(U2383 & R2358_U101); 
assign U6337 = ~(U2383 & R2358_U97); 
assign U6338 = ~(U2371 & R2099_U67); 
assign U6340 = ~(U2383 & R2358_U95); 
assign U6343 = ~(U2383 & R2358_U93); 
assign U6492 = ~(U2367 & R2358_U116); 
assign U6527 = ~(U2367 & R2358_U107); 
assign U6548 = ~(U2367 & R2358_U101); 
assign U6558 = ~(U2604 & R2099_U67); 
assign U6562 = ~(U2367 & R2358_U97); 
assign U6566 = ~(R2096_U72 & U7473); 
assign U6569 = ~(U2367 & R2358_U95); 
assign U6576 = ~(U2367 & R2358_U93); 
assign R2358_U99 = ~(R2358_U617 & R2358_U616); 
assign R2358_U109 = ~(R2358_U627 & R2358_U626); 
assign R2358_U623 = ~(R2358_U104 & R2358_U348); 
assign R2099_U135 = ~(R2099_U96 & R2099_U180); 
assign R2099_U136 = ~(R2099_U180 & R2099_U44); 
assign R2099_U298 = ~(R2099_U288 & R2099_U180); 
assign R2096_U93 = ~(R2096_U121 & REIP_REG_30__SCAN_IN); 
assign R2096_U140 = ~(R2096_U121 & R2096_U61); 
assign ADD_405_U95 = ~(ADD_405_U124 & INSTADDRPOINTER_REG_30__SCAN_IN); 
assign ADD_405_U144 = ~(ADD_405_U124 & ADD_405_U61); 
assign ADD_515_U93 = ~(ADD_515_U121 & INSTADDRPOINTER_REG_30__SCAN_IN); 
assign ADD_515_U140 = ~(ADD_515_U121 & ADD_515_U61); 
assign U2799 = ~(U6560 & U3930 & U3931 & U6558 & U6562); 
assign U2801 = ~(U6546 & U3926 & U3927 & U6544 & U6548); 
assign U2804 = ~(U6525 & U3920 & U3921 & U6523 & U6527); 
assign U2809 = ~(U3910 & U6490 & U3911 & U6488 & U6492); 
assign U2831 = ~(U6338 & U6339 & U6337); 
assign U2833 = ~(U6332 & U6333 & U6331); 
assign U2836 = ~(U6323 & U6324 & U6322); 
assign U2841 = ~(U6308 & U6309 & U6307); 
assign U2860 = ~(U4164 & U6250); 
assign U2861 = ~(U6247 & U6246 & U6249 & U6248); 
assign U2862 = ~(U6243 & U6242 & U6245 & U6244); 
assign U2863 = ~(U6239 & U6238 & U6241 & U6240); 
assign U2865 = ~(U6231 & U6230 & U6233 & U6232); 
assign U2868 = ~(U6219 & U6218 & U6221 & U6220); 
assign U2873 = ~(U6199 & U6198 & U6201 & U6200); 
assign U2955 = ~(U5944 & U5942 & U5946 & U5943 & U5945); 
assign U2956 = ~(U5939 & U5937 & U5941 & U5938 & U5940); 
assign U2957 = ~(U5934 & U5932 & U5936 & U5933 & U5935); 
assign U2958 = ~(U5929 & U5927 & U5931 & U5928 & U5930); 
assign U2960 = ~(U5919 & U5917 & U5921 & U5918 & U5920); 
assign U2963 = ~(U5904 & U5902 & U5906 & U5903 & U5905); 
assign U2968 = ~(U5879 & U5877 & U5881 & U5878 & U5880); 
assign U2990 = ~(U3840 & U3838 & U5754 & U5756); 
assign U2991 = ~(U3837 & U3835 & U5747 & U5749); 
assign U3841 = U5762 & U5764; 
assign U3843 = U3842 & U5765; 
assign U3932 = U6568 & U6566; 
assign U5900 = ~(R2358_U109 & U2364); 
assign U5925 = ~(R2358_U99 & U2364); 
assign U6216 = ~(U2386 & R2358_U109); 
assign U6236 = ~(U2386 & R2358_U99); 
assign U6319 = ~(U2383 & R2358_U109); 
assign U6334 = ~(U2383 & R2358_U99); 
assign U6520 = ~(U2367 & R2358_U109); 
assign U6555 = ~(U2367 & R2358_U99); 
assign R2358_U105 = ~(R2358_U623 & R2358_U622); 
assign R2099_U66 = ~(R2099_U299 & R2099_U298); 
assign R2099_U145 = ~R2099_U135; 
assign R2099_U181 = ~R2099_U136; 
assign R2099_U293 = ~(R2099_U97 & R2099_U135); 
assign R2099_U295 = ~(R2099_U43 & R2099_U136); 
assign R2096_U70 = ~(R2096_U140 & R2096_U139); 
assign R2096_U122 = ~R2096_U93; 
assign R2096_U137 = ~(R2096_U93 & REIP_REG_31__SCAN_IN); 
assign ADD_405_U70 = ~(ADD_405_U144 & ADD_405_U143); 
assign ADD_405_U125 = ~ADD_405_U95; 
assign ADD_405_U141 = ~(ADD_405_U95 & INSTADDRPOINTER_REG_31__SCAN_IN); 
assign ADD_515_U70 = ~(ADD_515_U140 & ADD_515_U139); 
assign ADD_515_U122 = ~ADD_515_U93; 
assign ADD_515_U137 = ~(ADD_515_U93 & INSTADDRPOINTER_REG_31__SCAN_IN); 
assign U2800 = ~(U6553 & U3928 & U3929 & U6551 & U6555); 
assign U2805 = ~(U6518 & U3918 & U3919 & U6516 & U6520); 
assign U2832 = ~(U6335 & U6336 & U6334); 
assign U2837 = ~(U6320 & U6321 & U6319); 
assign U2864 = ~(U6235 & U6234 & U6237 & U6236); 
assign U2869 = ~(U6215 & U6214 & U6217 & U6216); 
assign U2959 = ~(U5924 & U5922 & U5926 & U5923 & U5925); 
assign U2964 = ~(U5899 & U5897 & U5901 & U5898 & U5900); 
assign U5761 = ~(R2099_U66 & U2380); 
assign U5771 = ~(ADD_405_U70 & U2375); 
assign U5772 = ~(ADD_515_U70 & U2374); 
assign U5910 = ~(R2358_U105 & U2364); 
assign U6224 = ~(U2386 & R2358_U105); 
assign U6325 = ~(U2383 & R2358_U105); 
assign U6341 = ~(U2371 & R2099_U66); 
assign U6534 = ~(U2367 & R2358_U105); 
assign U6565 = ~(U2604 & R2099_U66); 
assign U6573 = ~(R2096_U70 & U7473); 
assign R2099_U292 = ~(R2099_U145 & R2099_U291); 
assign R2099_U294 = ~(R2099_U181 & R2099_U285); 
assign R2096_U138 = ~(R2096_U122 & R2096_U92); 
assign ADD_405_U142 = ~(ADD_405_U125 & ADD_405_U94); 
assign ADD_515_U138 = ~(ADD_515_U122 & ADD_515_U92); 
assign U2798 = ~(U6567 & U3932 & U3933 & U6565 & U6569); 
assign U2803 = ~(U6532 & U3922 & U3923 & U6530 & U6534); 
assign U2830 = ~(U6341 & U6342 & U6340); 
assign U2835 = ~(U6326 & U6327 & U6325); 
assign U2867 = ~(U6223 & U6222 & U6225 & U6224); 
assign U2962 = ~(U5909 & U5907 & U5911 & U5908 & U5910); 
assign U2989 = ~(U3843 & U3841 & U5761 & U5763); 
assign U3844 = U5769 & U5771; 
assign U3846 = U3845 & U5772; 
assign U3934 = U6575 & U6573; 
assign R2099_U64 = ~(R2099_U293 & R2099_U292); 
assign R2099_U65 = ~(R2099_U295 & R2099_U294); 
assign R2096_U69 = ~(R2096_U138 & R2096_U137); 
assign ADD_405_U69 = ~(ADD_405_U142 & ADD_405_U141); 
assign ADD_515_U69 = ~(ADD_515_U138 & ADD_515_U137); 
assign U5768 = ~(R2099_U65 & U2380); 
assign U5775 = ~(R2099_U64 & U2380); 
assign U5778 = ~(ADD_405_U69 & U2375); 
assign U5779 = ~(ADD_515_U69 & U2374); 
assign U6344 = ~(U2371 & R2099_U65); 
assign U6346 = ~(U2371 & R2099_U64); 
assign U6572 = ~(U2604 & R2099_U65); 
assign U6579 = ~(U2604 & R2099_U64); 
assign U6580 = ~(R2096_U69 & U7473); 
assign U2797 = ~(U6574 & U3934 & U3935 & U6572 & U6576); 
assign U2828 = ~(U6347 & U6346); 
assign U2829 = ~(U6344 & U6345 & U6343); 
assign U2988 = ~(U3846 & U3844 & U5768 & U5770); 
assign U3847 = U5776 & U5778; 
assign U3849 = U3848 & U5779; 
assign U3936 = U6582 & U6580; 
assign U2796 = ~(U6581 & U3936 & U3937 & U6579 & U6583); 
assign U2987 = ~(U3849 & U3847 & U5775 & U5777); 
endmodule 
