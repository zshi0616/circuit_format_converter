module b03_C( STATO_REG_0__SCAN_IN, REQUEST1, REQUEST2, REQUEST3, REQUEST4, CODA0_REG_2__SCAN_IN, CODA0_REG_1__SCAN_IN, CODA0_REG_0__SCAN_IN, CODA1_REG_2__SCAN_IN, CODA1_REG_1__SCAN_IN, CODA1_REG_0__SCAN_IN, CODA2_REG_2__SCAN_IN, CODA2_REG_1__SCAN_IN, CODA2_REG_0__SCAN_IN, CODA3_REG_2__SCAN_IN, CODA3_REG_1__SCAN_IN, CODA3_REG_0__SCAN_IN, GRANT_REG_3__SCAN_IN, GRANT_REG_2__SCAN_IN, GRANT_REG_1__SCAN_IN, GRANT_REG_0__SCAN_IN, GRANT_O_REG_3__SCAN_IN, GRANT_O_REG_2__SCAN_IN, GRANT_O_REG_1__SCAN_IN, GRANT_O_REG_0__SCAN_IN, RU3_REG_SCAN_IN, FU1_REG_SCAN_IN, FU3_REG_SCAN_IN, RU1_REG_SCAN_IN, RU4_REG_SCAN_IN, FU2_REG_SCAN_IN, FU4_REG_SCAN_IN, RU2_REG_SCAN_IN, STATO_REG_1__SCAN_IN, U204, U205, U206, U207, U208, U209, U210, U211, U212, U213, U214, U215, U216, U217, U229, U230, U231, U232, U233, U234, U235, U236, U237, U238, U239, U240, U241, U242); 
input STATO_REG_0__SCAN_IN, REQUEST1, REQUEST2, REQUEST3, REQUEST4, CODA0_REG_2__SCAN_IN, CODA0_REG_1__SCAN_IN, CODA0_REG_0__SCAN_IN, CODA1_REG_2__SCAN_IN, CODA1_REG_1__SCAN_IN, CODA1_REG_0__SCAN_IN, CODA2_REG_2__SCAN_IN, CODA2_REG_1__SCAN_IN, CODA2_REG_0__SCAN_IN, CODA3_REG_2__SCAN_IN, CODA3_REG_1__SCAN_IN, CODA3_REG_0__SCAN_IN, GRANT_REG_3__SCAN_IN, GRANT_REG_2__SCAN_IN, GRANT_REG_1__SCAN_IN, GRANT_REG_0__SCAN_IN, GRANT_O_REG_3__SCAN_IN, GRANT_O_REG_2__SCAN_IN, GRANT_O_REG_1__SCAN_IN, GRANT_O_REG_0__SCAN_IN, RU3_REG_SCAN_IN, FU1_REG_SCAN_IN, FU3_REG_SCAN_IN, RU1_REG_SCAN_IN, RU4_REG_SCAN_IN, FU2_REG_SCAN_IN, FU4_REG_SCAN_IN, RU2_REG_SCAN_IN, STATO_REG_1__SCAN_IN; 
output U204, U205, U206, U207, U208, U209, U210, U211, U212, U213, U214, U215, U216, U217, U229, U230, U231, U232, U233, U234, U235, U236, U237, U238, U239, U240, U241, U242; 
wire U201, U202, U203, U218, U219, U220, U221, U222, U223, U224, U225, U226, U227, U228, U243, U244, U245, U246, U247, U248, U249, U250, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, U280, U281, U282, U283, U284, U285, U286, U287, U288, U289, U290, U291, U292, U293, U294, U295, U296, U297, U298, U299, U300, U301, U302, U303, U304, U305, U306, U307, U308, U309, U310, U311, U312, U313, U314, U315, U316, U317, U318, U319, U320, U321, U322; 
assign U203 = ~STATO_REG_0__SCAN_IN; 
assign U218 = ~STATO_REG_1__SCAN_IN; 
assign U219 = ~RU3_REG_SCAN_IN; 
assign U221 = ~RU1_REG_SCAN_IN; 
assign U222 = ~(RU1_REG_SCAN_IN & STATO_REG_0__SCAN_IN); 
assign U224 = ~CODA0_REG_2__SCAN_IN; 
assign U225 = ~CODA0_REG_1__SCAN_IN; 
assign U226 = ~CODA0_REG_0__SCAN_IN; 
assign U227 = ~FU1_REG_SCAN_IN; 
assign U228 = ~FU2_REG_SCAN_IN; 
assign U243 = ~RU2_REG_SCAN_IN; 
assign U245 = ~FU3_REG_SCAN_IN; 
assign U246 = ~FU4_REG_SCAN_IN; 
assign U248 = FU1_REG_SCAN_IN | FU3_REG_SCAN_IN | FU2_REG_SCAN_IN | FU4_REG_SCAN_IN; 
assign U256 = RU3_REG_SCAN_IN | RU2_REG_SCAN_IN; 
assign U304 = ~(GRANT_REG_3__SCAN_IN & STATO_REG_0__SCAN_IN); 
assign U306 = ~(GRANT_REG_2__SCAN_IN & STATO_REG_0__SCAN_IN); 
assign U308 = ~(GRANT_REG_1__SCAN_IN & STATO_REG_0__SCAN_IN); 
assign U310 = ~(GRANT_REG_0__SCAN_IN & STATO_REG_0__SCAN_IN); 
assign U312 = ~(RU3_REG_SCAN_IN & STATO_REG_0__SCAN_IN); 
assign U314 = ~(RU3_REG_SCAN_IN & STATO_REG_0__SCAN_IN); 
assign U316 = ~(RU4_REG_SCAN_IN & STATO_REG_0__SCAN_IN); 
assign U318 = ~(RU2_REG_SCAN_IN & STATO_REG_0__SCAN_IN); 
assign U320 = ~(RU4_REG_SCAN_IN & STATO_REG_0__SCAN_IN); 
assign U322 = ~(RU2_REG_SCAN_IN & STATO_REG_0__SCAN_IN); 
assign U220 = ~(U243 & RU3_REG_SCAN_IN); 
assign U244 = ~(U248 & STATO_REG_1__SCAN_IN); 
assign U247 = ~U222; 
assign U257 = ~(U221 & U256); 
assign U291 = ~(U203 & FU1_REG_SCAN_IN); 
assign U292 = ~(REQUEST1 & U203); 
assign U293 = ~(U228 & RU2_REG_SCAN_IN); 
assign U294 = ~(U219 & U246 & U243 & RU4_REG_SCAN_IN); 
assign U303 = ~(U203 & GRANT_O_REG_3__SCAN_IN); 
assign U305 = ~(U203 & GRANT_O_REG_2__SCAN_IN); 
assign U307 = ~(U203 & GRANT_O_REG_1__SCAN_IN); 
assign U309 = ~(U203 & GRANT_O_REG_0__SCAN_IN); 
assign U311 = ~(REQUEST3 & U203); 
assign U313 = ~(U203 & FU3_REG_SCAN_IN); 
assign U315 = ~(REQUEST4 & U203); 
assign U317 = ~(U203 & FU2_REG_SCAN_IN); 
assign U319 = ~(U203 & FU4_REG_SCAN_IN); 
assign U321 = ~(REQUEST2 & U203); 
assign U204 = ~(U222 & U292); 
assign U205 = ~(U222 & U291); 
assign U233 = ~(U304 & U303); 
assign U234 = ~(U306 & U305); 
assign U235 = ~(U308 & U307); 
assign U236 = ~(U310 & U309); 
assign U237 = ~(U312 & U311); 
assign U238 = ~(U314 & U313); 
assign U239 = ~(U316 & U315); 
assign U240 = ~(U318 & U317); 
assign U241 = ~(U320 & U319); 
assign U242 = ~(U322 & U321); 
assign U249 = ~U244; 
assign U250 = ~U220; 
assign U254 = ~(U247 & U227); 
assign U295 = ~(U244 & GRANT_REG_3__SCAN_IN); 
assign U297 = ~(U244 & GRANT_REG_2__SCAN_IN); 
assign U299 = ~(U244 & GRANT_REG_1__SCAN_IN); 
assign U301 = ~(U244 & GRANT_REG_0__SCAN_IN); 
assign U251 = ~(U250 & U245); 
assign U296 = ~(U226 & U225 & U249 & CODA0_REG_2__SCAN_IN); 
assign U298 = ~(U226 & U224 & U249 & CODA0_REG_1__SCAN_IN); 
assign U300 = ~(U225 & U224 & U249 & CODA0_REG_0__SCAN_IN); 
assign U302 = ~(U249 & CODA0_REG_2__SCAN_IN & CODA0_REG_1__SCAN_IN & CODA0_REG_0__SCAN_IN); 
assign U229 = ~(U296 & U295); 
assign U230 = ~(U298 & U297); 
assign U231 = ~(U300 & U299); 
assign U232 = ~(U302 & U301); 
assign U252 = ~(U294 & U293 & U251); 
assign U253 = ~(U221 & U252 & STATO_REG_0__SCAN_IN); 
assign U223 = ~(U254 & U244 & U253); 
assign U201 = U223 & U218; 
assign U202 = U223 & STATO_REG_1__SCAN_IN; 
assign U255 = ~U223; 
assign U258 = ~(U201 & U257); 
assign U259 = ~(U202 & CODA1_REG_2__SCAN_IN); 
assign U260 = ~(U255 & CODA0_REG_2__SCAN_IN); 
assign U261 = ~(U220 & U221 & U201); 
assign U262 = ~(U202 & CODA1_REG_1__SCAN_IN); 
assign U263 = ~(U255 & CODA0_REG_1__SCAN_IN); 
assign U264 = ~(U221 & U243 & U201); 
assign U265 = ~(U202 & CODA1_REG_0__SCAN_IN); 
assign U266 = ~(U255 & CODA0_REG_0__SCAN_IN); 
assign U267 = ~(U202 & CODA2_REG_2__SCAN_IN); 
assign U268 = ~(U201 & CODA0_REG_2__SCAN_IN); 
assign U269 = ~(U255 & CODA1_REG_2__SCAN_IN); 
assign U270 = ~(U202 & CODA2_REG_1__SCAN_IN); 
assign U271 = ~(U201 & CODA0_REG_1__SCAN_IN); 
assign U272 = ~(U255 & CODA1_REG_1__SCAN_IN); 
assign U273 = ~(U202 & CODA2_REG_0__SCAN_IN); 
assign U274 = ~(U201 & CODA0_REG_0__SCAN_IN); 
assign U275 = ~(U255 & CODA1_REG_0__SCAN_IN); 
assign U276 = ~(U202 & CODA3_REG_2__SCAN_IN); 
assign U277 = ~(U201 & CODA1_REG_2__SCAN_IN); 
assign U278 = ~(U255 & CODA2_REG_2__SCAN_IN); 
assign U279 = ~(U202 & CODA3_REG_1__SCAN_IN); 
assign U280 = ~(U201 & CODA1_REG_1__SCAN_IN); 
assign U281 = ~(U255 & CODA2_REG_1__SCAN_IN); 
assign U282 = ~(U202 & CODA3_REG_0__SCAN_IN); 
assign U283 = ~(U201 & CODA1_REG_0__SCAN_IN); 
assign U284 = ~(U255 & CODA2_REG_0__SCAN_IN); 
assign U285 = ~(U201 & CODA2_REG_2__SCAN_IN); 
assign U286 = ~(U255 & CODA3_REG_2__SCAN_IN); 
assign U287 = ~(U201 & CODA2_REG_1__SCAN_IN); 
assign U288 = ~(U255 & CODA3_REG_1__SCAN_IN); 
assign U289 = ~(U201 & CODA2_REG_0__SCAN_IN); 
assign U290 = ~(U255 & CODA3_REG_0__SCAN_IN); 
assign U206 = ~(U290 & U289); 
assign U207 = ~(U288 & U287); 
assign U208 = ~(U286 & U285); 
assign U209 = ~(U283 & U282 & U284); 
assign U210 = ~(U280 & U279 & U281); 
assign U211 = ~(U277 & U276 & U278); 
assign U212 = ~(U274 & U273 & U275); 
assign U213 = ~(U271 & U270 & U272); 
assign U214 = ~(U268 & U267 & U269); 
assign U215 = ~(U265 & U264 & U266); 
assign U216 = ~(U262 & U261 & U263); 
assign U217 = ~(U259 & U258 & U260); 
endmodule 
